magic
tech sky130A
magscale 1 2
timestamp 1654258643
<< viali >>
rect 14289 47209 14323 47243
rect 22477 47209 22511 47243
rect 44097 47209 44131 47243
rect 3065 47141 3099 47175
rect 29929 47141 29963 47175
rect 47961 47141 47995 47175
rect 12357 47073 12391 47107
rect 12633 47073 12667 47107
rect 30757 47073 30791 47107
rect 47041 47073 47075 47107
rect 1777 47005 1811 47039
rect 3801 47005 3835 47039
rect 4721 47005 4755 47039
rect 6377 47005 6411 47039
rect 7297 47005 7331 47039
rect 9413 47005 9447 47039
rect 14105 47005 14139 47039
rect 14933 47005 14967 47039
rect 16681 47005 16715 47039
rect 16957 47005 16991 47039
rect 21005 47005 21039 47039
rect 22017 47005 22051 47039
rect 22661 47005 22695 47039
rect 24869 47005 24903 47039
rect 28549 47005 28583 47039
rect 29745 47005 29779 47039
rect 31033 47005 31067 47039
rect 38393 47005 38427 47039
rect 41521 47005 41555 47039
rect 42717 47005 42751 47039
rect 43269 47005 43303 47039
rect 43913 47005 43947 47039
rect 45201 47005 45235 47039
rect 47777 47005 47811 47039
rect 2053 46937 2087 46971
rect 2789 46937 2823 46971
rect 4077 46937 4111 46971
rect 4997 46937 5031 46971
rect 6653 46937 6687 46971
rect 9597 46937 9631 46971
rect 15117 46937 15151 46971
rect 19717 46937 19751 46971
rect 20085 46937 20119 46971
rect 28733 46937 28767 46971
rect 40325 46937 40359 46971
rect 40509 46937 40543 46971
rect 43453 46937 43487 46971
rect 45385 46937 45419 46971
rect 7481 46869 7515 46903
rect 1869 46597 1903 46631
rect 5825 46597 5859 46631
rect 19441 46529 19475 46563
rect 24593 46529 24627 46563
rect 38117 46529 38151 46563
rect 42441 46529 42475 46563
rect 47961 46529 47995 46563
rect 3985 46461 4019 46495
rect 4169 46461 4203 46495
rect 10977 46461 11011 46495
rect 11529 46461 11563 46495
rect 11713 46461 11747 46495
rect 11989 46461 12023 46495
rect 13829 46461 13863 46495
rect 14013 46461 14047 46495
rect 14289 46461 14323 46495
rect 19625 46461 19659 46495
rect 20637 46461 20671 46495
rect 24777 46461 24811 46495
rect 25145 46461 25179 46495
rect 32229 46461 32263 46495
rect 32413 46461 32447 46495
rect 32689 46461 32723 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46857 46461 46891 46495
rect 2145 46325 2179 46359
rect 41337 46325 41371 46359
rect 48053 46325 48087 46359
rect 4537 46121 4571 46155
rect 5181 46121 5215 46155
rect 13553 46121 13587 46155
rect 14197 46121 14231 46155
rect 19901 46121 19935 46155
rect 24685 46121 24719 46155
rect 32505 46121 32539 46155
rect 38301 46121 38335 46155
rect 11713 45985 11747 46019
rect 20821 45985 20855 46019
rect 21281 45985 21315 46019
rect 25789 45985 25823 46019
rect 41061 45985 41095 46019
rect 42533 45985 42567 46019
rect 47041 45985 47075 46019
rect 2053 45917 2087 45951
rect 5089 45917 5123 45951
rect 11989 45917 12023 45951
rect 14105 45917 14139 45951
rect 19809 45917 19843 45951
rect 24593 45917 24627 45951
rect 25237 45917 25271 45951
rect 38209 45917 38243 45951
rect 43361 45917 43395 45951
rect 44281 45917 44315 45951
rect 45661 45917 45695 45951
rect 46305 45917 46339 45951
rect 21005 45849 21039 45883
rect 25421 45849 25455 45883
rect 41245 45849 41279 45883
rect 44373 45849 44407 45883
rect 46489 45849 46523 45883
rect 43453 45781 43487 45815
rect 45753 45781 45787 45815
rect 11897 45577 11931 45611
rect 21005 45577 21039 45611
rect 33057 45577 33091 45611
rect 40417 45577 40451 45611
rect 41429 45577 41463 45611
rect 42901 45509 42935 45543
rect 47961 45509 47995 45543
rect 1777 45441 1811 45475
rect 11805 45441 11839 45475
rect 20913 45441 20947 45475
rect 25513 45441 25547 45475
rect 32965 45441 32999 45475
rect 40325 45441 40359 45475
rect 41337 45441 41371 45475
rect 42717 45441 42751 45475
rect 48145 45441 48179 45475
rect 1961 45373 1995 45407
rect 2789 45373 2823 45407
rect 43177 45373 43211 45407
rect 45017 45373 45051 45407
rect 45201 45373 45235 45407
rect 45569 45373 45603 45407
rect 2329 45033 2363 45067
rect 25421 45033 25455 45067
rect 43269 45033 43303 45067
rect 44097 45033 44131 45067
rect 45201 45033 45235 45067
rect 45753 45033 45787 45067
rect 46305 44897 46339 44931
rect 48145 44897 48179 44931
rect 2237 44829 2271 44863
rect 25329 44829 25363 44863
rect 43177 44829 43211 44863
rect 45661 44829 45695 44863
rect 46489 44761 46523 44795
rect 46305 44489 46339 44523
rect 47685 44489 47719 44523
rect 45109 44353 45143 44387
rect 45753 44353 45787 44387
rect 46213 44353 46247 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 38669 44285 38703 44319
rect 38853 44285 38887 44319
rect 40049 44285 40083 44319
rect 46949 44149 46983 44183
rect 38853 43945 38887 43979
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 26985 43741 27019 43775
rect 38761 43741 38795 43775
rect 45845 43741 45879 43775
rect 46305 43741 46339 43775
rect 27077 43605 27111 43639
rect 1409 43265 1443 43299
rect 47041 43265 47075 43299
rect 1685 43197 1719 43231
rect 47777 43061 47811 43095
rect 46305 42721 46339 42755
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 46949 42313 46983 42347
rect 46857 42177 46891 42211
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 47685 41973 47719 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46489 41633 46523 41667
rect 46305 41565 46339 41599
rect 48145 41565 48179 41599
rect 1593 41497 1627 41531
rect 2145 41225 2179 41259
rect 2053 41089 2087 41123
rect 47961 41089 47995 41123
rect 48053 40885 48087 40919
rect 47685 40681 47719 40715
rect 1869 40409 1903 40443
rect 1961 40341 1995 40375
rect 46765 40001 46799 40035
rect 46857 39797 46891 39831
rect 47777 39797 47811 39831
rect 24961 39457 24995 39491
rect 46305 39457 46339 39491
rect 46489 39457 46523 39491
rect 48145 39457 48179 39491
rect 22845 39389 22879 39423
rect 24869 39321 24903 39355
rect 22661 39253 22695 39287
rect 24409 39253 24443 39287
rect 24777 39253 24811 39287
rect 25513 39253 25547 39287
rect 24593 39049 24627 39083
rect 19809 38981 19843 39015
rect 22109 38981 22143 39015
rect 38761 38981 38795 39015
rect 19993 38913 20027 38947
rect 24225 38913 24259 38947
rect 39497 38913 39531 38947
rect 47869 38913 47903 38947
rect 21833 38845 21867 38879
rect 23581 38845 23615 38879
rect 24133 38845 24167 38879
rect 39957 38845 39991 38879
rect 48053 38777 48087 38811
rect 20177 38709 20211 38743
rect 38853 38709 38887 38743
rect 21557 38505 21591 38539
rect 23489 38437 23523 38471
rect 40693 38369 40727 38403
rect 19257 38301 19291 38335
rect 19441 38301 19475 38335
rect 20729 38301 20763 38335
rect 21465 38301 21499 38335
rect 23305 38301 23339 38335
rect 24409 38301 24443 38335
rect 38669 38301 38703 38335
rect 39865 38301 39899 38335
rect 46305 38301 46339 38335
rect 39221 38233 39255 38267
rect 46489 38233 46523 38267
rect 48145 38233 48179 38267
rect 19349 38165 19383 38199
rect 20821 38165 20855 38199
rect 24501 38165 24535 38199
rect 46857 37961 46891 37995
rect 19809 37893 19843 37927
rect 27077 37893 27111 37927
rect 39405 37893 39439 37927
rect 40233 37893 40267 37927
rect 17969 37825 18003 37859
rect 22477 37825 22511 37859
rect 24685 37825 24719 37859
rect 26985 37825 27019 37859
rect 27629 37825 27663 37859
rect 29377 37825 29411 37859
rect 38485 37825 38519 37859
rect 38761 37825 38795 37859
rect 46765 37825 46799 37859
rect 47777 37825 47811 37859
rect 19533 37757 19567 37791
rect 22753 37757 22787 37791
rect 24961 37757 24995 37791
rect 18153 37621 18187 37655
rect 21281 37621 21315 37655
rect 24225 37621 24259 37655
rect 26433 37621 26467 37655
rect 27721 37621 27755 37655
rect 29469 37621 29503 37655
rect 18613 37417 18647 37451
rect 21649 37417 21683 37451
rect 23397 37417 23431 37451
rect 24409 37417 24443 37451
rect 21189 37281 21223 37315
rect 21281 37281 21315 37315
rect 23213 37281 23247 37315
rect 24593 37281 24627 37315
rect 28641 37281 28675 37315
rect 29561 37281 29595 37315
rect 2053 37213 2087 37247
rect 18337 37213 18371 37247
rect 18429 37213 18463 37247
rect 18705 37213 18739 37247
rect 20913 37213 20947 37247
rect 21097 37213 21131 37247
rect 21465 37213 21499 37247
rect 23029 37213 23063 37247
rect 23397 37213 23431 37247
rect 24685 37213 24719 37247
rect 25973 37213 26007 37247
rect 28365 37213 28399 37247
rect 28457 37213 28491 37247
rect 28733 37213 28767 37247
rect 29745 37213 29779 37247
rect 24409 37145 24443 37179
rect 26249 37145 26283 37179
rect 29929 37145 29963 37179
rect 18153 37077 18187 37111
rect 23121 37077 23155 37111
rect 24869 37077 24903 37111
rect 27721 37077 27755 37111
rect 28181 37077 28215 37111
rect 26249 36873 26283 36907
rect 28457 36805 28491 36839
rect 1777 36737 1811 36771
rect 25605 36737 25639 36771
rect 26433 36737 26467 36771
rect 28181 36737 28215 36771
rect 30665 36737 30699 36771
rect 1961 36669 1995 36703
rect 2789 36669 2823 36703
rect 16681 36669 16715 36703
rect 16957 36669 16991 36703
rect 19533 36669 19567 36703
rect 19809 36669 19843 36703
rect 18429 36533 18463 36567
rect 21281 36533 21315 36567
rect 25697 36533 25731 36567
rect 29929 36533 29963 36567
rect 30757 36533 30791 36567
rect 2237 36329 2271 36363
rect 17693 36329 17727 36363
rect 18613 36329 18647 36363
rect 20729 36329 20763 36363
rect 21741 36329 21775 36363
rect 23765 36329 23799 36363
rect 25237 36329 25271 36363
rect 28365 36329 28399 36363
rect 17509 36193 17543 36227
rect 18245 36193 18279 36227
rect 23857 36193 23891 36227
rect 26433 36193 26467 36227
rect 28917 36193 28951 36227
rect 2145 36125 2179 36159
rect 17417 36125 17451 36159
rect 18429 36125 18463 36159
rect 18705 36125 18739 36159
rect 20913 36125 20947 36159
rect 21097 36125 21131 36159
rect 21189 36125 21223 36159
rect 21649 36125 21683 36159
rect 22385 36125 22419 36159
rect 23581 36125 23615 36159
rect 23673 36125 23707 36159
rect 25421 36125 25455 36159
rect 25605 36125 25639 36159
rect 25697 36125 25731 36159
rect 26157 36125 26191 36159
rect 26249 36125 26283 36159
rect 28490 36125 28524 36159
rect 29009 36125 29043 36159
rect 29745 36125 29779 36159
rect 26433 36057 26467 36091
rect 29561 36057 29595 36091
rect 22569 35989 22603 36023
rect 28549 35989 28583 36023
rect 29929 35989 29963 36023
rect 17601 35785 17635 35819
rect 22661 35785 22695 35819
rect 24225 35785 24259 35819
rect 22385 35717 22419 35751
rect 1593 35649 1627 35683
rect 17509 35649 17543 35683
rect 22109 35649 22143 35683
rect 22293 35649 22327 35683
rect 22477 35649 22511 35683
rect 24041 35649 24075 35683
rect 24409 35649 24443 35683
rect 24593 35649 24627 35683
rect 27445 35649 27479 35683
rect 28181 35649 28215 35683
rect 28917 35649 28951 35683
rect 29101 35649 29135 35683
rect 29837 35649 29871 35683
rect 48145 35649 48179 35683
rect 25697 35581 25731 35615
rect 26157 35581 26191 35615
rect 28457 35581 28491 35615
rect 30113 35581 30147 35615
rect 26065 35513 26099 35547
rect 27629 35513 27663 35547
rect 28365 35513 28399 35547
rect 1409 35445 1443 35479
rect 24501 35445 24535 35479
rect 28273 35445 28307 35479
rect 29009 35445 29043 35479
rect 31585 35445 31619 35479
rect 47961 35445 47995 35479
rect 21833 35241 21867 35275
rect 26341 35241 26375 35275
rect 27905 35241 27939 35275
rect 28825 35241 28859 35275
rect 31033 35241 31067 35275
rect 30021 35173 30055 35207
rect 17141 35105 17175 35139
rect 21649 35105 21683 35139
rect 25237 35105 25271 35139
rect 25605 35105 25639 35139
rect 26801 35105 26835 35139
rect 28641 35105 28675 35139
rect 30573 35105 30607 35139
rect 30665 35105 30699 35139
rect 16865 35037 16899 35071
rect 17049 35037 17083 35071
rect 19349 35037 19383 35071
rect 20545 35037 20579 35071
rect 21557 35037 21591 35071
rect 24409 35037 24443 35071
rect 25697 35037 25731 35071
rect 26525 35037 26559 35071
rect 26617 35037 26651 35071
rect 26893 35037 26927 35071
rect 27721 35037 27755 35071
rect 27997 35037 28031 35071
rect 28825 35037 28859 35071
rect 30297 35037 30331 35071
rect 30481 35037 30515 35071
rect 30849 35037 30883 35071
rect 48145 35037 48179 35071
rect 24593 34969 24627 35003
rect 28549 34969 28583 35003
rect 16681 34901 16715 34935
rect 19441 34901 19475 34935
rect 20729 34901 20763 34935
rect 24777 34901 24811 34935
rect 25881 34901 25915 34935
rect 27537 34901 27571 34935
rect 29009 34901 29043 34935
rect 47961 34901 47995 34935
rect 17233 34697 17267 34731
rect 24501 34697 24535 34731
rect 25053 34697 25087 34731
rect 27721 34697 27755 34731
rect 29377 34697 29411 34731
rect 23121 34629 23155 34663
rect 24041 34629 24075 34663
rect 25421 34629 25455 34663
rect 28825 34629 28859 34663
rect 15945 34561 15979 34595
rect 17417 34561 17451 34595
rect 17509 34561 17543 34595
rect 17785 34561 17819 34595
rect 20913 34561 20947 34595
rect 21097 34561 21131 34595
rect 22201 34561 22235 34595
rect 22385 34561 22419 34595
rect 22937 34561 22971 34595
rect 24317 34561 24351 34595
rect 25237 34561 25271 34595
rect 25329 34561 25363 34595
rect 25539 34561 25573 34595
rect 26249 34561 26283 34595
rect 27905 34561 27939 34595
rect 27997 34561 28031 34595
rect 28273 34561 28307 34595
rect 28733 34561 28767 34595
rect 28917 34561 28951 34595
rect 29561 34561 29595 34595
rect 29653 34561 29687 34595
rect 29837 34561 29871 34595
rect 29929 34561 29963 34595
rect 47777 34561 47811 34595
rect 16037 34493 16071 34527
rect 17693 34493 17727 34527
rect 18429 34493 18463 34527
rect 20177 34493 20211 34527
rect 21189 34493 21223 34527
rect 22477 34493 22511 34527
rect 23305 34493 23339 34527
rect 24133 34493 24167 34527
rect 25697 34493 25731 34527
rect 26433 34493 26467 34527
rect 28181 34493 28215 34527
rect 18692 34357 18726 34391
rect 20729 34357 20763 34391
rect 22017 34357 22051 34391
rect 24317 34357 24351 34391
rect 47593 34357 47627 34391
rect 19993 34153 20027 34187
rect 21465 34153 21499 34187
rect 22293 34153 22327 34187
rect 23673 34153 23707 34187
rect 25145 34153 25179 34187
rect 25329 34153 25363 34187
rect 29009 34153 29043 34187
rect 21649 34085 21683 34119
rect 15761 34017 15795 34051
rect 19625 34017 19659 34051
rect 22293 34017 22327 34051
rect 27261 34017 27295 34051
rect 47133 34017 47167 34051
rect 47685 34017 47719 34051
rect 1593 33949 1627 33983
rect 19257 33949 19291 33983
rect 19441 33949 19475 33983
rect 19533 33949 19567 33983
rect 19809 33949 19843 33983
rect 21097 33949 21131 33983
rect 21373 33949 21407 33983
rect 22109 33949 22143 33983
rect 22385 33949 22419 33983
rect 23581 33949 23615 33983
rect 25789 33949 25823 33983
rect 30481 33949 30515 33983
rect 30849 33949 30883 33983
rect 16037 33881 16071 33915
rect 24961 33881 24995 33915
rect 25177 33881 25211 33915
rect 27537 33881 27571 33915
rect 30665 33881 30699 33915
rect 30757 33881 30791 33915
rect 47225 33881 47259 33915
rect 1409 33813 1443 33847
rect 17509 33813 17543 33847
rect 22569 33813 22603 33847
rect 25973 33813 26007 33847
rect 31033 33813 31067 33847
rect 17509 33609 17543 33643
rect 20085 33609 20119 33643
rect 28825 33609 28859 33643
rect 48053 33609 48087 33643
rect 16957 33541 16991 33575
rect 22017 33541 22051 33575
rect 16681 33473 16715 33507
rect 17417 33473 17451 33507
rect 17601 33473 17635 33507
rect 19533 33473 19567 33507
rect 19901 33473 19935 33507
rect 21833 33473 21867 33507
rect 22753 33473 22787 33507
rect 24501 33473 24535 33507
rect 24961 33473 24995 33507
rect 28457 33473 28491 33507
rect 28641 33473 28675 33507
rect 30941 33473 30975 33507
rect 46857 33473 46891 33507
rect 47593 33473 47627 33507
rect 1409 33405 1443 33439
rect 1685 33405 1719 33439
rect 16957 33405 16991 33439
rect 30849 33405 30883 33439
rect 22937 33337 22971 33371
rect 31309 33337 31343 33371
rect 16773 33269 16807 33303
rect 19901 33269 19935 33303
rect 22201 33269 22235 33303
rect 24317 33269 24351 33303
rect 25053 33269 25087 33303
rect 28457 33269 28491 33303
rect 46949 33269 46983 33303
rect 47869 33269 47903 33303
rect 1961 33065 1995 33099
rect 17233 33065 17267 33099
rect 17601 33065 17635 33099
rect 21189 33065 21223 33099
rect 21649 33065 21683 33099
rect 24961 33065 24995 33099
rect 26249 33065 26283 33099
rect 28641 33065 28675 33099
rect 29653 33065 29687 33099
rect 19625 32997 19659 33031
rect 2329 32929 2363 32963
rect 17325 32929 17359 32963
rect 21373 32929 21407 32963
rect 25605 32929 25639 32963
rect 27445 32929 27479 32963
rect 27905 32929 27939 32963
rect 31125 32929 31159 32963
rect 1869 32861 1903 32895
rect 2973 32861 3007 32895
rect 17233 32861 17267 32895
rect 18521 32861 18555 32895
rect 19441 32861 19475 32895
rect 19717 32861 19751 32895
rect 21465 32861 21499 32895
rect 22109 32861 22143 32895
rect 24685 32861 24719 32895
rect 25329 32861 25363 32895
rect 26157 32861 26191 32895
rect 27537 32861 27571 32895
rect 29561 32861 29595 32895
rect 46305 32861 46339 32895
rect 18337 32793 18371 32827
rect 21189 32793 21223 32827
rect 28549 32793 28583 32827
rect 31401 32793 31435 32827
rect 46489 32793 46523 32827
rect 48145 32793 48179 32827
rect 2789 32725 2823 32759
rect 18705 32725 18739 32759
rect 19257 32725 19291 32759
rect 22201 32725 22235 32759
rect 25421 32725 25455 32759
rect 32873 32725 32907 32759
rect 21281 32521 21315 32555
rect 23029 32521 23063 32555
rect 27537 32521 27571 32555
rect 30573 32521 30607 32555
rect 31125 32521 31159 32555
rect 33701 32521 33735 32555
rect 46949 32521 46983 32555
rect 48053 32521 48087 32555
rect 2329 32453 2363 32487
rect 23857 32453 23891 32487
rect 25789 32453 25823 32487
rect 25989 32453 26023 32487
rect 27445 32453 27479 32487
rect 2145 32385 2179 32419
rect 16865 32385 16899 32419
rect 17785 32385 17819 32419
rect 19073 32385 19107 32419
rect 19349 32385 19383 32419
rect 20821 32385 20855 32419
rect 21097 32385 21131 32419
rect 22201 32385 22235 32419
rect 22937 32385 22971 32419
rect 23581 32385 23615 32419
rect 28181 32385 28215 32419
rect 28365 32385 28399 32419
rect 28825 32385 28859 32419
rect 29009 32385 29043 32419
rect 29929 32385 29963 32419
rect 30076 32385 30110 32419
rect 31309 32385 31343 32419
rect 31493 32385 31527 32419
rect 31585 32385 31619 32419
rect 32137 32385 32171 32419
rect 32321 32385 32355 32419
rect 32965 32385 32999 32419
rect 33609 32385 33643 32419
rect 46857 32385 46891 32419
rect 47961 32385 47995 32419
rect 3985 32317 4019 32351
rect 16957 32317 16991 32351
rect 18061 32317 18095 32351
rect 20913 32317 20947 32351
rect 22017 32317 22051 32351
rect 25329 32317 25363 32351
rect 30297 32317 30331 32351
rect 32505 32317 32539 32351
rect 26157 32249 26191 32283
rect 33057 32249 33091 32283
rect 1685 32181 1719 32215
rect 17233 32181 17267 32215
rect 19257 32181 19291 32215
rect 19625 32181 19659 32215
rect 21097 32181 21131 32215
rect 22385 32181 22419 32215
rect 25973 32181 26007 32215
rect 28825 32181 28859 32215
rect 30205 32181 30239 32215
rect 18245 31977 18279 32011
rect 26249 31977 26283 32011
rect 30389 31977 30423 32011
rect 47685 31977 47719 32011
rect 17601 31909 17635 31943
rect 21189 31909 21223 31943
rect 30757 31909 30791 31943
rect 34161 31909 34195 31943
rect 1409 31841 1443 31875
rect 1593 31841 1627 31875
rect 3893 31841 3927 31875
rect 15853 31841 15887 31875
rect 18337 31841 18371 31875
rect 19441 31841 19475 31875
rect 22477 31841 22511 31875
rect 23765 31841 23799 31875
rect 27169 31841 27203 31875
rect 28917 31841 28951 31875
rect 29653 31841 29687 31875
rect 32413 31841 32447 31875
rect 32689 31841 32723 31875
rect 3249 31773 3283 31807
rect 3801 31773 3835 31807
rect 7481 31773 7515 31807
rect 18521 31773 18555 31807
rect 22261 31773 22295 31807
rect 22385 31773 22419 31807
rect 23029 31773 23063 31807
rect 23673 31773 23707 31807
rect 23857 31773 23891 31807
rect 24961 31773 24995 31807
rect 29561 31773 29595 31807
rect 30389 31773 30423 31807
rect 30481 31773 30515 31807
rect 31309 31773 31343 31807
rect 31401 31773 31435 31807
rect 31539 31773 31573 31807
rect 31677 31773 31711 31807
rect 16129 31705 16163 31739
rect 18245 31705 18279 31739
rect 19717 31705 19751 31739
rect 27445 31705 27479 31739
rect 7573 31637 7607 31671
rect 18705 31637 18739 31671
rect 22017 31637 22051 31671
rect 23121 31637 23155 31671
rect 31769 31637 31803 31671
rect 17325 31433 17359 31467
rect 17877 31433 17911 31467
rect 19717 31433 19751 31467
rect 23581 31433 23615 31467
rect 28089 31433 28123 31467
rect 28917 31433 28951 31467
rect 33149 31433 33183 31467
rect 33793 31433 33827 31467
rect 2789 31365 2823 31399
rect 17049 31365 17083 31399
rect 20913 31365 20947 31399
rect 27813 31365 27847 31399
rect 15945 31297 15979 31331
rect 16129 31297 16163 31331
rect 16681 31297 16715 31331
rect 16801 31297 16835 31331
rect 16957 31297 16991 31331
rect 17146 31297 17180 31331
rect 17785 31297 17819 31331
rect 18981 31297 19015 31331
rect 19165 31297 19199 31331
rect 19533 31297 19567 31331
rect 24685 31297 24719 31331
rect 25513 31297 25547 31331
rect 27445 31297 27479 31331
rect 27538 31297 27572 31331
rect 27721 31297 27755 31331
rect 27951 31297 27985 31331
rect 28825 31297 28859 31331
rect 29009 31297 29043 31331
rect 31033 31297 31067 31331
rect 32413 31297 32447 31331
rect 32597 31297 32631 31331
rect 32689 31297 32723 31331
rect 32965 31297 32999 31331
rect 33701 31297 33735 31331
rect 2605 31229 2639 31263
rect 4445 31229 4479 31263
rect 16037 31229 16071 31263
rect 19257 31229 19291 31263
rect 19349 31229 19383 31263
rect 21833 31229 21867 31263
rect 22109 31229 22143 31263
rect 24777 31229 24811 31263
rect 25053 31229 25087 31263
rect 30757 31229 30791 31263
rect 32781 31229 32815 31263
rect 21097 31161 21131 31195
rect 6929 31093 6963 31127
rect 25697 31093 25731 31127
rect 21925 30889 21959 30923
rect 22477 30889 22511 30923
rect 24593 30889 24627 30923
rect 25329 30889 25363 30923
rect 25513 30889 25547 30923
rect 30205 30889 30239 30923
rect 30757 30889 30791 30923
rect 26249 30821 26283 30855
rect 26985 30821 27019 30855
rect 6561 30753 6595 30787
rect 6745 30753 6779 30787
rect 8217 30753 8251 30787
rect 28825 30753 28859 30787
rect 30941 30753 30975 30787
rect 32781 30753 32815 30787
rect 47133 30753 47167 30787
rect 21281 30685 21315 30719
rect 21429 30685 21463 30719
rect 21557 30685 21591 30719
rect 21746 30685 21780 30719
rect 22385 30685 22419 30719
rect 24409 30685 24443 30719
rect 26065 30685 26099 30719
rect 27997 30685 28031 30719
rect 28733 30685 28767 30719
rect 30021 30685 30055 30719
rect 30665 30685 30699 30719
rect 32413 30685 32447 30719
rect 32597 30685 32631 30719
rect 32689 30685 32723 30719
rect 32965 30685 32999 30719
rect 21649 30617 21683 30651
rect 25145 30617 25179 30651
rect 25345 30617 25379 30651
rect 26801 30617 26835 30651
rect 29837 30617 29871 30651
rect 46857 30617 46891 30651
rect 46949 30617 46983 30651
rect 28181 30549 28215 30583
rect 30941 30549 30975 30583
rect 33149 30549 33183 30583
rect 29653 30345 29687 30379
rect 30573 30345 30607 30379
rect 27537 30277 27571 30311
rect 33149 30277 33183 30311
rect 16957 30209 16991 30243
rect 19257 30209 19291 30243
rect 19441 30209 19475 30243
rect 19625 30209 19659 30243
rect 19809 30209 19843 30243
rect 24133 30209 24167 30243
rect 24869 30209 24903 30243
rect 25789 30209 25823 30243
rect 25973 30209 26007 30243
rect 26065 30209 26099 30243
rect 28365 30209 28399 30243
rect 28457 30209 28491 30243
rect 28733 30209 28767 30243
rect 29469 30209 29503 30243
rect 30205 30209 30239 30243
rect 31033 30209 31067 30243
rect 17233 30141 17267 30175
rect 19533 30141 19567 30175
rect 25605 30141 25639 30175
rect 28641 30141 28675 30175
rect 30297 30141 30331 30175
rect 31309 30141 31343 30175
rect 32873 30141 32907 30175
rect 19993 30073 20027 30107
rect 24317 30073 24351 30107
rect 31585 30073 31619 30107
rect 18705 30005 18739 30039
rect 25053 30005 25087 30039
rect 27629 30005 27663 30039
rect 28181 30005 28215 30039
rect 30389 30005 30423 30039
rect 31401 30005 31435 30039
rect 34621 30005 34655 30039
rect 18061 29801 18095 29835
rect 19717 29801 19751 29835
rect 20545 29801 20579 29835
rect 28825 29801 28859 29835
rect 29929 29801 29963 29835
rect 33793 29801 33827 29835
rect 19533 29665 19567 29699
rect 24777 29665 24811 29699
rect 30481 29665 30515 29699
rect 17969 29597 18003 29631
rect 19441 29597 19475 29631
rect 20453 29597 20487 29631
rect 20729 29597 20763 29631
rect 24501 29597 24535 29631
rect 25789 29597 25823 29631
rect 27077 29597 27111 29631
rect 29745 29597 29779 29631
rect 30021 29597 30055 29631
rect 33701 29597 33735 29631
rect 48145 29597 48179 29631
rect 27353 29529 27387 29563
rect 29561 29529 29595 29563
rect 30757 29529 30791 29563
rect 21005 29461 21039 29495
rect 25973 29461 26007 29495
rect 32229 29461 32263 29495
rect 47961 29461 47995 29495
rect 19533 29257 19567 29291
rect 25421 29257 25455 29291
rect 27445 29257 27479 29291
rect 30205 29257 30239 29291
rect 32229 29257 32263 29291
rect 18981 29189 19015 29223
rect 29009 29189 29043 29223
rect 16681 29121 16715 29155
rect 18889 29121 18923 29155
rect 19717 29121 19751 29155
rect 19993 29121 20027 29155
rect 20545 29121 20579 29155
rect 20729 29121 20763 29155
rect 20821 29121 20855 29155
rect 21097 29121 21131 29155
rect 22661 29121 22695 29155
rect 24869 29121 24903 29155
rect 25881 29121 25915 29155
rect 27629 29121 27663 29155
rect 27721 29121 27755 29155
rect 27997 29121 28031 29155
rect 28825 29121 28859 29155
rect 30389 29121 30423 29155
rect 30481 29121 30515 29155
rect 30665 29121 30699 29155
rect 30757 29121 30791 29155
rect 32137 29121 32171 29155
rect 18429 29053 18463 29087
rect 20913 29053 20947 29087
rect 22937 29053 22971 29087
rect 25145 29053 25179 29087
rect 28641 29053 28675 29087
rect 19901 28985 19935 29019
rect 26065 28985 26099 29019
rect 27905 28985 27939 29019
rect 16944 28917 16978 28951
rect 21281 28917 21315 28951
rect 24409 28917 24443 28951
rect 25237 28917 25271 28951
rect 19993 28713 20027 28747
rect 23305 28713 23339 28747
rect 27077 28713 27111 28747
rect 28365 28713 28399 28747
rect 30113 28713 30147 28747
rect 25421 28645 25455 28679
rect 19901 28577 19935 28611
rect 21189 28577 21223 28611
rect 22845 28577 22879 28611
rect 17693 28509 17727 28543
rect 19809 28509 19843 28543
rect 21465 28509 21499 28543
rect 22569 28509 22603 28543
rect 22753 28509 22787 28543
rect 22937 28509 22971 28543
rect 23121 28509 23155 28543
rect 25237 28509 25271 28543
rect 26893 28509 26927 28543
rect 28273 28509 28307 28543
rect 30389 28509 30423 28543
rect 18337 28441 18371 28475
rect 18521 28441 18555 28475
rect 30113 28441 30147 28475
rect 30297 28441 30331 28475
rect 17785 28373 17819 28407
rect 18705 28373 18739 28407
rect 20177 28373 20211 28407
rect 18613 28169 18647 28203
rect 22201 28169 22235 28203
rect 25697 28169 25731 28203
rect 19809 28101 19843 28135
rect 20637 28101 20671 28135
rect 20821 28101 20855 28135
rect 23765 28101 23799 28135
rect 29377 28101 29411 28135
rect 29561 28101 29595 28135
rect 16865 28033 16899 28067
rect 19533 28033 19567 28067
rect 19626 28033 19660 28067
rect 19909 28033 19943 28067
rect 20039 28033 20073 28067
rect 21833 28033 21867 28067
rect 22845 28033 22879 28067
rect 23581 28033 23615 28067
rect 24685 28033 24719 28067
rect 25513 28033 25547 28067
rect 30021 28033 30055 28067
rect 30205 28033 30239 28067
rect 30297 28033 30331 28067
rect 46857 28033 46891 28067
rect 17141 27965 17175 27999
rect 21925 27965 21959 27999
rect 23121 27965 23155 27999
rect 24777 27965 24811 27999
rect 20177 27897 20211 27931
rect 20913 27829 20947 27863
rect 22017 27829 22051 27863
rect 22661 27829 22695 27863
rect 23029 27829 23063 27863
rect 23949 27829 23983 27863
rect 24777 27829 24811 27863
rect 25053 27829 25087 27863
rect 30021 27829 30055 27863
rect 46949 27829 46983 27863
rect 47777 27829 47811 27863
rect 21005 27625 21039 27659
rect 21465 27625 21499 27659
rect 23765 27625 23799 27659
rect 24777 27625 24811 27659
rect 30941 27625 30975 27659
rect 26249 27557 26283 27591
rect 31125 27557 31159 27591
rect 31585 27557 31619 27591
rect 16129 27489 16163 27523
rect 17049 27489 17083 27523
rect 21189 27489 21223 27523
rect 28457 27489 28491 27523
rect 30849 27489 30883 27523
rect 46305 27489 46339 27523
rect 46489 27489 46523 27523
rect 48145 27489 48179 27523
rect 14289 27421 14323 27455
rect 16589 27421 16623 27455
rect 19257 27421 19291 27455
rect 19441 27421 19475 27455
rect 20269 27421 20303 27455
rect 20361 27421 20395 27455
rect 21281 27421 21315 27455
rect 22753 27421 22787 27455
rect 22937 27421 22971 27455
rect 23581 27421 23615 27455
rect 25053 27421 25087 27455
rect 25145 27421 25179 27455
rect 25237 27421 25271 27455
rect 25421 27421 25455 27455
rect 25973 27421 26007 27455
rect 26065 27421 26099 27455
rect 27077 27421 27111 27455
rect 27353 27421 27387 27455
rect 28181 27421 28215 27455
rect 29837 27421 29871 27455
rect 30021 27421 30055 27455
rect 30205 27421 30239 27455
rect 30941 27421 30975 27455
rect 31769 27421 31803 27455
rect 31953 27421 31987 27455
rect 32045 27421 32079 27455
rect 14473 27353 14507 27387
rect 16773 27353 16807 27387
rect 21005 27353 21039 27387
rect 23397 27353 23431 27387
rect 30665 27353 30699 27387
rect 19349 27285 19383 27319
rect 20545 27285 20579 27319
rect 22845 27285 22879 27319
rect 26893 27285 26927 27319
rect 27261 27285 27295 27319
rect 27813 27285 27847 27319
rect 28273 27285 28307 27319
rect 10977 27081 11011 27115
rect 13277 27081 13311 27115
rect 14381 27081 14415 27115
rect 15669 27081 15703 27115
rect 19441 27081 19475 27115
rect 27721 27081 27755 27115
rect 28641 27081 28675 27115
rect 30941 27081 30975 27115
rect 31493 27081 31527 27115
rect 11805 27013 11839 27047
rect 22201 27013 22235 27047
rect 25170 27013 25204 27047
rect 30665 27013 30699 27047
rect 10609 26945 10643 26979
rect 14289 26945 14323 26979
rect 14933 26945 14967 26979
rect 15577 26945 15611 26979
rect 19349 26945 19383 26979
rect 19533 26945 19567 26979
rect 20453 26945 20487 26979
rect 20637 26945 20671 26979
rect 20821 26945 20855 26979
rect 21833 26945 21867 26979
rect 21926 26945 21960 26979
rect 22109 26945 22143 26979
rect 22339 26945 22373 26979
rect 24685 26945 24719 26979
rect 25053 26945 25087 26979
rect 25987 26935 26021 26969
rect 26138 26945 26172 26979
rect 26234 26945 26268 26979
rect 26341 26945 26375 26979
rect 27537 26945 27571 26979
rect 28457 26945 28491 26979
rect 29653 26945 29687 26979
rect 29837 26945 29871 26979
rect 29929 26945 29963 26979
rect 30389 26945 30423 26979
rect 30573 26945 30607 26979
rect 30757 26945 30791 26979
rect 31401 26945 31435 26979
rect 31585 26945 31619 26979
rect 32321 26945 32355 26979
rect 10701 26877 10735 26911
rect 11529 26877 11563 26911
rect 24961 26877 24995 26911
rect 32229 26877 32263 26911
rect 20545 26809 20579 26843
rect 25329 26809 25363 26843
rect 32689 26809 32723 26843
rect 15025 26741 15059 26775
rect 20177 26741 20211 26775
rect 20729 26741 20763 26775
rect 22477 26741 22511 26775
rect 25789 26741 25823 26775
rect 29469 26741 29503 26775
rect 11253 26537 11287 26571
rect 20361 26537 20395 26571
rect 21373 26537 21407 26571
rect 27426 26537 27460 26571
rect 28917 26537 28951 26571
rect 32781 26537 32815 26571
rect 25237 26469 25271 26503
rect 26065 26469 26099 26503
rect 15209 26401 15243 26435
rect 15485 26401 15519 26435
rect 19993 26401 20027 26435
rect 21189 26401 21223 26435
rect 31033 26401 31067 26435
rect 31309 26401 31343 26435
rect 11161 26333 11195 26367
rect 11345 26333 11379 26367
rect 13277 26333 13311 26367
rect 15025 26333 15059 26367
rect 20177 26333 20211 26367
rect 21097 26333 21131 26367
rect 24685 26333 24719 26367
rect 24869 26333 24903 26367
rect 25053 26333 25087 26367
rect 27169 26333 27203 26367
rect 29561 26333 29595 26367
rect 29745 26333 29779 26367
rect 29837 26333 29871 26367
rect 29929 26333 29963 26367
rect 47685 26333 47719 26367
rect 13369 26265 13403 26299
rect 24961 26265 24995 26299
rect 25697 26265 25731 26299
rect 25881 26265 25915 26299
rect 30113 26197 30147 26231
rect 10793 25993 10827 26027
rect 12081 25993 12115 26027
rect 23581 25993 23615 26027
rect 24133 25993 24167 26027
rect 27537 25993 27571 26027
rect 29101 25993 29135 26027
rect 31493 25993 31527 26027
rect 22109 25925 22143 25959
rect 28549 25925 28583 25959
rect 30021 25925 30055 25959
rect 10701 25857 10735 25891
rect 11989 25857 12023 25891
rect 12817 25857 12851 25891
rect 13829 25857 13863 25891
rect 15025 25857 15059 25891
rect 16681 25857 16715 25891
rect 16865 25857 16899 25891
rect 17693 25857 17727 25891
rect 18429 25857 18463 25891
rect 18613 25857 18647 25891
rect 21833 25857 21867 25891
rect 24041 25857 24075 25891
rect 24777 25857 24811 25891
rect 25421 25857 25455 25891
rect 27261 25857 27295 25891
rect 27629 25857 27663 25891
rect 28365 25857 28399 25891
rect 29009 25857 29043 25891
rect 29837 25857 29871 25891
rect 30205 25857 30239 25891
rect 30849 25857 30883 25891
rect 31401 25857 31435 25891
rect 46305 25857 46339 25891
rect 13093 25789 13127 25823
rect 13737 25789 13771 25823
rect 27077 25789 27111 25823
rect 13001 25721 13035 25755
rect 12633 25653 12667 25687
rect 14105 25653 14139 25687
rect 15117 25653 15151 25687
rect 17049 25653 17083 25687
rect 17877 25653 17911 25687
rect 18429 25653 18463 25687
rect 24869 25653 24903 25687
rect 25513 25653 25547 25687
rect 30665 25653 30699 25687
rect 46397 25653 46431 25687
rect 47777 25653 47811 25687
rect 11805 25449 11839 25483
rect 16773 25449 16807 25483
rect 17785 25449 17819 25483
rect 18245 25449 18279 25483
rect 22937 25449 22971 25483
rect 24672 25449 24706 25483
rect 31401 25449 31435 25483
rect 17233 25381 17267 25415
rect 26157 25381 26191 25415
rect 9413 25313 9447 25347
rect 14473 25313 14507 25347
rect 24409 25313 24443 25347
rect 29653 25313 29687 25347
rect 29929 25313 29963 25347
rect 46489 25313 46523 25347
rect 48145 25313 48179 25347
rect 8953 25245 8987 25279
rect 11437 25245 11471 25279
rect 12725 25245 12759 25279
rect 14197 25245 14231 25279
rect 16497 25245 16531 25279
rect 16589 25245 16623 25279
rect 17601 25245 17635 25279
rect 18521 25245 18555 25279
rect 22845 25245 22879 25279
rect 46305 25245 46339 25279
rect 1869 25177 1903 25211
rect 9137 25177 9171 25211
rect 11253 25177 11287 25211
rect 12449 25177 12483 25211
rect 18245 25177 18279 25211
rect 1961 25109 1995 25143
rect 11529 25109 11563 25143
rect 11621 25109 11655 25143
rect 12633 25109 12667 25143
rect 12817 25109 12851 25143
rect 13001 25109 13035 25143
rect 15945 25109 15979 25143
rect 17417 25109 17451 25143
rect 17509 25109 17543 25143
rect 18429 25109 18463 25143
rect 8861 24905 8895 24939
rect 11621 24905 11655 24939
rect 14933 24905 14967 24939
rect 17049 24905 17083 24939
rect 19809 24905 19843 24939
rect 23121 24905 23155 24939
rect 26157 24905 26191 24939
rect 12817 24837 12851 24871
rect 16957 24837 16991 24871
rect 18337 24837 18371 24871
rect 39589 24837 39623 24871
rect 8769 24769 8803 24803
rect 9689 24769 9723 24803
rect 9873 24769 9907 24803
rect 10517 24769 10551 24803
rect 11529 24769 11563 24803
rect 11897 24769 11931 24803
rect 12541 24769 12575 24803
rect 14749 24769 14783 24803
rect 15945 24769 15979 24803
rect 16681 24769 16715 24803
rect 16865 24769 16899 24803
rect 18061 24769 18095 24803
rect 20269 24769 20303 24803
rect 20913 24769 20947 24803
rect 22201 24769 22235 24803
rect 22937 24769 22971 24803
rect 27629 24769 27663 24803
rect 28273 24769 28307 24803
rect 30665 24769 30699 24803
rect 30757 24769 30791 24803
rect 38761 24769 38795 24803
rect 38853 24769 38887 24803
rect 45201 24769 45235 24803
rect 47593 24769 47627 24803
rect 11713 24701 11747 24735
rect 14289 24701 14323 24735
rect 20361 24701 20395 24735
rect 24409 24701 24443 24735
rect 24685 24701 24719 24735
rect 39405 24701 39439 24735
rect 40969 24701 41003 24735
rect 45385 24701 45419 24735
rect 46857 24701 46891 24735
rect 11897 24633 11931 24667
rect 9689 24565 9723 24599
rect 10333 24565 10367 24599
rect 16037 24565 16071 24599
rect 17233 24565 17267 24599
rect 21005 24565 21039 24599
rect 22385 24565 22419 24599
rect 27721 24565 27755 24599
rect 28365 24565 28399 24599
rect 47685 24565 47719 24599
rect 13461 24361 13495 24395
rect 14197 24361 14231 24395
rect 10333 24225 10367 24259
rect 10609 24225 10643 24259
rect 16589 24225 16623 24259
rect 17141 24225 17175 24259
rect 20453 24225 20487 24259
rect 22109 24225 22143 24259
rect 27353 24225 27387 24259
rect 29009 24225 29043 24259
rect 46305 24225 46339 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 12541 24157 12575 24191
rect 13369 24157 13403 24191
rect 13553 24157 13587 24191
rect 14105 24157 14139 24191
rect 17601 24157 17635 24191
rect 17969 24157 18003 24191
rect 18061 24157 18095 24191
rect 19533 24157 19567 24191
rect 20269 24157 20303 24191
rect 22661 24157 22695 24191
rect 24409 24157 24443 24191
rect 27169 24157 27203 24191
rect 43085 24157 43119 24191
rect 43269 24157 43303 24191
rect 45845 24157 45879 24191
rect 12633 24089 12667 24123
rect 16865 24089 16899 24123
rect 16957 24089 16991 24123
rect 12081 24021 12115 24055
rect 16773 24021 16807 24055
rect 17877 24021 17911 24055
rect 19625 24021 19659 24055
rect 22753 24021 22787 24055
rect 24501 24021 24535 24055
rect 43177 24021 43211 24055
rect 45661 24021 45695 24055
rect 26341 23817 26375 23851
rect 40601 23817 40635 23851
rect 41337 23817 41371 23851
rect 47685 23817 47719 23851
rect 16681 23749 16715 23783
rect 18337 23749 18371 23783
rect 20729 23749 20763 23783
rect 26065 23749 26099 23783
rect 27721 23749 27755 23783
rect 42717 23749 42751 23783
rect 1869 23681 1903 23715
rect 8401 23681 8435 23715
rect 14565 23681 14599 23715
rect 16865 23681 16899 23715
rect 17049 23681 17083 23715
rect 17141 23681 17175 23715
rect 20361 23681 20395 23715
rect 21925 23681 21959 23715
rect 23029 23681 23063 23715
rect 25329 23681 25363 23715
rect 37749 23681 37783 23715
rect 39221 23681 39255 23715
rect 40233 23681 40267 23715
rect 41153 23681 41187 23715
rect 42441 23681 42475 23715
rect 43361 23681 43395 23715
rect 43545 23681 43579 23715
rect 47593 23681 47627 23715
rect 8585 23613 8619 23647
rect 9781 23613 9815 23647
rect 18061 23613 18095 23647
rect 19809 23613 19843 23647
rect 22477 23613 22511 23647
rect 27537 23613 27571 23647
rect 27997 23613 28031 23647
rect 39129 23613 39163 23647
rect 39589 23613 39623 23647
rect 40141 23613 40175 23647
rect 45201 23613 45235 23647
rect 45385 23613 45419 23647
rect 46673 23613 46707 23647
rect 14749 23545 14783 23579
rect 1961 23477 1995 23511
rect 23121 23477 23155 23511
rect 25421 23477 25455 23511
rect 38025 23477 38059 23511
rect 43453 23477 43487 23511
rect 9045 23273 9079 23307
rect 43453 23273 43487 23307
rect 47961 23273 47995 23307
rect 17877 23205 17911 23239
rect 20085 23205 20119 23239
rect 42901 23205 42935 23239
rect 16497 23137 16531 23171
rect 16773 23137 16807 23171
rect 23489 23137 23523 23171
rect 25237 23137 25271 23171
rect 25421 23137 25455 23171
rect 27905 23137 27939 23171
rect 28181 23137 28215 23171
rect 38393 23137 38427 23171
rect 40049 23137 40083 23171
rect 45385 23137 45419 23171
rect 8953 23069 8987 23103
rect 10701 23069 10735 23103
rect 14749 23069 14783 23103
rect 15393 23069 15427 23103
rect 16405 23069 16439 23103
rect 17693 23069 17727 23103
rect 19901 23069 19935 23103
rect 20637 23069 20671 23103
rect 21741 23069 21775 23103
rect 27813 23069 27847 23103
rect 36829 23069 36863 23103
rect 37749 23069 37783 23103
rect 43026 23069 43060 23103
rect 43545 23069 43579 23103
rect 44005 23069 44039 23103
rect 44189 23069 44223 23103
rect 47685 23069 47719 23103
rect 22017 23001 22051 23035
rect 27077 23001 27111 23035
rect 40233 23001 40267 23035
rect 41889 23001 41923 23035
rect 45569 23001 45603 23035
rect 47225 23001 47259 23035
rect 10885 22933 10919 22967
rect 14841 22933 14875 22967
rect 15485 22933 15519 22967
rect 20821 22933 20855 22967
rect 37013 22933 37047 22967
rect 43085 22933 43119 22967
rect 44097 22933 44131 22967
rect 48145 22933 48179 22967
rect 23765 22729 23799 22763
rect 26249 22729 26283 22763
rect 29285 22729 29319 22763
rect 39497 22729 39531 22763
rect 40785 22729 40819 22763
rect 42809 22729 42843 22763
rect 44281 22729 44315 22763
rect 45661 22729 45695 22763
rect 13553 22661 13587 22695
rect 14657 22661 14691 22695
rect 22099 22661 22133 22695
rect 22845 22661 22879 22695
rect 27813 22661 27847 22695
rect 35909 22661 35943 22695
rect 37565 22661 37599 22695
rect 39221 22661 39255 22695
rect 23075 22627 23109 22661
rect 8493 22593 8527 22627
rect 11529 22593 11563 22627
rect 14381 22593 14415 22627
rect 22293 22593 22327 22627
rect 22385 22593 22419 22627
rect 23673 22593 23707 22627
rect 23857 22593 23891 22627
rect 34713 22593 34747 22627
rect 35817 22593 35851 22627
rect 36461 22593 36495 22627
rect 39865 22593 39899 22627
rect 40969 22593 41003 22627
rect 42993 22593 43027 22627
rect 43177 22593 43211 22627
rect 44465 22593 44499 22627
rect 45109 22593 45143 22627
rect 45569 22593 45603 22627
rect 47593 22593 47627 22627
rect 8677 22525 8711 22559
rect 8953 22525 8987 22559
rect 11805 22525 11839 22559
rect 16129 22525 16163 22559
rect 17601 22525 17635 22559
rect 17785 22525 17819 22559
rect 19073 22525 19107 22559
rect 24501 22525 24535 22559
rect 24777 22525 24811 22559
rect 27537 22525 27571 22559
rect 37381 22525 37415 22559
rect 40325 22525 40359 22559
rect 43269 22525 43303 22559
rect 46213 22525 46247 22559
rect 46489 22525 46523 22559
rect 47869 22525 47903 22559
rect 22109 22457 22143 22491
rect 23213 22457 23247 22491
rect 48145 22457 48179 22491
rect 23029 22389 23063 22423
rect 34529 22389 34563 22423
rect 36645 22389 36679 22423
rect 39957 22389 39991 22423
rect 44925 22389 44959 22423
rect 47685 22389 47719 22423
rect 9045 22185 9079 22219
rect 17785 22185 17819 22219
rect 21833 22185 21867 22219
rect 22385 22185 22419 22219
rect 24501 22185 24535 22219
rect 27261 22185 27295 22219
rect 34713 22185 34747 22219
rect 34897 22185 34931 22219
rect 35449 22185 35483 22219
rect 43085 22117 43119 22151
rect 10701 22049 10735 22083
rect 10977 22049 11011 22083
rect 12081 22049 12115 22083
rect 14110 22049 14144 22083
rect 19533 22049 19567 22083
rect 19809 22049 19843 22083
rect 25605 22049 25639 22083
rect 34069 22049 34103 22083
rect 46029 22049 46063 22083
rect 8953 21981 8987 22015
rect 10609 21981 10643 22015
rect 11989 21981 12023 22015
rect 12633 21981 12667 22015
rect 13277 21981 13311 22015
rect 16405 21981 16439 22015
rect 17693 21981 17727 22015
rect 19441 21981 19475 22015
rect 20453 21981 20487 22015
rect 21005 21981 21039 22015
rect 21649 21981 21683 22015
rect 22661 21981 22695 22015
rect 23121 21981 23155 22015
rect 23489 21981 23523 22015
rect 24501 21981 24535 22015
rect 25513 21981 25547 22015
rect 27169 21981 27203 22015
rect 28733 21981 28767 22015
rect 29561 21981 29595 22015
rect 30297 21981 30331 22015
rect 32229 21981 32263 22015
rect 35173 21981 35207 22015
rect 36277 21981 36311 22015
rect 37565 21981 37599 22015
rect 39129 21981 39163 22015
rect 39865 21981 39899 22015
rect 40049 21981 40083 22015
rect 45201 21981 45235 22015
rect 45385 21981 45419 22015
rect 45845 21981 45879 22015
rect 12725 21913 12759 21947
rect 14289 21913 14323 21947
rect 15945 21913 15979 21947
rect 22385 21913 22419 21947
rect 32413 21913 32447 21947
rect 36921 21913 36955 21947
rect 40233 21913 40267 21947
rect 42717 21913 42751 21947
rect 47685 21913 47719 21947
rect 13461 21845 13495 21879
rect 16589 21845 16623 21879
rect 20453 21845 20487 21879
rect 21097 21845 21131 21879
rect 22569 21845 22603 21879
rect 23305 21845 23339 21879
rect 23397 21845 23431 21879
rect 23673 21845 23707 21879
rect 28825 21845 28859 21879
rect 29745 21845 29779 21879
rect 30389 21845 30423 21879
rect 43177 21845 43211 21879
rect 45385 21845 45419 21879
rect 11713 21641 11747 21675
rect 24409 21641 24443 21675
rect 28365 21641 28399 21675
rect 42717 21641 42751 21675
rect 45569 21641 45603 21675
rect 47777 21641 47811 21675
rect 47961 21641 47995 21675
rect 19717 21573 19751 21607
rect 23857 21573 23891 21607
rect 28181 21573 28215 21607
rect 33517 21573 33551 21607
rect 34621 21573 34655 21607
rect 34713 21573 34747 21607
rect 43729 21573 43763 21607
rect 46673 21573 46707 21607
rect 46857 21573 46891 21607
rect 10793 21505 10827 21539
rect 10977 21505 11011 21539
rect 11529 21505 11563 21539
rect 12265 21505 12299 21539
rect 16865 21505 16899 21539
rect 19441 21505 19475 21539
rect 21833 21505 21867 21539
rect 22569 21505 22603 21539
rect 23581 21505 23615 21539
rect 23673 21505 23707 21539
rect 24317 21505 24351 21539
rect 24501 21505 24535 21539
rect 25421 21505 25455 21539
rect 26985 21505 27019 21539
rect 27997 21505 28031 21539
rect 28089 21505 28123 21539
rect 28825 21505 28859 21539
rect 29009 21505 29043 21539
rect 29469 21505 29503 21539
rect 32229 21505 32263 21539
rect 36369 21505 36403 21539
rect 37749 21505 37783 21539
rect 41705 21505 41739 21539
rect 41889 21505 41923 21539
rect 42901 21505 42935 21539
rect 43637 21505 43671 21539
rect 43821 21505 43855 21539
rect 44741 21505 44775 21539
rect 46213 21505 46247 21539
rect 47593 21505 47627 21539
rect 47869 21505 47903 21539
rect 13553 21437 13587 21471
rect 13737 21437 13771 21471
rect 14013 21437 14047 21471
rect 29745 21437 29779 21471
rect 31217 21437 31251 21471
rect 32781 21437 32815 21471
rect 33425 21437 33459 21471
rect 35633 21437 35667 21471
rect 38301 21437 38335 21471
rect 41797 21437 41831 21471
rect 43177 21437 43211 21471
rect 45017 21437 45051 21471
rect 47041 21437 47075 21471
rect 17049 21369 17083 21403
rect 27813 21369 27847 21403
rect 33977 21369 34011 21403
rect 48145 21369 48179 21403
rect 10793 21301 10827 21335
rect 12357 21301 12391 21335
rect 21189 21301 21223 21335
rect 21833 21301 21867 21335
rect 22661 21301 22695 21335
rect 25513 21301 25547 21335
rect 27077 21301 27111 21335
rect 28825 21301 28859 21335
rect 36645 21301 36679 21335
rect 43085 21301 43119 21335
rect 46029 21301 46063 21335
rect 12173 21097 12207 21131
rect 12633 21097 12667 21131
rect 14933 21097 14967 21131
rect 16221 21097 16255 21131
rect 16405 21097 16439 21131
rect 23305 21097 23339 21131
rect 24685 21097 24719 21131
rect 28273 21097 28307 21131
rect 30113 21097 30147 21131
rect 32689 21097 32723 21131
rect 33425 21097 33459 21131
rect 20545 20961 20579 20995
rect 21557 20961 21591 20995
rect 25513 20961 25547 20995
rect 26709 20961 26743 20995
rect 29653 20961 29687 20995
rect 31401 20961 31435 20995
rect 32965 20961 32999 20995
rect 35265 20961 35299 20995
rect 45201 20961 45235 20995
rect 46305 20961 46339 20995
rect 48145 20961 48179 20995
rect 10425 20893 10459 20927
rect 12633 20893 12667 20927
rect 12909 20893 12943 20927
rect 14105 20893 14139 20927
rect 14841 20893 14875 20927
rect 17417 20893 17451 20927
rect 18153 20893 18187 20927
rect 20269 20893 20303 20927
rect 24501 20893 24535 20927
rect 25329 20893 25363 20927
rect 29745 20893 29779 20927
rect 32045 20893 32079 20927
rect 32505 20893 32539 20927
rect 33609 20893 33643 20927
rect 36737 20893 36771 20927
rect 42901 20893 42935 20927
rect 43269 20893 43303 20927
rect 45661 20893 45695 20927
rect 10701 20825 10735 20859
rect 16037 20825 16071 20859
rect 21833 20825 21867 20859
rect 28089 20825 28123 20859
rect 28289 20825 28323 20859
rect 31493 20825 31527 20859
rect 35357 20825 35391 20859
rect 36277 20825 36311 20859
rect 45753 20825 45787 20859
rect 46489 20825 46523 20859
rect 12817 20757 12851 20791
rect 14289 20757 14323 20791
rect 16247 20757 16281 20791
rect 17601 20757 17635 20791
rect 18245 20757 18279 20791
rect 28457 20757 28491 20791
rect 36829 20757 36863 20791
rect 43913 20757 43947 20791
rect 10517 20553 10551 20587
rect 12817 20553 12851 20587
rect 32413 20553 32447 20587
rect 43269 20553 43303 20587
rect 44097 20553 44131 20587
rect 14105 20485 14139 20519
rect 14321 20485 14355 20519
rect 16865 20485 16899 20519
rect 17081 20485 17115 20519
rect 18337 20485 18371 20519
rect 19993 20485 20027 20519
rect 27997 20485 28031 20519
rect 30021 20485 30055 20519
rect 35081 20485 35115 20519
rect 43729 20485 43763 20519
rect 45385 20485 45419 20519
rect 47961 20485 47995 20519
rect 10517 20417 10551 20451
rect 11713 20417 11747 20451
rect 12814 20417 12848 20451
rect 13185 20417 13219 20451
rect 15025 20417 15059 20451
rect 15669 20417 15703 20451
rect 22017 20417 22051 20451
rect 25145 20417 25179 20451
rect 25881 20417 25915 20451
rect 26985 20417 27019 20451
rect 29929 20417 29963 20451
rect 32321 20417 32355 20451
rect 33517 20417 33551 20451
rect 43085 20417 43119 20451
rect 43269 20417 43303 20451
rect 43913 20417 43947 20451
rect 44189 20417 44223 20451
rect 13277 20349 13311 20383
rect 18153 20349 18187 20383
rect 22109 20349 22143 20383
rect 25973 20349 26007 20383
rect 27261 20349 27295 20383
rect 27721 20349 27755 20383
rect 34897 20349 34931 20383
rect 35357 20349 35391 20383
rect 45201 20349 45235 20383
rect 45661 20349 45695 20383
rect 14473 20281 14507 20315
rect 17233 20281 17267 20315
rect 48145 20281 48179 20315
rect 11529 20213 11563 20247
rect 12633 20213 12667 20247
rect 14289 20213 14323 20247
rect 15117 20213 15151 20247
rect 15761 20213 15795 20247
rect 17049 20213 17083 20247
rect 22385 20213 22419 20247
rect 25145 20213 25179 20247
rect 26249 20213 26283 20247
rect 29469 20213 29503 20247
rect 33609 20213 33643 20247
rect 12817 20009 12851 20043
rect 14289 20009 14323 20043
rect 14473 20009 14507 20043
rect 27353 20009 27387 20043
rect 28181 20009 28215 20043
rect 45017 20009 45051 20043
rect 46857 20009 46891 20043
rect 34713 19941 34747 19975
rect 45661 19941 45695 19975
rect 15761 19873 15795 19907
rect 16957 19873 16991 19907
rect 20085 19873 20119 19907
rect 25605 19873 25639 19907
rect 29561 19873 29595 19907
rect 32965 19873 32999 19907
rect 35909 19873 35943 19907
rect 2053 19805 2087 19839
rect 11069 19805 11103 19839
rect 13277 19805 13311 19839
rect 15577 19805 15611 19839
rect 17877 19805 17911 19839
rect 19625 19805 19659 19839
rect 24409 19805 24443 19839
rect 28181 19805 28215 19839
rect 28457 19805 28491 19839
rect 32597 19805 32631 19839
rect 33425 19805 33459 19839
rect 33609 19805 33643 19839
rect 33793 19805 33827 19839
rect 34897 19805 34931 19839
rect 35449 19805 35483 19839
rect 44005 19805 44039 19839
rect 44097 19805 44131 19839
rect 45017 19805 45051 19839
rect 45201 19805 45235 19839
rect 45845 19805 45879 19839
rect 46581 19805 46615 19839
rect 47409 19805 47443 19839
rect 11345 19737 11379 19771
rect 13369 19737 13403 19771
rect 14105 19737 14139 19771
rect 19809 19737 19843 19771
rect 25881 19737 25915 19771
rect 29745 19737 29779 19771
rect 31401 19737 31435 19771
rect 32229 19737 32263 19771
rect 32781 19737 32815 19771
rect 35633 19737 35667 19771
rect 44281 19737 44315 19771
rect 46305 19737 46339 19771
rect 46673 19737 46707 19771
rect 14305 19669 14339 19703
rect 18061 19669 18095 19703
rect 24593 19669 24627 19703
rect 28365 19669 28399 19703
rect 46489 19669 46523 19703
rect 47501 19669 47535 19703
rect 13369 19465 13403 19499
rect 20453 19465 20487 19499
rect 24501 19465 24535 19499
rect 28273 19465 28307 19499
rect 28917 19465 28951 19499
rect 44005 19465 44039 19499
rect 47685 19465 47719 19499
rect 12909 19397 12943 19431
rect 19809 19397 19843 19431
rect 33517 19397 33551 19431
rect 1777 19329 1811 19363
rect 12173 19329 12207 19363
rect 14013 19329 14047 19363
rect 14197 19329 14231 19363
rect 14289 19329 14323 19363
rect 14933 19329 14967 19363
rect 19717 19329 19751 19363
rect 20361 19329 20395 19363
rect 21005 19329 21039 19363
rect 28089 19329 28123 19363
rect 28825 19329 28859 19363
rect 32505 19329 32539 19363
rect 33333 19329 33367 19363
rect 35817 19329 35851 19363
rect 43913 19329 43947 19363
rect 44097 19329 44131 19363
rect 45937 19329 45971 19363
rect 46305 19329 46339 19363
rect 46581 19329 46615 19363
rect 46857 19329 46891 19363
rect 47593 19329 47627 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 17509 19261 17543 19295
rect 17785 19261 17819 19295
rect 19257 19261 19291 19295
rect 22753 19261 22787 19295
rect 23029 19261 23063 19295
rect 32597 19261 32631 19295
rect 32873 19261 32907 19295
rect 33793 19261 33827 19295
rect 13277 19193 13311 19227
rect 13829 19193 13863 19227
rect 12357 19125 12391 19159
rect 15025 19125 15059 19159
rect 21097 19125 21131 19159
rect 35633 19125 35667 19159
rect 45477 19125 45511 19159
rect 46213 19125 46247 19159
rect 2237 18921 2271 18955
rect 18613 18921 18647 18955
rect 23673 18921 23707 18955
rect 33517 18921 33551 18955
rect 32873 18853 32907 18887
rect 15945 18785 15979 18819
rect 18153 18785 18187 18819
rect 20729 18785 20763 18819
rect 32321 18785 32355 18819
rect 42625 18785 42659 18819
rect 46305 18785 46339 18819
rect 46489 18785 46523 18819
rect 48145 18785 48179 18819
rect 2145 18717 2179 18751
rect 13001 18717 13035 18751
rect 14105 18717 14139 18751
rect 14933 18717 14967 18751
rect 15761 18717 15795 18751
rect 18245 18717 18279 18751
rect 20545 18717 20579 18751
rect 22845 18717 22879 18751
rect 23581 18717 23615 18751
rect 27261 18717 27295 18751
rect 31033 18717 31067 18751
rect 31125 18717 31159 18751
rect 31309 18717 31343 18751
rect 31401 18717 31435 18751
rect 32137 18717 32171 18751
rect 32781 18717 32815 18751
rect 32965 18717 32999 18751
rect 33425 18717 33459 18751
rect 33609 18717 33643 18751
rect 37105 18717 37139 18751
rect 37197 18717 37231 18751
rect 37289 18717 37323 18751
rect 45109 18717 45143 18751
rect 45293 18717 45327 18751
rect 17601 18649 17635 18683
rect 22385 18649 22419 18683
rect 27537 18649 27571 18683
rect 31953 18649 31987 18683
rect 36645 18649 36679 18683
rect 42809 18649 42843 18683
rect 44465 18649 44499 18683
rect 13185 18581 13219 18615
rect 14197 18581 14231 18615
rect 14749 18581 14783 18615
rect 23029 18581 23063 18615
rect 31401 18581 31435 18615
rect 37473 18581 37507 18615
rect 45201 18581 45235 18615
rect 1593 18377 1627 18411
rect 31309 18377 31343 18411
rect 31401 18377 31435 18411
rect 37105 18377 37139 18411
rect 42809 18377 42843 18411
rect 47961 18377 47995 18411
rect 17233 18309 17267 18343
rect 31217 18309 31251 18343
rect 34897 18309 34931 18343
rect 37473 18309 37507 18343
rect 45385 18309 45419 18343
rect 47777 18309 47811 18343
rect 1409 18241 1443 18275
rect 13093 18241 13127 18275
rect 17141 18241 17175 18275
rect 17877 18241 17911 18275
rect 18061 18241 18095 18275
rect 21097 18241 21131 18275
rect 24961 18241 24995 18275
rect 26157 18241 26191 18275
rect 27169 18241 27203 18275
rect 27813 18241 27847 18275
rect 28733 18241 28767 18275
rect 30297 18241 30331 18275
rect 30481 18241 30515 18275
rect 31585 18241 31619 18275
rect 32321 18241 32355 18275
rect 32965 18241 32999 18275
rect 34713 18241 34747 18275
rect 36645 18241 36679 18275
rect 42717 18241 42751 18275
rect 47593 18241 47627 18275
rect 13369 18173 13403 18207
rect 14841 18173 14875 18207
rect 21189 18173 21223 18207
rect 21833 18173 21867 18207
rect 22109 18173 22143 18207
rect 26985 18173 27019 18207
rect 32137 18173 32171 18207
rect 35909 18173 35943 18207
rect 37289 18173 37323 18207
rect 37749 18173 37783 18207
rect 43913 18173 43947 18207
rect 44741 18173 44775 18207
rect 45201 18173 45235 18207
rect 45661 18173 45695 18207
rect 26341 18105 26375 18139
rect 27353 18105 27387 18139
rect 31033 18105 31067 18139
rect 17877 18037 17911 18071
rect 23581 18037 23615 18071
rect 24777 18037 24811 18071
rect 27813 18037 27847 18071
rect 28825 18037 28859 18071
rect 30389 18037 30423 18071
rect 32505 18037 32539 18071
rect 33057 18037 33091 18071
rect 36921 18037 36955 18071
rect 17417 17833 17451 17867
rect 21189 17833 21223 17867
rect 22569 17833 22603 17867
rect 26617 17833 26651 17867
rect 28917 17833 28951 17867
rect 31217 17833 31251 17867
rect 45661 17833 45695 17867
rect 18429 17697 18463 17731
rect 20913 17697 20947 17731
rect 25237 17697 25271 17731
rect 25421 17697 25455 17731
rect 27169 17697 27203 17731
rect 30481 17697 30515 17731
rect 32965 17697 32999 17731
rect 45477 17697 45511 17731
rect 46305 17697 46339 17731
rect 12817 17629 12851 17663
rect 13369 17629 13403 17663
rect 15485 17629 15519 17663
rect 15761 17629 15795 17663
rect 15945 17629 15979 17663
rect 16865 17629 16899 17663
rect 17141 17629 17175 17663
rect 18153 17629 18187 17663
rect 20821 17629 20855 17663
rect 22477 17629 22511 17663
rect 23581 17629 23615 17663
rect 25145 17629 25179 17663
rect 25329 17629 25363 17663
rect 26433 17629 26467 17663
rect 29561 17629 29595 17663
rect 30389 17629 30423 17663
rect 30573 17629 30607 17663
rect 31125 17629 31159 17663
rect 31309 17629 31343 17663
rect 31953 17629 31987 17663
rect 32321 17629 32355 17663
rect 35449 17629 35483 17663
rect 36185 17629 36219 17663
rect 45017 17629 45051 17663
rect 45385 17629 45419 17663
rect 17233 17561 17267 17595
rect 17877 17561 17911 17595
rect 18061 17561 18095 17595
rect 26249 17561 26283 17595
rect 27445 17561 27479 17595
rect 35541 17561 35575 17595
rect 36369 17561 36403 17595
rect 38025 17561 38059 17595
rect 46489 17561 46523 17595
rect 48145 17561 48179 17595
rect 12817 17493 12851 17527
rect 13461 17493 13495 17527
rect 15301 17493 15335 17527
rect 17049 17493 17083 17527
rect 18245 17493 18279 17527
rect 23765 17493 23799 17527
rect 24961 17493 24995 17527
rect 29653 17493 29687 17527
rect 17141 17289 17175 17323
rect 22937 17289 22971 17323
rect 27077 17289 27111 17323
rect 31493 17289 31527 17323
rect 46305 17289 46339 17323
rect 46949 17289 46983 17323
rect 16773 17221 16807 17255
rect 16989 17221 17023 17255
rect 17877 17221 17911 17255
rect 21833 17221 21867 17255
rect 23121 17221 23155 17255
rect 12449 17153 12483 17187
rect 15117 17153 15151 17187
rect 15945 17153 15979 17187
rect 22017 17153 22051 17187
rect 22109 17153 22143 17187
rect 23029 17153 23063 17187
rect 24133 17153 24167 17187
rect 26985 17153 27019 17187
rect 27169 17153 27203 17187
rect 27629 17153 27663 17187
rect 31401 17153 31435 17187
rect 31585 17153 31619 17187
rect 43729 17153 43763 17187
rect 46213 17153 46247 17187
rect 46397 17153 46431 17187
rect 46857 17153 46891 17187
rect 47593 17153 47627 17187
rect 12725 17085 12759 17119
rect 17601 17085 17635 17119
rect 24409 17085 24443 17119
rect 27905 17085 27939 17119
rect 29653 17085 29687 17119
rect 43913 17085 43947 17119
rect 45385 17085 45419 17119
rect 22753 17017 22787 17051
rect 2053 16949 2087 16983
rect 14197 16949 14231 16983
rect 15117 16949 15151 16983
rect 16037 16949 16071 16983
rect 16957 16949 16991 16983
rect 19349 16949 19383 16983
rect 21833 16949 21867 16983
rect 23305 16949 23339 16983
rect 25881 16949 25915 16983
rect 47685 16949 47719 16983
rect 13001 16745 13035 16779
rect 16773 16745 16807 16779
rect 17417 16745 17451 16779
rect 18337 16745 18371 16779
rect 22661 16745 22695 16779
rect 22845 16745 22879 16779
rect 25053 16745 25087 16779
rect 25605 16745 25639 16779
rect 27077 16745 27111 16779
rect 27629 16745 27663 16779
rect 43913 16745 43947 16779
rect 23305 16677 23339 16711
rect 1409 16609 1443 16643
rect 1869 16609 1903 16643
rect 12725 16609 12759 16643
rect 15025 16609 15059 16643
rect 15301 16609 15335 16643
rect 19717 16609 19751 16643
rect 23857 16609 23891 16643
rect 24501 16609 24535 16643
rect 26893 16609 26927 16643
rect 46305 16609 46339 16643
rect 12633 16541 12667 16575
rect 17233 16541 17267 16575
rect 18061 16541 18095 16575
rect 18153 16541 18187 16575
rect 23581 16541 23615 16575
rect 23673 16541 23707 16575
rect 24685 16541 24719 16575
rect 25513 16541 25547 16575
rect 26801 16541 26835 16575
rect 27813 16541 27847 16575
rect 43821 16541 43855 16575
rect 1593 16473 1627 16507
rect 19901 16473 19935 16507
rect 21557 16473 21591 16507
rect 22477 16473 22511 16507
rect 24777 16473 24811 16507
rect 46489 16473 46523 16507
rect 48145 16473 48179 16507
rect 22687 16405 22721 16439
rect 23489 16405 23523 16439
rect 24869 16405 24903 16439
rect 2145 16201 2179 16235
rect 18153 16201 18187 16235
rect 18797 16201 18831 16235
rect 19901 16201 19935 16235
rect 17969 16133 18003 16167
rect 24409 16133 24443 16167
rect 2053 16065 2087 16099
rect 15301 16065 15335 16099
rect 18245 16065 18279 16099
rect 18705 16065 18739 16099
rect 19809 16065 19843 16099
rect 21005 16065 21039 16099
rect 25513 16065 25547 16099
rect 44741 16065 44775 16099
rect 47777 16065 47811 16099
rect 21097 15997 21131 16031
rect 21833 15997 21867 16031
rect 22109 15997 22143 16031
rect 24869 15997 24903 16031
rect 44925 15997 44959 16031
rect 46121 15997 46155 16031
rect 17969 15929 18003 15963
rect 24777 15929 24811 15963
rect 25329 15929 25363 15963
rect 15393 15861 15427 15895
rect 23581 15861 23615 15895
rect 21005 15657 21039 15691
rect 22477 15657 22511 15691
rect 45109 15657 45143 15691
rect 47685 15657 47719 15691
rect 15209 15521 15243 15555
rect 15393 15521 15427 15555
rect 2053 15453 2087 15487
rect 14289 15453 14323 15487
rect 18429 15453 18463 15487
rect 19257 15453 19291 15487
rect 21005 15453 21039 15487
rect 21189 15453 21223 15487
rect 21649 15453 21683 15487
rect 22385 15453 22419 15487
rect 24869 15453 24903 15487
rect 45017 15453 45051 15487
rect 17049 15385 17083 15419
rect 14381 15317 14415 15351
rect 18521 15317 18555 15351
rect 19349 15317 19383 15351
rect 21833 15317 21867 15351
rect 24961 15317 24995 15351
rect 22201 15113 22235 15147
rect 13553 15045 13587 15079
rect 21833 15045 21867 15079
rect 22033 15045 22067 15079
rect 1777 14977 1811 15011
rect 13369 14977 13403 15011
rect 15669 14977 15703 15011
rect 19165 14977 19199 15011
rect 19441 14977 19475 15011
rect 19625 14977 19659 15011
rect 22845 14977 22879 15011
rect 46581 14977 46615 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 13829 14909 13863 14943
rect 16681 14909 16715 14943
rect 16865 14909 16899 14943
rect 18061 14909 18095 14943
rect 15761 14773 15795 14807
rect 18981 14773 19015 14807
rect 22017 14773 22051 14807
rect 22937 14773 22971 14807
rect 46673 14773 46707 14807
rect 2237 14569 2271 14603
rect 21005 14569 21039 14603
rect 22293 14569 22327 14603
rect 22477 14569 22511 14603
rect 15301 14433 15335 14467
rect 15485 14433 15519 14467
rect 17877 14433 17911 14467
rect 18153 14433 18187 14467
rect 19533 14433 19567 14467
rect 23581 14433 23615 14467
rect 23857 14433 23891 14467
rect 24685 14433 24719 14467
rect 2145 14365 2179 14399
rect 14657 14365 14691 14399
rect 17785 14365 17819 14399
rect 19257 14365 19291 14399
rect 21465 14365 21499 14399
rect 21649 14365 21683 14399
rect 23489 14365 23523 14399
rect 24409 14365 24443 14399
rect 31217 14365 31251 14399
rect 45017 14365 45051 14399
rect 17141 14297 17175 14331
rect 22109 14297 22143 14331
rect 22309 14297 22343 14331
rect 45201 14297 45235 14331
rect 46857 14297 46891 14331
rect 14749 14229 14783 14263
rect 21649 14229 21683 14263
rect 26157 14229 26191 14263
rect 31309 14229 31343 14263
rect 15577 14025 15611 14059
rect 23581 14025 23615 14059
rect 24317 14025 24351 14059
rect 25053 14025 25087 14059
rect 45201 14025 45235 14059
rect 17877 13957 17911 13991
rect 15485 13889 15519 13923
rect 21833 13889 21867 13923
rect 24317 13889 24351 13923
rect 24961 13889 24995 13923
rect 45109 13889 45143 13923
rect 17601 13821 17635 13855
rect 19625 13821 19659 13855
rect 22090 13685 22124 13719
rect 47777 13685 47811 13719
rect 17969 13481 18003 13515
rect 19441 13481 19475 13515
rect 21833 13481 21867 13515
rect 15209 13345 15243 13379
rect 15485 13345 15519 13379
rect 21649 13345 21683 13379
rect 30389 13345 30423 13379
rect 30573 13345 30607 13379
rect 46305 13345 46339 13379
rect 46489 13345 46523 13379
rect 15025 13277 15059 13311
rect 18153 13277 18187 13311
rect 19441 13277 19475 13311
rect 21557 13277 21591 13311
rect 32229 13209 32263 13243
rect 48145 13209 48179 13243
rect 1409 12801 1443 12835
rect 1593 12597 1627 12631
rect 47685 12189 47719 12223
rect 22109 11713 22143 11747
rect 22293 11645 22327 11679
rect 23949 11645 23983 11679
rect 22293 11305 22327 11339
rect 46305 11169 46339 11203
rect 22201 11101 22235 11135
rect 46489 11033 46523 11067
rect 48145 11033 48179 11067
rect 47593 10625 47627 10659
rect 47041 10421 47075 10455
rect 47685 10421 47719 10455
rect 46305 10081 46339 10115
rect 46489 10081 46523 10115
rect 48145 10081 48179 10115
rect 47869 9537 47903 9571
rect 48053 9401 48087 9435
rect 47777 8857 47811 8891
rect 47869 8789 47903 8823
rect 46949 8449 46983 8483
rect 46765 8313 46799 8347
rect 46489 7905 46523 7939
rect 47317 7905 47351 7939
rect 45477 7769 45511 7803
rect 45569 7769 45603 7803
rect 47041 7769 47075 7803
rect 47133 7769 47167 7803
rect 46673 7497 46707 7531
rect 47961 7497 47995 7531
rect 46213 7361 46247 7395
rect 48145 7361 48179 7395
rect 45937 7157 45971 7191
rect 46305 7157 46339 7191
rect 47317 6817 47351 6851
rect 47593 6749 47627 6783
rect 48053 6409 48087 6443
rect 47961 6273 47995 6307
rect 41705 5729 41739 5763
rect 42165 5729 42199 5763
rect 43177 5729 43211 5763
rect 36737 5661 36771 5695
rect 37197 5593 37231 5627
rect 37289 5593 37323 5627
rect 38209 5593 38243 5627
rect 42257 5593 42291 5627
rect 42441 5321 42475 5355
rect 48053 5321 48087 5355
rect 37749 5253 37783 5287
rect 39773 5185 39807 5219
rect 40417 5185 40451 5219
rect 42625 5185 42659 5219
rect 47869 5185 47903 5219
rect 37657 5117 37691 5151
rect 38485 5117 38519 5151
rect 39865 4981 39899 5015
rect 40509 4981 40543 5015
rect 37105 4777 37139 4811
rect 39221 4777 39255 4811
rect 39957 4641 39991 4675
rect 41797 4641 41831 4675
rect 42625 4641 42659 4675
rect 43177 4641 43211 4675
rect 47593 4641 47627 4675
rect 14289 4573 14323 4607
rect 18337 4573 18371 4607
rect 20637 4573 20671 4607
rect 37289 4573 37323 4607
rect 39129 4573 39163 4607
rect 46673 4573 46707 4607
rect 47317 4573 47351 4607
rect 40141 4505 40175 4539
rect 42717 4505 42751 4539
rect 14381 4437 14415 4471
rect 18429 4437 18463 4471
rect 20729 4437 20763 4471
rect 46765 4437 46799 4471
rect 37749 4233 37783 4267
rect 27169 4165 27203 4199
rect 40325 4165 40359 4199
rect 46673 4165 46707 4199
rect 47777 4165 47811 4199
rect 2053 4097 2087 4131
rect 7205 4097 7239 4131
rect 11897 4097 11931 4131
rect 13277 4097 13311 4131
rect 13369 4097 13403 4131
rect 13921 4097 13955 4131
rect 14013 4097 14047 4131
rect 14565 4097 14599 4131
rect 15209 4097 15243 4131
rect 15853 4097 15887 4131
rect 16681 4097 16715 4131
rect 17325 4097 17359 4131
rect 17969 4097 18003 4131
rect 18613 4097 18647 4131
rect 19257 4097 19291 4131
rect 19901 4097 19935 4131
rect 20545 4097 20579 4131
rect 21833 4097 21867 4131
rect 21925 4097 21959 4131
rect 22753 4097 22787 4131
rect 24133 4097 24167 4131
rect 24777 4097 24811 4131
rect 37289 4097 37323 4131
rect 39221 4097 39255 4131
rect 39405 4097 39439 4131
rect 40509 4097 40543 4131
rect 41153 4097 41187 4131
rect 41245 4097 41279 4131
rect 42441 4097 42475 4131
rect 27077 4029 27111 4063
rect 28089 4029 28123 4063
rect 39865 4029 39899 4063
rect 42901 4029 42935 4063
rect 46857 3961 46891 3995
rect 2145 3893 2179 3927
rect 2881 3893 2915 3927
rect 7297 3893 7331 3927
rect 11989 3893 12023 3927
rect 14657 3893 14691 3927
rect 15301 3893 15335 3927
rect 15945 3893 15979 3927
rect 16773 3893 16807 3927
rect 17417 3893 17451 3927
rect 18061 3893 18095 3927
rect 18705 3893 18739 3927
rect 19349 3893 19383 3927
rect 19993 3893 20027 3927
rect 20637 3893 20671 3927
rect 22845 3893 22879 3927
rect 24225 3893 24259 3927
rect 24869 3893 24903 3927
rect 25605 3893 25639 3927
rect 37381 3893 37415 3927
rect 40693 3893 40727 3927
rect 42533 3893 42567 3927
rect 46121 3893 46155 3927
rect 47869 3893 47903 3927
rect 14841 3621 14875 3655
rect 15485 3621 15519 3655
rect 17417 3621 17451 3655
rect 18061 3621 18095 3655
rect 22753 3621 22787 3655
rect 40049 3621 40083 3655
rect 3985 3553 4019 3587
rect 11253 3553 11287 3587
rect 11529 3553 11563 3587
rect 16129 3553 16163 3587
rect 24685 3553 24719 3587
rect 24869 3553 24903 3587
rect 25145 3553 25179 3587
rect 33885 3553 33919 3587
rect 41797 3553 41831 3587
rect 44189 3553 44223 3587
rect 46305 3553 46339 3587
rect 46489 3553 46523 3587
rect 2697 3485 2731 3519
rect 6193 3485 6227 3519
rect 6653 3485 6687 3519
rect 7481 3485 7515 3519
rect 10425 3485 10459 3519
rect 11069 3485 11103 3519
rect 13553 3485 13587 3519
rect 14105 3485 14139 3519
rect 14749 3485 14783 3519
rect 15393 3485 15427 3519
rect 16037 3485 16071 3519
rect 16681 3485 16715 3519
rect 17325 3485 17359 3519
rect 17969 3485 18003 3519
rect 19441 3485 19475 3519
rect 19533 3485 19567 3519
rect 20269 3485 20303 3519
rect 20729 3485 20763 3519
rect 20821 3485 20855 3519
rect 22017 3485 22051 3519
rect 22845 3485 22879 3519
rect 23673 3485 23707 3519
rect 27169 3485 27203 3519
rect 33057 3485 33091 3519
rect 40233 3485 40267 3519
rect 41061 3485 41095 3519
rect 43361 3485 43395 3519
rect 45201 3485 45235 3519
rect 45661 3485 45695 3519
rect 1869 3417 1903 3451
rect 2237 3417 2271 3451
rect 9413 3417 9447 3451
rect 16773 3417 16807 3451
rect 41245 3417 41279 3451
rect 48145 3417 48179 3451
rect 2789 3349 2823 3383
rect 6745 3349 6779 3383
rect 9689 3349 9723 3383
rect 10517 3349 10551 3383
rect 14197 3349 14231 3383
rect 26985 3349 27019 3383
rect 33149 3349 33183 3383
rect 43453 3349 43487 3383
rect 45753 3349 45787 3383
rect 13001 3145 13035 3179
rect 18337 3145 18371 3179
rect 21925 3145 21959 3179
rect 22569 3145 22603 3179
rect 39865 3145 39899 3179
rect 41153 3145 41187 3179
rect 1961 3077 1995 3111
rect 7389 3077 7423 3111
rect 13829 3077 13863 3111
rect 19533 3077 19567 3111
rect 23397 3077 23431 3111
rect 27169 3077 27203 3111
rect 28089 3077 28123 3111
rect 33149 3077 33183 3111
rect 42625 3077 42659 3111
rect 45385 3077 45419 3111
rect 1777 3009 1811 3043
rect 7205 3009 7239 3043
rect 10977 3009 11011 3043
rect 12081 3009 12115 3043
rect 12909 3009 12943 3043
rect 13645 3009 13679 3043
rect 18253 3015 18287 3049
rect 21189 3009 21223 3043
rect 21833 3009 21867 3043
rect 22485 3009 22519 3043
rect 23213 3009 23247 3043
rect 26249 3009 26283 3043
rect 32965 3009 32999 3043
rect 39405 3009 39439 3043
rect 40049 3009 40083 3043
rect 41797 3009 41831 3043
rect 42441 3009 42475 3043
rect 45201 3009 45235 3043
rect 47777 3009 47811 3043
rect 2237 2941 2271 2975
rect 7757 2941 7791 2975
rect 11989 2941 12023 2975
rect 12449 2941 12483 2975
rect 15117 2941 15151 2975
rect 19349 2941 19383 2975
rect 23673 2941 23707 2975
rect 27077 2941 27111 2975
rect 33517 2941 33551 2975
rect 40509 2941 40543 2975
rect 40693 2941 40727 2975
rect 43177 2941 43211 2975
rect 47041 2941 47075 2975
rect 39221 2873 39255 2907
rect 41613 2873 41647 2907
rect 47961 2873 47995 2907
rect 9781 2805 9815 2839
rect 26341 2805 26375 2839
rect 3985 2601 4019 2635
rect 14289 2601 14323 2635
rect 19349 2601 19383 2635
rect 20913 2601 20947 2635
rect 22385 2601 22419 2635
rect 23397 2601 23431 2635
rect 27261 2601 27295 2635
rect 27445 2601 27479 2635
rect 39221 2601 39255 2635
rect 40325 2601 40359 2635
rect 40601 2601 40635 2635
rect 48053 2601 48087 2635
rect 25053 2533 25087 2567
rect 35541 2533 35575 2567
rect 36461 2533 36495 2567
rect 38301 2533 38335 2567
rect 41337 2533 41371 2567
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2789 2465 2823 2499
rect 6561 2465 6595 2499
rect 6745 2465 6779 2499
rect 7113 2465 7147 2499
rect 9137 2465 9171 2499
rect 9873 2465 9907 2499
rect 26433 2465 26467 2499
rect 40325 2465 40359 2499
rect 46489 2465 46523 2499
rect 3801 2397 3835 2431
rect 5457 2397 5491 2431
rect 14197 2397 14231 2431
rect 14841 2397 14875 2431
rect 16681 2397 16715 2431
rect 19257 2397 19291 2431
rect 23581 2397 23615 2431
rect 26985 2397 27019 2431
rect 28457 2397 28491 2431
rect 29929 2397 29963 2431
rect 35725 2397 35759 2431
rect 38117 2397 38151 2431
rect 40049 2397 40083 2431
rect 41153 2397 41187 2431
rect 43637 2397 43671 2431
rect 43913 2397 43947 2431
rect 46213 2397 46247 2431
rect 9321 2329 9355 2363
rect 15669 2329 15703 2363
rect 20821 2329 20855 2363
rect 22293 2329 22327 2363
rect 24869 2329 24903 2363
rect 26249 2329 26283 2363
rect 36277 2329 36311 2363
rect 39129 2329 39163 2363
rect 45385 2329 45419 2363
rect 47777 2329 47811 2363
rect 5273 2261 5307 2295
rect 14933 2261 14967 2295
rect 15761 2261 15795 2295
rect 16865 2261 16899 2295
rect 28641 2261 28675 2295
rect 29745 2261 29779 2295
rect 45477 2261 45511 2295
<< metal1 >>
rect 18598 47404 18604 47456
rect 18656 47444 18662 47456
rect 22554 47444 22560 47456
rect 18656 47416 22560 47444
rect 18656 47404 18662 47416
rect 22554 47404 22560 47416
rect 22612 47404 22618 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 14277 47243 14335 47249
rect 14277 47209 14289 47243
rect 14323 47240 14335 47243
rect 17218 47240 17224 47252
rect 14323 47212 17224 47240
rect 14323 47209 14335 47212
rect 14277 47203 14335 47209
rect 17218 47200 17224 47212
rect 17276 47200 17282 47252
rect 20806 47200 20812 47252
rect 20864 47240 20870 47252
rect 22465 47243 22523 47249
rect 22465 47240 22477 47243
rect 20864 47212 22477 47240
rect 20864 47200 20870 47212
rect 22465 47209 22477 47212
rect 22511 47209 22523 47243
rect 22465 47203 22523 47209
rect 22554 47200 22560 47252
rect 22612 47240 22618 47252
rect 44085 47243 44143 47249
rect 44085 47240 44097 47243
rect 22612 47212 44097 47240
rect 22612 47200 22618 47212
rect 44085 47209 44097 47212
rect 44131 47209 44143 47243
rect 44085 47203 44143 47209
rect 3053 47175 3111 47181
rect 3053 47141 3065 47175
rect 3099 47172 3111 47175
rect 29917 47175 29975 47181
rect 3099 47144 26234 47172
rect 3099 47141 3111 47144
rect 3053 47135 3111 47141
rect 12250 47064 12256 47116
rect 12308 47104 12314 47116
rect 12345 47107 12403 47113
rect 12345 47104 12357 47107
rect 12308 47076 12357 47104
rect 12308 47064 12314 47076
rect 12345 47073 12357 47076
rect 12391 47073 12403 47107
rect 12345 47067 12403 47073
rect 12621 47107 12679 47113
rect 12621 47073 12633 47107
rect 12667 47104 12679 47107
rect 19242 47104 19248 47116
rect 12667 47076 19248 47104
rect 12667 47073 12679 47076
rect 12621 47067 12679 47073
rect 19242 47064 19248 47076
rect 19300 47064 19306 47116
rect 26206 47104 26234 47144
rect 29917 47141 29929 47175
rect 29963 47172 29975 47175
rect 30098 47172 30104 47184
rect 29963 47144 30104 47172
rect 29963 47141 29975 47144
rect 29917 47135 29975 47141
rect 30098 47132 30104 47144
rect 30156 47132 30162 47184
rect 34790 47172 34796 47184
rect 30208 47144 34796 47172
rect 30208 47104 30236 47144
rect 34790 47132 34796 47144
rect 34848 47132 34854 47184
rect 47394 47132 47400 47184
rect 47452 47172 47458 47184
rect 47949 47175 48007 47181
rect 47949 47172 47961 47175
rect 47452 47144 47961 47172
rect 47452 47132 47458 47144
rect 47949 47141 47961 47144
rect 47995 47141 48007 47175
rect 47949 47135 48007 47141
rect 30742 47104 30748 47116
rect 26206 47076 30236 47104
rect 30703 47076 30748 47104
rect 30742 47064 30748 47076
rect 30800 47064 30806 47116
rect 44450 47104 44456 47116
rect 43272 47076 44456 47104
rect 1765 47039 1823 47045
rect 1765 47005 1777 47039
rect 1811 47036 1823 47039
rect 1946 47036 1952 47048
rect 1811 47008 1952 47036
rect 1811 47005 1823 47008
rect 1765 46999 1823 47005
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4706 47036 4712 47048
rect 4667 47008 4712 47036
rect 3789 46999 3847 47005
rect 4706 46996 4712 47008
rect 4764 46996 4770 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6365 47039 6423 47045
rect 6365 47036 6377 47039
rect 5868 47008 6377 47036
rect 5868 46996 5874 47008
rect 6365 47005 6377 47008
rect 6411 47005 6423 47039
rect 7282 47036 7288 47048
rect 7243 47008 7288 47036
rect 6365 46999 6423 47005
rect 7282 46996 7288 47008
rect 7340 46996 7346 47048
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 9088 47008 9413 47036
rect 9088 46996 9094 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 9401 46999 9459 47005
rect 14093 47039 14151 47045
rect 14093 47005 14105 47039
rect 14139 47005 14151 47039
rect 14093 46999 14151 47005
rect 2038 46968 2044 46980
rect 1999 46940 2044 46968
rect 2038 46928 2044 46940
rect 2096 46928 2102 46980
rect 2777 46971 2835 46977
rect 2777 46937 2789 46971
rect 2823 46937 2835 46971
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 2777 46931 2835 46937
rect 2590 46860 2596 46912
rect 2648 46900 2654 46912
rect 2792 46900 2820 46931
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 4982 46968 4988 46980
rect 4943 46940 4988 46968
rect 4982 46928 4988 46940
rect 5040 46928 5046 46980
rect 6638 46968 6644 46980
rect 6599 46940 6644 46968
rect 6638 46928 6644 46940
rect 6696 46928 6702 46980
rect 9490 46928 9496 46980
rect 9548 46968 9554 46980
rect 9585 46971 9643 46977
rect 9585 46968 9597 46971
rect 9548 46940 9597 46968
rect 9548 46928 9554 46940
rect 9585 46937 9597 46940
rect 9631 46937 9643 46971
rect 9585 46931 9643 46937
rect 7466 46900 7472 46912
rect 2648 46872 2820 46900
rect 7427 46872 7472 46900
rect 2648 46860 2654 46872
rect 7466 46860 7472 46872
rect 7524 46860 7530 46912
rect 12894 46860 12900 46912
rect 12952 46900 12958 46912
rect 14108 46900 14136 46999
rect 14182 46996 14188 47048
rect 14240 47036 14246 47048
rect 14921 47039 14979 47045
rect 14921 47036 14933 47039
rect 14240 47008 14933 47036
rect 14240 46996 14246 47008
rect 14921 47005 14933 47008
rect 14967 47005 14979 47039
rect 14921 46999 14979 47005
rect 16482 46996 16488 47048
rect 16540 47036 16546 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16540 47008 16681 47036
rect 16540 46996 16546 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16669 46999 16727 47005
rect 16945 47039 17003 47045
rect 16945 47005 16957 47039
rect 16991 47036 17003 47039
rect 20162 47036 20168 47048
rect 16991 47008 20168 47036
rect 16991 47005 17003 47008
rect 16945 46999 17003 47005
rect 20162 46996 20168 47008
rect 20220 46996 20226 47048
rect 20990 47036 20996 47048
rect 20951 47008 20996 47036
rect 20990 46996 20996 47008
rect 21048 46996 21054 47048
rect 22002 47036 22008 47048
rect 21963 47008 22008 47036
rect 22002 46996 22008 47008
rect 22060 46996 22066 47048
rect 22649 47039 22707 47045
rect 22649 47005 22661 47039
rect 22695 47005 22707 47039
rect 24854 47036 24860 47048
rect 24815 47008 24860 47036
rect 22649 46999 22707 47005
rect 15010 46928 15016 46980
rect 15068 46968 15074 46980
rect 15105 46971 15163 46977
rect 15105 46968 15117 46971
rect 15068 46940 15117 46968
rect 15068 46928 15074 46940
rect 15105 46937 15117 46940
rect 15151 46937 15163 46971
rect 15105 46931 15163 46937
rect 19705 46971 19763 46977
rect 19705 46937 19717 46971
rect 19751 46937 19763 46971
rect 19705 46931 19763 46937
rect 20073 46971 20131 46977
rect 20073 46937 20085 46971
rect 20119 46968 20131 46971
rect 20530 46968 20536 46980
rect 20119 46940 20536 46968
rect 20119 46937 20131 46940
rect 20073 46931 20131 46937
rect 12952 46872 14136 46900
rect 12952 46860 12958 46872
rect 18690 46860 18696 46912
rect 18748 46900 18754 46912
rect 19720 46900 19748 46931
rect 20530 46928 20536 46940
rect 20588 46928 20594 46980
rect 22664 46968 22692 46999
rect 24854 46996 24860 47008
rect 24912 46996 24918 47048
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28537 47039 28595 47045
rect 28537 47036 28549 47039
rect 28408 47008 28549 47036
rect 28408 46996 28414 47008
rect 28537 47005 28549 47008
rect 28583 47005 28595 47039
rect 28537 46999 28595 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 30834 46996 30840 47048
rect 30892 47036 30898 47048
rect 31021 47039 31079 47045
rect 31021 47036 31033 47039
rect 30892 47008 31033 47036
rect 30892 46996 30898 47008
rect 31021 47005 31033 47008
rect 31067 47005 31079 47039
rect 31021 46999 31079 47005
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38381 47039 38439 47045
rect 38381 47036 38393 47039
rect 38160 47008 38393 47036
rect 38160 46996 38166 47008
rect 38381 47005 38393 47008
rect 38427 47005 38439 47039
rect 41506 47036 41512 47048
rect 41467 47008 41512 47036
rect 38381 46999 38439 47005
rect 41506 46996 41512 47008
rect 41564 46996 41570 47048
rect 42702 47036 42708 47048
rect 42663 47008 42708 47036
rect 42702 46996 42708 47008
rect 42760 46996 42766 47048
rect 43272 47045 43300 47076
rect 44450 47064 44456 47076
rect 44508 47064 44514 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 43257 47039 43315 47045
rect 43257 47005 43269 47039
rect 43303 47005 43315 47039
rect 43257 46999 43315 47005
rect 43806 46996 43812 47048
rect 43864 47036 43870 47048
rect 43901 47039 43959 47045
rect 43901 47036 43913 47039
rect 43864 47008 43913 47036
rect 43864 46996 43870 47008
rect 43901 47005 43913 47008
rect 43947 47005 43959 47039
rect 43901 46999 43959 47005
rect 45094 46996 45100 47048
rect 45152 47036 45158 47048
rect 45189 47039 45247 47045
rect 45189 47036 45201 47039
rect 45152 47008 45201 47036
rect 45152 46996 45158 47008
rect 45189 47005 45201 47008
rect 45235 47005 45247 47039
rect 45189 46999 45247 47005
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47765 47039 47823 47045
rect 47765 47036 47777 47039
rect 47728 47008 47777 47036
rect 47728 46996 47734 47008
rect 47765 47005 47777 47008
rect 47811 47005 47823 47039
rect 47765 46999 47823 47005
rect 22020 46940 22692 46968
rect 28721 46971 28779 46977
rect 18748 46872 19748 46900
rect 18748 46860 18754 46872
rect 19978 46860 19984 46912
rect 20036 46900 20042 46912
rect 22020 46900 22048 46940
rect 28721 46937 28733 46971
rect 28767 46968 28779 46971
rect 34606 46968 34612 46980
rect 28767 46940 34612 46968
rect 28767 46937 28779 46940
rect 28721 46931 28779 46937
rect 34606 46928 34612 46940
rect 34664 46928 34670 46980
rect 40313 46971 40371 46977
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 40313 46931 40371 46937
rect 20036 46872 22048 46900
rect 20036 46860 20042 46872
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 40402 46928 40408 46980
rect 40460 46968 40466 46980
rect 40497 46971 40555 46977
rect 40497 46968 40509 46971
rect 40460 46940 40509 46968
rect 40460 46928 40466 46940
rect 40497 46937 40509 46940
rect 40543 46937 40555 46971
rect 40497 46931 40555 46937
rect 43346 46928 43352 46980
rect 43404 46968 43410 46980
rect 43441 46971 43499 46977
rect 43441 46968 43453 46971
rect 43404 46940 43453 46968
rect 43404 46928 43410 46940
rect 43441 46937 43453 46940
rect 43487 46937 43499 46971
rect 45370 46968 45376 46980
rect 45331 46940 45376 46968
rect 43441 46931 43499 46937
rect 45370 46928 45376 46940
rect 45428 46928 45434 46980
rect 39356 46872 40356 46900
rect 39356 46860 39362 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 1854 46628 1860 46640
rect 1815 46600 1860 46628
rect 1854 46588 1860 46600
rect 1912 46588 1918 46640
rect 3878 46588 3884 46640
rect 3936 46628 3942 46640
rect 5813 46631 5871 46637
rect 5813 46628 5825 46631
rect 3936 46600 5825 46628
rect 3936 46588 3942 46600
rect 5813 46597 5825 46600
rect 5859 46597 5871 46631
rect 22002 46628 22008 46640
rect 5813 46591 5871 46597
rect 19444 46600 22008 46628
rect 19444 46569 19472 46600
rect 22002 46588 22008 46600
rect 22060 46588 22066 46640
rect 24854 46628 24860 46640
rect 24596 46600 24860 46628
rect 24596 46569 24624 46600
rect 24854 46588 24860 46600
rect 24912 46588 24918 46640
rect 19429 46563 19487 46569
rect 19429 46529 19441 46563
rect 19475 46529 19487 46563
rect 19429 46523 19487 46529
rect 24581 46563 24639 46569
rect 24581 46529 24593 46563
rect 24627 46529 24639 46563
rect 38102 46560 38108 46572
rect 38063 46532 38108 46560
rect 24581 46523 24639 46529
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 41506 46520 41512 46572
rect 41564 46560 41570 46572
rect 42429 46563 42487 46569
rect 42429 46560 42441 46563
rect 41564 46532 42441 46560
rect 41564 46520 41570 46532
rect 42429 46529 42441 46532
rect 42475 46529 42487 46563
rect 47946 46560 47952 46572
rect 47907 46532 47952 46560
rect 42429 46523 42487 46529
rect 47946 46520 47952 46532
rect 48004 46520 48010 46572
rect 3970 46492 3976 46504
rect 3931 46464 3976 46492
rect 3970 46452 3976 46464
rect 4028 46452 4034 46504
rect 4157 46495 4215 46501
rect 4157 46461 4169 46495
rect 4203 46492 4215 46495
rect 5166 46492 5172 46504
rect 4203 46464 5172 46492
rect 4203 46461 4215 46464
rect 4157 46455 4215 46461
rect 5166 46452 5172 46464
rect 5224 46452 5230 46504
rect 10965 46495 11023 46501
rect 10965 46461 10977 46495
rect 11011 46492 11023 46495
rect 11517 46495 11575 46501
rect 11517 46492 11529 46495
rect 11011 46464 11529 46492
rect 11011 46461 11023 46464
rect 10965 46455 11023 46461
rect 11517 46461 11529 46464
rect 11563 46461 11575 46495
rect 11517 46455 11575 46461
rect 11701 46495 11759 46501
rect 11701 46461 11713 46495
rect 11747 46492 11759 46495
rect 11882 46492 11888 46504
rect 11747 46464 11888 46492
rect 11747 46461 11759 46464
rect 11701 46455 11759 46461
rect 11882 46452 11888 46464
rect 11940 46452 11946 46504
rect 11977 46495 12035 46501
rect 11977 46461 11989 46495
rect 12023 46461 12035 46495
rect 11977 46455 12035 46461
rect 11992 46424 12020 46455
rect 13538 46452 13544 46504
rect 13596 46492 13602 46504
rect 13817 46495 13875 46501
rect 13817 46492 13829 46495
rect 13596 46464 13829 46492
rect 13596 46452 13602 46464
rect 13817 46461 13829 46464
rect 13863 46461 13875 46495
rect 13817 46455 13875 46461
rect 14001 46495 14059 46501
rect 14001 46461 14013 46495
rect 14047 46492 14059 46495
rect 14182 46492 14188 46504
rect 14047 46464 14188 46492
rect 14047 46461 14059 46464
rect 14001 46455 14059 46461
rect 14182 46452 14188 46464
rect 14240 46452 14246 46504
rect 14274 46452 14280 46504
rect 14332 46492 14338 46504
rect 19613 46495 19671 46501
rect 14332 46464 14377 46492
rect 14332 46452 14338 46464
rect 19613 46461 19625 46495
rect 19659 46492 19671 46495
rect 19886 46492 19892 46504
rect 19659 46464 19892 46492
rect 19659 46461 19671 46464
rect 19613 46455 19671 46461
rect 19886 46452 19892 46464
rect 19944 46452 19950 46504
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 24762 46492 24768 46504
rect 24723 46464 24768 46492
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 25130 46492 25136 46504
rect 25091 46464 25136 46492
rect 25130 46452 25136 46464
rect 25188 46452 25194 46504
rect 32214 46492 32220 46504
rect 32175 46464 32220 46492
rect 32214 46452 32220 46464
rect 32272 46452 32278 46504
rect 32398 46492 32404 46504
rect 32359 46464 32404 46492
rect 32398 46452 32404 46464
rect 32456 46452 32462 46504
rect 32677 46495 32735 46501
rect 32677 46461 32689 46495
rect 32723 46461 32735 46495
rect 38286 46492 38292 46504
rect 38247 46464 38292 46492
rect 32677 46455 32735 46461
rect 10980 46396 12020 46424
rect 10980 46368 11008 46396
rect 32306 46384 32312 46436
rect 32364 46424 32370 46436
rect 32692 46424 32720 46455
rect 38286 46452 38292 46464
rect 38344 46452 38350 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 42610 46492 42616 46504
rect 42571 46464 42616 46492
rect 42610 46452 42616 46464
rect 42668 46452 42674 46504
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46461 42947 46495
rect 45186 46492 45192 46504
rect 45147 46464 45192 46492
rect 42889 46455 42947 46461
rect 32364 46396 32720 46424
rect 32364 46384 32370 46396
rect 41874 46384 41880 46436
rect 41932 46424 41938 46436
rect 42904 46424 42932 46455
rect 45186 46452 45192 46464
rect 45244 46452 45250 46504
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 45646 46492 45652 46504
rect 45419 46464 45652 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 45646 46452 45652 46464
rect 45704 46452 45710 46504
rect 46842 46492 46848 46504
rect 46803 46464 46848 46492
rect 46842 46452 46848 46464
rect 46900 46452 46906 46504
rect 41932 46396 42932 46424
rect 41932 46384 41938 46396
rect 2130 46356 2136 46368
rect 2091 46328 2136 46356
rect 2130 46316 2136 46328
rect 2188 46316 2194 46368
rect 10962 46316 10968 46368
rect 11020 46316 11026 46368
rect 41046 46316 41052 46368
rect 41104 46356 41110 46368
rect 41325 46359 41383 46365
rect 41325 46356 41337 46359
rect 41104 46328 41337 46356
rect 41104 46316 41110 46328
rect 41325 46325 41337 46328
rect 41371 46325 41383 46359
rect 48038 46356 48044 46368
rect 47999 46328 48044 46356
rect 41325 46319 41383 46325
rect 48038 46316 48044 46328
rect 48096 46316 48102 46368
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 3970 46112 3976 46164
rect 4028 46152 4034 46164
rect 4525 46155 4583 46161
rect 4525 46152 4537 46155
rect 4028 46124 4537 46152
rect 4028 46112 4034 46124
rect 4525 46121 4537 46124
rect 4571 46121 4583 46155
rect 5166 46152 5172 46164
rect 5127 46124 5172 46152
rect 4525 46115 4583 46121
rect 5166 46112 5172 46124
rect 5224 46112 5230 46164
rect 13538 46152 13544 46164
rect 13499 46124 13544 46152
rect 13538 46112 13544 46124
rect 13596 46112 13602 46164
rect 14182 46152 14188 46164
rect 14143 46124 14188 46152
rect 14182 46112 14188 46124
rect 14240 46112 14246 46164
rect 19886 46152 19892 46164
rect 19847 46124 19892 46152
rect 19886 46112 19892 46124
rect 19944 46112 19950 46164
rect 24673 46155 24731 46161
rect 24673 46121 24685 46155
rect 24719 46152 24731 46155
rect 24762 46152 24768 46164
rect 24719 46124 24768 46152
rect 24719 46121 24731 46124
rect 24673 46115 24731 46121
rect 24762 46112 24768 46124
rect 24820 46112 24826 46164
rect 32214 46112 32220 46164
rect 32272 46152 32278 46164
rect 32493 46155 32551 46161
rect 32493 46152 32505 46155
rect 32272 46124 32505 46152
rect 32272 46112 32278 46124
rect 32493 46121 32505 46124
rect 32539 46121 32551 46155
rect 38286 46152 38292 46164
rect 38247 46124 38292 46152
rect 32493 46115 32551 46121
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 46842 46152 46848 46164
rect 43364 46124 46848 46152
rect 11606 45976 11612 46028
rect 11664 46016 11670 46028
rect 11701 46019 11759 46025
rect 11701 46016 11713 46019
rect 11664 45988 11713 46016
rect 11664 45976 11670 45988
rect 11701 45985 11713 45988
rect 11747 45985 11759 46019
rect 11701 45979 11759 45985
rect 20809 46019 20867 46025
rect 20809 45985 20821 46019
rect 20855 46016 20867 46019
rect 20990 46016 20996 46028
rect 20855 45988 20996 46016
rect 20855 45985 20867 45988
rect 20809 45979 20867 45985
rect 20990 45976 20996 45988
rect 21048 45976 21054 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 25774 46016 25780 46028
rect 25735 45988 25780 46016
rect 25774 45976 25780 45988
rect 25832 45976 25838 46028
rect 41046 46016 41052 46028
rect 41007 45988 41052 46016
rect 41046 45976 41052 45988
rect 41104 45976 41110 46028
rect 42518 46016 42524 46028
rect 42479 45988 42524 46016
rect 42518 45976 42524 45988
rect 42576 45976 42582 46028
rect 1762 45908 1768 45960
rect 1820 45948 1826 45960
rect 2041 45951 2099 45957
rect 2041 45948 2053 45951
rect 1820 45920 2053 45948
rect 1820 45908 1826 45920
rect 2041 45917 2053 45920
rect 2087 45917 2099 45951
rect 2041 45911 2099 45917
rect 5077 45951 5135 45957
rect 5077 45917 5089 45951
rect 5123 45948 5135 45951
rect 11974 45948 11980 45960
rect 5123 45920 6914 45948
rect 11935 45920 11980 45948
rect 5123 45917 5135 45920
rect 5077 45911 5135 45917
rect 6886 45812 6914 45920
rect 11974 45908 11980 45920
rect 12032 45908 12038 45960
rect 14090 45948 14096 45960
rect 14003 45920 14096 45948
rect 14090 45908 14096 45920
rect 14148 45948 14154 45960
rect 19797 45951 19855 45957
rect 19797 45948 19809 45951
rect 14148 45920 19809 45948
rect 14148 45908 14154 45920
rect 19797 45917 19809 45920
rect 19843 45948 19855 45951
rect 20254 45948 20260 45960
rect 19843 45920 20260 45948
rect 19843 45917 19855 45920
rect 19797 45911 19855 45917
rect 20254 45908 20260 45920
rect 20312 45908 20318 45960
rect 24581 45951 24639 45957
rect 24581 45917 24593 45951
rect 24627 45917 24639 45951
rect 25222 45948 25228 45960
rect 25183 45920 25228 45948
rect 24581 45911 24639 45917
rect 20990 45880 20996 45892
rect 20951 45852 20996 45880
rect 20990 45840 20996 45852
rect 21048 45840 21054 45892
rect 24486 45812 24492 45824
rect 6886 45784 24492 45812
rect 24486 45772 24492 45784
rect 24544 45812 24550 45824
rect 24596 45812 24624 45911
rect 25222 45908 25228 45920
rect 25280 45908 25286 45960
rect 38194 45948 38200 45960
rect 38155 45920 38200 45948
rect 38194 45908 38200 45920
rect 38252 45908 38258 45960
rect 43364 45957 43392 46124
rect 46842 46112 46848 46124
rect 46900 46112 46906 46164
rect 47578 46084 47584 46096
rect 44284 46056 47584 46084
rect 44284 45957 44312 46056
rect 47578 46044 47584 46056
rect 47636 46044 47642 46096
rect 47026 46016 47032 46028
rect 46987 45988 47032 46016
rect 47026 45976 47032 45988
rect 47084 45976 47090 46028
rect 43349 45951 43407 45957
rect 43349 45917 43361 45951
rect 43395 45917 43407 45951
rect 43349 45911 43407 45917
rect 44269 45951 44327 45957
rect 44269 45917 44281 45951
rect 44315 45917 44327 45951
rect 44269 45911 44327 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45948 45707 45951
rect 45738 45948 45744 45960
rect 45695 45920 45744 45948
rect 45695 45917 45707 45920
rect 45649 45911 45707 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 45830 45908 45836 45960
rect 45888 45948 45894 45960
rect 46293 45951 46351 45957
rect 46293 45948 46305 45951
rect 45888 45920 46305 45948
rect 45888 45908 45894 45920
rect 46293 45917 46305 45920
rect 46339 45917 46351 45951
rect 46293 45911 46351 45917
rect 25406 45880 25412 45892
rect 25367 45852 25412 45880
rect 25406 45840 25412 45852
rect 25464 45840 25470 45892
rect 41230 45880 41236 45892
rect 41191 45852 41236 45880
rect 41230 45840 41236 45852
rect 41288 45840 41294 45892
rect 44361 45883 44419 45889
rect 41386 45852 43576 45880
rect 24544 45784 24624 45812
rect 24544 45772 24550 45784
rect 38194 45772 38200 45824
rect 38252 45812 38258 45824
rect 41386 45812 41414 45852
rect 43438 45812 43444 45824
rect 38252 45784 41414 45812
rect 43399 45784 43444 45812
rect 38252 45772 38258 45784
rect 43438 45772 43444 45784
rect 43496 45772 43502 45824
rect 43548 45812 43576 45852
rect 44361 45849 44373 45883
rect 44407 45880 44419 45883
rect 46477 45883 46535 45889
rect 46477 45880 46489 45883
rect 44407 45852 46489 45880
rect 44407 45849 44419 45852
rect 44361 45843 44419 45849
rect 46477 45849 46489 45852
rect 46523 45849 46535 45883
rect 46477 45843 46535 45849
rect 45462 45812 45468 45824
rect 43548 45784 45468 45812
rect 45462 45772 45468 45784
rect 45520 45772 45526 45824
rect 45741 45815 45799 45821
rect 45741 45781 45753 45815
rect 45787 45812 45799 45815
rect 46014 45812 46020 45824
rect 45787 45784 46020 45812
rect 45787 45781 45799 45784
rect 45741 45775 45799 45781
rect 46014 45772 46020 45784
rect 46072 45772 46078 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 11882 45608 11888 45620
rect 11843 45580 11888 45608
rect 11882 45568 11888 45580
rect 11940 45568 11946 45620
rect 20990 45608 20996 45620
rect 20951 45580 20996 45608
rect 20990 45568 20996 45580
rect 21048 45568 21054 45620
rect 32398 45568 32404 45620
rect 32456 45608 32462 45620
rect 33045 45611 33103 45617
rect 33045 45608 33057 45611
rect 32456 45580 33057 45608
rect 32456 45568 32462 45580
rect 33045 45577 33057 45580
rect 33091 45577 33103 45611
rect 33045 45571 33103 45577
rect 40405 45611 40463 45617
rect 40405 45577 40417 45611
rect 40451 45608 40463 45611
rect 41230 45608 41236 45620
rect 40451 45580 41236 45608
rect 40451 45577 40463 45580
rect 40405 45571 40463 45577
rect 41230 45568 41236 45580
rect 41288 45568 41294 45620
rect 41417 45611 41475 45617
rect 41417 45577 41429 45611
rect 41463 45608 41475 45611
rect 42610 45608 42616 45620
rect 41463 45580 42616 45608
rect 41463 45577 41475 45580
rect 41417 45571 41475 45577
rect 42610 45568 42616 45580
rect 42668 45568 42674 45620
rect 46382 45568 46388 45620
rect 46440 45608 46446 45620
rect 46440 45580 47992 45608
rect 46440 45568 46446 45580
rect 42889 45543 42947 45549
rect 42889 45509 42901 45543
rect 42935 45540 42947 45543
rect 43438 45540 43444 45552
rect 42935 45512 43444 45540
rect 42935 45509 42947 45512
rect 42889 45503 42947 45509
rect 43438 45500 43444 45512
rect 43496 45500 43502 45552
rect 44818 45500 44824 45552
rect 44876 45540 44882 45552
rect 47964 45549 47992 45580
rect 47949 45543 48007 45549
rect 44876 45512 46428 45540
rect 44876 45500 44882 45512
rect 1762 45472 1768 45484
rect 1723 45444 1768 45472
rect 1762 45432 1768 45444
rect 1820 45432 1826 45484
rect 11793 45475 11851 45481
rect 11793 45441 11805 45475
rect 11839 45472 11851 45475
rect 20898 45472 20904 45484
rect 11839 45444 20904 45472
rect 11839 45441 11851 45444
rect 11793 45435 11851 45441
rect 20898 45432 20904 45444
rect 20956 45432 20962 45484
rect 25222 45432 25228 45484
rect 25280 45472 25286 45484
rect 25501 45475 25559 45481
rect 25501 45472 25513 45475
rect 25280 45444 25513 45472
rect 25280 45432 25286 45444
rect 25501 45441 25513 45444
rect 25547 45441 25559 45475
rect 25501 45435 25559 45441
rect 32953 45475 33011 45481
rect 32953 45441 32965 45475
rect 32999 45472 33011 45475
rect 38746 45472 38752 45484
rect 32999 45444 38752 45472
rect 32999 45441 33011 45444
rect 32953 45435 33011 45441
rect 38746 45432 38752 45444
rect 38804 45432 38810 45484
rect 40218 45432 40224 45484
rect 40276 45472 40282 45484
rect 40313 45475 40371 45481
rect 40313 45472 40325 45475
rect 40276 45444 40325 45472
rect 40276 45432 40282 45444
rect 40313 45441 40325 45444
rect 40359 45441 40371 45475
rect 40313 45435 40371 45441
rect 41325 45475 41383 45481
rect 41325 45441 41337 45475
rect 41371 45441 41383 45475
rect 42702 45472 42708 45484
rect 42663 45444 42708 45472
rect 41325 45435 41383 45441
rect 1949 45407 2007 45413
rect 1949 45373 1961 45407
rect 1995 45404 2007 45407
rect 2314 45404 2320 45416
rect 1995 45376 2320 45404
rect 1995 45373 2007 45376
rect 1949 45367 2007 45373
rect 2314 45364 2320 45376
rect 2372 45364 2378 45416
rect 2774 45404 2780 45416
rect 2735 45376 2780 45404
rect 2774 45364 2780 45376
rect 2832 45364 2838 45416
rect 41340 45268 41368 45435
rect 42702 45432 42708 45444
rect 42760 45432 42766 45484
rect 46400 45472 46428 45512
rect 47949 45509 47961 45543
rect 47995 45509 48007 45543
rect 47949 45503 48007 45509
rect 48133 45475 48191 45481
rect 48133 45472 48145 45475
rect 46400 45444 48145 45472
rect 48133 45441 48145 45444
rect 48179 45441 48191 45475
rect 48133 45435 48191 45441
rect 43162 45404 43168 45416
rect 43123 45376 43168 45404
rect 43162 45364 43168 45376
rect 43220 45364 43226 45416
rect 45002 45404 45008 45416
rect 44963 45376 45008 45404
rect 45002 45364 45008 45376
rect 45060 45364 45066 45416
rect 45189 45407 45247 45413
rect 45189 45373 45201 45407
rect 45235 45373 45247 45407
rect 45554 45404 45560 45416
rect 45515 45376 45560 45404
rect 45189 45367 45247 45373
rect 43254 45296 43260 45348
rect 43312 45336 43318 45348
rect 45204 45336 45232 45367
rect 45554 45364 45560 45376
rect 45612 45364 45618 45416
rect 43312 45308 45232 45336
rect 43312 45296 43318 45308
rect 46750 45268 46756 45280
rect 41340 45240 46756 45268
rect 46750 45228 46756 45240
rect 46808 45228 46814 45280
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 2314 45064 2320 45076
rect 2275 45036 2320 45064
rect 2314 45024 2320 45036
rect 2372 45024 2378 45076
rect 25406 45064 25412 45076
rect 25367 45036 25412 45064
rect 25406 45024 25412 45036
rect 25464 45024 25470 45076
rect 43254 45064 43260 45076
rect 43215 45036 43260 45064
rect 43254 45024 43260 45036
rect 43312 45024 43318 45076
rect 44085 45067 44143 45073
rect 44085 45033 44097 45067
rect 44131 45064 44143 45067
rect 45002 45064 45008 45076
rect 44131 45036 45008 45064
rect 44131 45033 44143 45036
rect 44085 45027 44143 45033
rect 45002 45024 45008 45036
rect 45060 45024 45066 45076
rect 45186 45064 45192 45076
rect 45147 45036 45192 45064
rect 45186 45024 45192 45036
rect 45244 45024 45250 45076
rect 45646 45024 45652 45076
rect 45704 45064 45710 45076
rect 45741 45067 45799 45073
rect 45741 45064 45753 45067
rect 45704 45036 45753 45064
rect 45704 45024 45710 45036
rect 45741 45033 45753 45036
rect 45787 45033 45799 45067
rect 45741 45027 45799 45033
rect 46293 44931 46351 44937
rect 46293 44897 46305 44931
rect 46339 44928 46351 44931
rect 47026 44928 47032 44940
rect 46339 44900 47032 44928
rect 46339 44897 46351 44900
rect 46293 44891 46351 44897
rect 47026 44888 47032 44900
rect 47084 44888 47090 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 2225 44863 2283 44869
rect 2225 44829 2237 44863
rect 2271 44860 2283 44863
rect 3786 44860 3792 44872
rect 2271 44832 3792 44860
rect 2271 44829 2283 44832
rect 2225 44823 2283 44829
rect 3786 44820 3792 44832
rect 3844 44820 3850 44872
rect 25314 44860 25320 44872
rect 25275 44832 25320 44860
rect 25314 44820 25320 44832
rect 25372 44820 25378 44872
rect 43162 44860 43168 44872
rect 43123 44832 43168 44860
rect 43162 44820 43168 44832
rect 43220 44820 43226 44872
rect 45554 44820 45560 44872
rect 45612 44860 45618 44872
rect 45649 44863 45707 44869
rect 45649 44860 45661 44863
rect 45612 44832 45661 44860
rect 45612 44820 45618 44832
rect 45649 44829 45661 44832
rect 45695 44829 45707 44863
rect 45649 44823 45707 44829
rect 46477 44795 46535 44801
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 47670 44792 47676 44804
rect 46523 44764 47676 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 47670 44752 47676 44764
rect 47728 44752 47734 44804
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 45370 44480 45376 44532
rect 45428 44520 45434 44532
rect 46293 44523 46351 44529
rect 46293 44520 46305 44523
rect 45428 44492 46305 44520
rect 45428 44480 45434 44492
rect 46293 44489 46305 44492
rect 46339 44489 46351 44523
rect 47670 44520 47676 44532
rect 47631 44492 47676 44520
rect 46293 44483 46351 44489
rect 47670 44480 47676 44492
rect 47728 44480 47734 44532
rect 45094 44384 45100 44396
rect 45055 44356 45100 44384
rect 45094 44344 45100 44356
rect 45152 44344 45158 44396
rect 45741 44387 45799 44393
rect 45741 44353 45753 44387
rect 45787 44384 45799 44387
rect 45830 44384 45836 44396
rect 45787 44356 45836 44384
rect 45787 44353 45799 44356
rect 45741 44347 45799 44353
rect 45830 44344 45836 44356
rect 45888 44344 45894 44396
rect 46198 44384 46204 44396
rect 46159 44356 46204 44384
rect 46198 44344 46204 44356
rect 46256 44384 46262 44396
rect 46845 44387 46903 44393
rect 46845 44384 46857 44387
rect 46256 44356 46857 44384
rect 46256 44344 46262 44356
rect 46845 44353 46857 44356
rect 46891 44384 46903 44387
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 46891 44356 47593 44384
rect 46891 44353 46903 44356
rect 46845 44347 46903 44353
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 38654 44316 38660 44328
rect 38615 44288 38660 44316
rect 38654 44276 38660 44288
rect 38712 44276 38718 44328
rect 38838 44316 38844 44328
rect 38799 44288 38844 44316
rect 38838 44276 38844 44288
rect 38896 44276 38902 44328
rect 40034 44316 40040 44328
rect 39995 44288 40040 44316
rect 40034 44276 40040 44288
rect 40092 44276 40098 44328
rect 46934 44180 46940 44192
rect 46895 44152 46940 44180
rect 46934 44140 46940 44152
rect 46992 44140 46998 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 38838 43976 38844 43988
rect 38799 43948 38844 43976
rect 38838 43936 38844 43948
rect 38896 43936 38902 43988
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 46934 43840 46940 43852
rect 46523 43812 46940 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 46934 43800 46940 43812
rect 46992 43800 46998 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 25774 43732 25780 43784
rect 25832 43772 25838 43784
rect 26973 43775 27031 43781
rect 26973 43772 26985 43775
rect 25832 43744 26985 43772
rect 25832 43732 25838 43744
rect 26973 43741 26985 43744
rect 27019 43741 27031 43775
rect 38749 43775 38807 43781
rect 38749 43772 38761 43775
rect 26973 43735 27031 43741
rect 31726 43744 38761 43772
rect 25314 43664 25320 43716
rect 25372 43704 25378 43716
rect 31726 43704 31754 43744
rect 38749 43741 38761 43744
rect 38795 43772 38807 43775
rect 38930 43772 38936 43784
rect 38795 43744 38936 43772
rect 38795 43741 38807 43744
rect 38749 43735 38807 43741
rect 38930 43732 38936 43744
rect 38988 43732 38994 43784
rect 45833 43775 45891 43781
rect 45833 43741 45845 43775
rect 45879 43772 45891 43775
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 45879 43744 46305 43772
rect 45879 43741 45891 43744
rect 45833 43735 45891 43741
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 25372 43676 31754 43704
rect 25372 43664 25378 43676
rect 27065 43639 27123 43645
rect 27065 43605 27077 43639
rect 27111 43636 27123 43639
rect 38654 43636 38660 43648
rect 27111 43608 38660 43636
rect 27111 43605 27123 43608
rect 27065 43599 27123 43605
rect 38654 43596 38660 43608
rect 38712 43596 38718 43648
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 47026 43296 47032 43308
rect 46987 43268 47032 43296
rect 47026 43256 47032 43268
rect 47084 43256 47090 43308
rect 1670 43228 1676 43240
rect 1631 43200 1676 43228
rect 1670 43188 1676 43200
rect 1728 43188 1734 43240
rect 47762 43092 47768 43104
rect 47723 43064 47768 43092
rect 47762 43052 47768 43064
rect 47820 43052 47826 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46293 42755 46351 42761
rect 46293 42721 46305 42755
rect 46339 42752 46351 42755
rect 47762 42752 47768 42764
rect 46339 42724 47768 42752
rect 46339 42721 46351 42724
rect 46293 42715 46351 42721
rect 47762 42712 47768 42724
rect 47820 42712 47826 42764
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 46934 42616 46940 42628
rect 46523 42588 46940 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 46934 42576 46940 42588
rect 46992 42576 46998 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 46934 42344 46940 42356
rect 46895 42316 46940 42344
rect 46934 42304 46940 42316
rect 46992 42304 46998 42356
rect 46566 42168 46572 42220
rect 46624 42208 46630 42220
rect 46842 42208 46848 42220
rect 46624 42180 46848 42208
rect 46624 42168 46630 42180
rect 46842 42168 46848 42180
rect 46900 42168 46906 42220
rect 47578 42208 47584 42220
rect 47539 42180 47584 42208
rect 47578 42168 47584 42180
rect 47636 42168 47642 42220
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 46474 41964 46480 42016
rect 46532 42004 46538 42016
rect 47673 42007 47731 42013
rect 47673 42004 47685 42007
rect 46532 41976 47685 42004
rect 46532 41964 46538 41976
rect 47673 41973 47685 41976
rect 47719 41973 47731 42007
rect 47673 41967 47731 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46474 41664 46480 41676
rect 46435 41636 46480 41664
rect 46474 41624 46480 41636
rect 46532 41624 46538 41676
rect 46293 41599 46351 41605
rect 46293 41565 46305 41599
rect 46339 41565 46351 41599
rect 48130 41596 48136 41608
rect 48091 41568 48136 41596
rect 46293 41559 46351 41565
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46308 41528 46336 41559
rect 48130 41556 48136 41568
rect 48188 41556 48194 41608
rect 47670 41528 47676 41540
rect 46308 41500 47676 41528
rect 47670 41488 47676 41500
rect 47728 41488 47734 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2133 41259 2191 41265
rect 2133 41256 2145 41259
rect 1636 41228 2145 41256
rect 1636 41216 1642 41228
rect 2133 41225 2145 41228
rect 2179 41225 2191 41259
rect 2133 41219 2191 41225
rect 2041 41123 2099 41129
rect 2041 41089 2053 41123
rect 2087 41120 2099 41123
rect 14090 41120 14096 41132
rect 2087 41092 14096 41120
rect 2087 41089 2099 41092
rect 2041 41083 2099 41089
rect 14090 41080 14096 41092
rect 14148 41080 14154 41132
rect 47946 41120 47952 41132
rect 47907 41092 47952 41120
rect 47946 41080 47952 41092
rect 48004 41080 48010 41132
rect 47486 40876 47492 40928
rect 47544 40916 47550 40928
rect 48041 40919 48099 40925
rect 48041 40916 48053 40919
rect 47544 40888 48053 40916
rect 47544 40876 47550 40888
rect 48041 40885 48053 40888
rect 48087 40885 48099 40919
rect 48041 40879 48099 40885
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 47670 40712 47676 40724
rect 47631 40684 47676 40712
rect 47670 40672 47676 40684
rect 47728 40672 47734 40724
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 1946 40372 1952 40384
rect 1907 40344 1952 40372
rect 1946 40332 1952 40344
rect 2004 40332 2010 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 46750 40032 46756 40044
rect 46711 40004 46756 40032
rect 46750 39992 46756 40004
rect 46808 39992 46814 40044
rect 46474 39788 46480 39840
rect 46532 39828 46538 39840
rect 46845 39831 46903 39837
rect 46845 39828 46857 39831
rect 46532 39800 46857 39828
rect 46532 39788 46538 39800
rect 46845 39797 46857 39800
rect 46891 39797 46903 39831
rect 47762 39828 47768 39840
rect 47723 39800 47768 39828
rect 46845 39791 46903 39797
rect 47762 39788 47768 39800
rect 47820 39788 47826 39840
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 47762 39556 47768 39568
rect 46308 39528 47768 39556
rect 20346 39448 20352 39500
rect 20404 39488 20410 39500
rect 46308 39497 46336 39528
rect 47762 39516 47768 39528
rect 47820 39516 47826 39568
rect 24949 39491 25007 39497
rect 24949 39488 24961 39491
rect 20404 39460 24961 39488
rect 20404 39448 20410 39460
rect 24949 39457 24961 39460
rect 24995 39457 25007 39491
rect 24949 39451 25007 39457
rect 46293 39491 46351 39497
rect 46293 39457 46305 39491
rect 46339 39457 46351 39491
rect 46474 39488 46480 39500
rect 46435 39460 46480 39488
rect 46293 39451 46351 39457
rect 46474 39448 46480 39460
rect 46532 39448 46538 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 22833 39423 22891 39429
rect 22833 39389 22845 39423
rect 22879 39420 22891 39423
rect 22879 39392 24440 39420
rect 22879 39389 22891 39392
rect 22833 39383 22891 39389
rect 22094 39244 22100 39296
rect 22152 39284 22158 39296
rect 24412 39293 24440 39392
rect 24578 39312 24584 39364
rect 24636 39352 24642 39364
rect 24857 39355 24915 39361
rect 24857 39352 24869 39355
rect 24636 39324 24869 39352
rect 24636 39312 24642 39324
rect 24857 39321 24869 39324
rect 24903 39321 24915 39355
rect 24857 39315 24915 39321
rect 22649 39287 22707 39293
rect 22649 39284 22661 39287
rect 22152 39256 22661 39284
rect 22152 39244 22158 39256
rect 22649 39253 22661 39256
rect 22695 39253 22707 39287
rect 22649 39247 22707 39253
rect 24397 39287 24455 39293
rect 24397 39253 24409 39287
rect 24443 39253 24455 39287
rect 24397 39247 24455 39253
rect 24765 39287 24823 39293
rect 24765 39253 24777 39287
rect 24811 39284 24823 39287
rect 25501 39287 25559 39293
rect 25501 39284 25513 39287
rect 24811 39256 25513 39284
rect 24811 39253 24823 39256
rect 24765 39247 24823 39253
rect 25501 39253 25513 39256
rect 25547 39284 25559 39287
rect 46014 39284 46020 39296
rect 25547 39256 46020 39284
rect 25547 39253 25559 39256
rect 25501 39247 25559 39253
rect 46014 39244 46020 39256
rect 46072 39244 46078 39296
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 24578 39080 24584 39092
rect 24539 39052 24584 39080
rect 24578 39040 24584 39052
rect 24636 39040 24642 39092
rect 19797 39015 19855 39021
rect 19797 38981 19809 39015
rect 19843 39012 19855 39015
rect 20806 39012 20812 39024
rect 19843 38984 20812 39012
rect 19843 38981 19855 38984
rect 19797 38975 19855 38981
rect 20806 38972 20812 38984
rect 20864 38972 20870 39024
rect 22094 38972 22100 39024
rect 22152 39012 22158 39024
rect 22152 38984 22197 39012
rect 22152 38972 22158 38984
rect 22554 38972 22560 39024
rect 22612 38972 22618 39024
rect 38749 39015 38807 39021
rect 38749 38981 38761 39015
rect 38795 39012 38807 39015
rect 38795 38984 39804 39012
rect 38795 38981 38807 38984
rect 38749 38975 38807 38981
rect 19981 38947 20039 38953
rect 19981 38913 19993 38947
rect 20027 38944 20039 38947
rect 20346 38944 20352 38956
rect 20027 38916 20352 38944
rect 20027 38913 20039 38916
rect 19981 38907 20039 38913
rect 20346 38904 20352 38916
rect 20404 38904 20410 38956
rect 24213 38947 24271 38953
rect 24213 38944 24225 38947
rect 23584 38916 24225 38944
rect 20530 38836 20536 38888
rect 20588 38876 20594 38888
rect 23584 38885 23612 38916
rect 24213 38913 24225 38916
rect 24259 38944 24271 38947
rect 24670 38944 24676 38956
rect 24259 38916 24676 38944
rect 24259 38913 24271 38916
rect 24213 38907 24271 38913
rect 24670 38904 24676 38916
rect 24728 38904 24734 38956
rect 39485 38947 39543 38953
rect 39485 38944 39497 38947
rect 38856 38916 39497 38944
rect 21821 38879 21879 38885
rect 21821 38876 21833 38879
rect 20588 38848 21833 38876
rect 20588 38836 20594 38848
rect 21821 38845 21833 38848
rect 21867 38845 21879 38879
rect 21821 38839 21879 38845
rect 23569 38879 23627 38885
rect 23569 38845 23581 38879
rect 23615 38845 23627 38879
rect 24118 38876 24124 38888
rect 24079 38848 24124 38876
rect 23569 38839 23627 38845
rect 24118 38836 24124 38848
rect 24176 38836 24182 38888
rect 19058 38700 19064 38752
rect 19116 38740 19122 38752
rect 20165 38743 20223 38749
rect 20165 38740 20177 38743
rect 19116 38712 20177 38740
rect 19116 38700 19122 38712
rect 20165 38709 20177 38712
rect 20211 38709 20223 38743
rect 20165 38703 20223 38709
rect 38654 38700 38660 38752
rect 38712 38740 38718 38752
rect 38856 38749 38884 38916
rect 39485 38913 39497 38916
rect 39531 38913 39543 38947
rect 39485 38907 39543 38913
rect 39776 38808 39804 38984
rect 47854 38944 47860 38956
rect 47815 38916 47860 38944
rect 47854 38904 47860 38916
rect 47912 38904 47918 38956
rect 39850 38836 39856 38888
rect 39908 38876 39914 38888
rect 39945 38879 40003 38885
rect 39945 38876 39957 38879
rect 39908 38848 39957 38876
rect 39908 38836 39914 38848
rect 39945 38845 39957 38848
rect 39991 38876 40003 38879
rect 46198 38876 46204 38888
rect 39991 38848 46204 38876
rect 39991 38845 40003 38848
rect 39945 38839 40003 38845
rect 46198 38836 46204 38848
rect 46256 38836 46262 38888
rect 41138 38808 41144 38820
rect 39776 38780 41144 38808
rect 41138 38768 41144 38780
rect 41196 38808 41202 38820
rect 48041 38811 48099 38817
rect 48041 38808 48053 38811
rect 41196 38780 48053 38808
rect 41196 38768 41202 38780
rect 48041 38777 48053 38780
rect 48087 38777 48099 38811
rect 48041 38771 48099 38777
rect 38841 38743 38899 38749
rect 38841 38740 38853 38743
rect 38712 38712 38853 38740
rect 38712 38700 38718 38712
rect 38841 38709 38853 38712
rect 38887 38709 38899 38743
rect 38841 38703 38899 38709
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 21358 38536 21364 38548
rect 12406 38508 21364 38536
rect 9490 38360 9496 38412
rect 9548 38400 9554 38412
rect 12406 38400 12434 38508
rect 21358 38496 21364 38508
rect 21416 38496 21422 38548
rect 21545 38539 21603 38545
rect 21545 38505 21557 38539
rect 21591 38536 21603 38539
rect 22554 38536 22560 38548
rect 21591 38508 22560 38536
rect 21591 38505 21603 38508
rect 21545 38499 21603 38505
rect 22554 38496 22560 38508
rect 22612 38496 22618 38548
rect 38930 38496 38936 38548
rect 38988 38536 38994 38548
rect 46750 38536 46756 38548
rect 38988 38508 46756 38536
rect 38988 38496 38994 38508
rect 46750 38496 46756 38508
rect 46808 38496 46814 38548
rect 18138 38428 18144 38480
rect 18196 38468 18202 38480
rect 23477 38471 23535 38477
rect 18196 38440 20760 38468
rect 18196 38428 18202 38440
rect 9548 38372 12434 38400
rect 9548 38360 9554 38372
rect 19242 38332 19248 38344
rect 19203 38304 19248 38332
rect 19242 38292 19248 38304
rect 19300 38292 19306 38344
rect 20732 38341 20760 38440
rect 23477 38437 23489 38471
rect 23523 38468 23535 38471
rect 23523 38440 24440 38468
rect 23523 38437 23535 38440
rect 23477 38431 23535 38437
rect 24412 38400 24440 38440
rect 26970 38400 26976 38412
rect 24412 38372 26976 38400
rect 19429 38335 19487 38341
rect 19429 38301 19441 38335
rect 19475 38301 19487 38335
rect 19429 38295 19487 38301
rect 20717 38335 20775 38341
rect 20717 38301 20729 38335
rect 20763 38332 20775 38335
rect 21453 38335 21511 38341
rect 21453 38332 21465 38335
rect 20763 38304 21465 38332
rect 20763 38301 20775 38304
rect 20717 38295 20775 38301
rect 21453 38301 21465 38304
rect 21499 38301 21511 38335
rect 21453 38295 21511 38301
rect 19444 38264 19472 38295
rect 22830 38292 22836 38344
rect 22888 38332 22894 38344
rect 24412 38341 24440 38372
rect 26970 38360 26976 38372
rect 27028 38360 27034 38412
rect 40678 38400 40684 38412
rect 40591 38372 40684 38400
rect 40678 38360 40684 38372
rect 40736 38400 40742 38412
rect 43162 38400 43168 38412
rect 40736 38372 43168 38400
rect 40736 38360 40742 38372
rect 43162 38360 43168 38372
rect 43220 38360 43226 38412
rect 23293 38335 23351 38341
rect 23293 38332 23305 38335
rect 22888 38304 23305 38332
rect 22888 38292 22894 38304
rect 23293 38301 23305 38304
rect 23339 38301 23351 38335
rect 23293 38295 23351 38301
rect 24397 38335 24455 38341
rect 24397 38301 24409 38335
rect 24443 38301 24455 38335
rect 24397 38295 24455 38301
rect 24486 38292 24492 38344
rect 24544 38292 24550 38344
rect 38654 38332 38660 38344
rect 38615 38304 38660 38332
rect 38654 38292 38660 38304
rect 38712 38332 38718 38344
rect 39853 38335 39911 38341
rect 39853 38332 39865 38335
rect 38712 38304 39865 38332
rect 38712 38292 38718 38304
rect 39853 38301 39865 38304
rect 39899 38301 39911 38335
rect 46290 38332 46296 38344
rect 46251 38304 46296 38332
rect 39853 38295 39911 38301
rect 46290 38292 46296 38304
rect 46348 38292 46354 38344
rect 23198 38264 23204 38276
rect 19444 38236 23204 38264
rect 23198 38224 23204 38236
rect 23256 38224 23262 38276
rect 24504 38264 24532 38292
rect 39209 38267 39267 38273
rect 39209 38264 39221 38267
rect 24504 38236 39221 38264
rect 39209 38233 39221 38236
rect 39255 38233 39267 38267
rect 39209 38227 39267 38233
rect 46477 38267 46535 38273
rect 46477 38233 46489 38267
rect 46523 38264 46535 38267
rect 46842 38264 46848 38276
rect 46523 38236 46848 38264
rect 46523 38233 46535 38236
rect 46477 38227 46535 38233
rect 19334 38196 19340 38208
rect 19295 38168 19340 38196
rect 19334 38156 19340 38168
rect 19392 38156 19398 38208
rect 20806 38196 20812 38208
rect 20767 38168 20812 38196
rect 20806 38156 20812 38168
rect 20864 38156 20870 38208
rect 24486 38196 24492 38208
rect 24447 38168 24492 38196
rect 24486 38156 24492 38168
rect 24544 38156 24550 38208
rect 39224 38196 39252 38227
rect 46842 38224 46848 38236
rect 46900 38224 46906 38276
rect 48130 38264 48136 38276
rect 48091 38236 48136 38264
rect 48130 38224 48136 38236
rect 48188 38224 48194 38276
rect 47302 38196 47308 38208
rect 39224 38168 47308 38196
rect 47302 38156 47308 38168
rect 47360 38196 47366 38208
rect 47578 38196 47584 38208
rect 47360 38168 47584 38196
rect 47360 38156 47366 38168
rect 47578 38156 47584 38168
rect 47636 38156 47642 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 22370 37992 22376 38004
rect 17972 37964 22376 37992
rect 17218 37816 17224 37868
rect 17276 37856 17282 37868
rect 17972 37865 18000 37964
rect 22370 37952 22376 37964
rect 22428 37952 22434 38004
rect 46842 37992 46848 38004
rect 22480 37964 24716 37992
rect 46803 37964 46848 37992
rect 19794 37924 19800 37936
rect 19755 37896 19800 37924
rect 19794 37884 19800 37896
rect 19852 37884 19858 37936
rect 20806 37884 20812 37936
rect 20864 37884 20870 37936
rect 22480 37865 22508 37964
rect 24486 37924 24492 37936
rect 23966 37896 24492 37924
rect 24486 37884 24492 37896
rect 24544 37884 24550 37936
rect 24688 37865 24716 37964
rect 46842 37952 46848 37964
rect 46900 37952 46906 38004
rect 27065 37927 27123 37933
rect 27065 37924 27077 37927
rect 26174 37896 27077 37924
rect 27065 37893 27077 37896
rect 27111 37893 27123 37927
rect 38654 37924 38660 37936
rect 27065 37887 27123 37893
rect 38488 37896 38660 37924
rect 17957 37859 18015 37865
rect 17957 37856 17969 37859
rect 17276 37828 17969 37856
rect 17276 37816 17282 37828
rect 17957 37825 17969 37828
rect 18003 37825 18015 37859
rect 22465 37859 22523 37865
rect 22465 37856 22477 37859
rect 17957 37819 18015 37825
rect 22066 37828 22477 37856
rect 19426 37748 19432 37800
rect 19484 37788 19490 37800
rect 19521 37791 19579 37797
rect 19521 37788 19533 37791
rect 19484 37760 19533 37788
rect 19484 37748 19490 37760
rect 19521 37757 19533 37760
rect 19567 37788 19579 37791
rect 20530 37788 20536 37800
rect 19567 37760 20536 37788
rect 19567 37757 19579 37760
rect 19521 37751 19579 37757
rect 20530 37748 20536 37760
rect 20588 37788 20594 37800
rect 22066 37788 22094 37828
rect 22465 37825 22477 37828
rect 22511 37825 22523 37859
rect 22465 37819 22523 37825
rect 24673 37859 24731 37865
rect 24673 37825 24685 37859
rect 24719 37825 24731 37859
rect 26970 37856 26976 37868
rect 26883 37828 26976 37856
rect 24673 37819 24731 37825
rect 26970 37816 26976 37828
rect 27028 37856 27034 37868
rect 27617 37859 27675 37865
rect 27617 37856 27629 37859
rect 27028 37828 27629 37856
rect 27028 37816 27034 37828
rect 27617 37825 27629 37828
rect 27663 37856 27675 37859
rect 29365 37859 29423 37865
rect 29365 37856 29377 37859
rect 27663 37828 29377 37856
rect 27663 37825 27675 37828
rect 27617 37819 27675 37825
rect 29365 37825 29377 37828
rect 29411 37856 29423 37859
rect 30650 37856 30656 37868
rect 29411 37828 30656 37856
rect 29411 37825 29423 37828
rect 29365 37819 29423 37825
rect 30650 37816 30656 37828
rect 30708 37816 30714 37868
rect 38488 37865 38516 37896
rect 38654 37884 38660 37896
rect 38712 37924 38718 37936
rect 39393 37927 39451 37933
rect 39393 37924 39405 37927
rect 38712 37896 39405 37924
rect 38712 37884 38718 37896
rect 39393 37893 39405 37896
rect 39439 37893 39451 37927
rect 39393 37887 39451 37893
rect 39942 37884 39948 37936
rect 40000 37924 40006 37936
rect 40218 37924 40224 37936
rect 40000 37896 40224 37924
rect 40000 37884 40006 37896
rect 40218 37884 40224 37896
rect 40276 37884 40282 37936
rect 46290 37884 46296 37936
rect 46348 37924 46354 37936
rect 46348 37896 47808 37924
rect 46348 37884 46354 37896
rect 38473 37859 38531 37865
rect 38473 37825 38485 37859
rect 38519 37825 38531 37859
rect 38746 37856 38752 37868
rect 38707 37828 38752 37856
rect 38473 37819 38531 37825
rect 38746 37816 38752 37828
rect 38804 37816 38810 37868
rect 46750 37856 46756 37868
rect 46711 37828 46756 37856
rect 46750 37816 46756 37828
rect 46808 37816 46814 37868
rect 47780 37865 47808 37896
rect 47765 37859 47823 37865
rect 47765 37825 47777 37859
rect 47811 37825 47823 37859
rect 47765 37819 47823 37825
rect 22738 37788 22744 37800
rect 20588 37760 22094 37788
rect 22699 37760 22744 37788
rect 20588 37748 20594 37760
rect 22738 37748 22744 37760
rect 22796 37748 22802 37800
rect 24946 37788 24952 37800
rect 24907 37760 24952 37788
rect 24946 37748 24952 37760
rect 25004 37748 25010 37800
rect 18138 37652 18144 37664
rect 18099 37624 18144 37652
rect 18138 37612 18144 37624
rect 18196 37612 18202 37664
rect 21174 37612 21180 37664
rect 21232 37652 21238 37664
rect 21269 37655 21327 37661
rect 21269 37652 21281 37655
rect 21232 37624 21281 37652
rect 21232 37612 21238 37624
rect 21269 37621 21281 37624
rect 21315 37652 21327 37655
rect 22186 37652 22192 37664
rect 21315 37624 22192 37652
rect 21315 37621 21327 37624
rect 21269 37615 21327 37621
rect 22186 37612 22192 37624
rect 22244 37612 22250 37664
rect 22370 37612 22376 37664
rect 22428 37652 22434 37664
rect 22830 37652 22836 37664
rect 22428 37624 22836 37652
rect 22428 37612 22434 37624
rect 22830 37612 22836 37624
rect 22888 37612 22894 37664
rect 24213 37655 24271 37661
rect 24213 37621 24225 37655
rect 24259 37652 24271 37655
rect 24394 37652 24400 37664
rect 24259 37624 24400 37652
rect 24259 37621 24271 37624
rect 24213 37615 24271 37621
rect 24394 37612 24400 37624
rect 24452 37612 24458 37664
rect 25498 37612 25504 37664
rect 25556 37652 25562 37664
rect 26421 37655 26479 37661
rect 26421 37652 26433 37655
rect 25556 37624 26433 37652
rect 25556 37612 25562 37624
rect 26421 37621 26433 37624
rect 26467 37621 26479 37655
rect 26421 37615 26479 37621
rect 27614 37612 27620 37664
rect 27672 37652 27678 37664
rect 27709 37655 27767 37661
rect 27709 37652 27721 37655
rect 27672 37624 27721 37652
rect 27672 37612 27678 37624
rect 27709 37621 27721 37624
rect 27755 37621 27767 37655
rect 29454 37652 29460 37664
rect 29415 37624 29460 37652
rect 27709 37615 27767 37621
rect 29454 37612 29460 37624
rect 29512 37612 29518 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 18598 37448 18604 37460
rect 18559 37420 18604 37448
rect 18598 37408 18604 37420
rect 18656 37408 18662 37460
rect 19794 37408 19800 37460
rect 19852 37448 19858 37460
rect 21637 37451 21695 37457
rect 21637 37448 21649 37451
rect 19852 37420 21649 37448
rect 19852 37408 19858 37420
rect 21637 37417 21649 37420
rect 21683 37417 21695 37451
rect 21637 37411 21695 37417
rect 22738 37408 22744 37460
rect 22796 37448 22802 37460
rect 23385 37451 23443 37457
rect 23385 37448 23397 37451
rect 22796 37420 23397 37448
rect 22796 37408 22802 37420
rect 23385 37417 23397 37420
rect 23431 37417 23443 37451
rect 24394 37448 24400 37460
rect 24355 37420 24400 37448
rect 23385 37411 23443 37417
rect 24394 37408 24400 37420
rect 24452 37408 24458 37460
rect 20162 37340 20168 37392
rect 20220 37380 20226 37392
rect 20220 37352 21312 37380
rect 20220 37340 20226 37352
rect 21174 37312 21180 37324
rect 21135 37284 21180 37312
rect 21174 37272 21180 37284
rect 21232 37272 21238 37324
rect 21284 37321 21312 37352
rect 21358 37340 21364 37392
rect 21416 37380 21422 37392
rect 21416 37352 25360 37380
rect 21416 37340 21422 37352
rect 21269 37315 21327 37321
rect 21269 37281 21281 37315
rect 21315 37281 21327 37315
rect 23198 37312 23204 37324
rect 23159 37284 23204 37312
rect 21269 37275 21327 37281
rect 23198 37272 23204 37284
rect 23256 37272 23262 37324
rect 24581 37315 24639 37321
rect 24581 37281 24593 37315
rect 24627 37312 24639 37315
rect 25332 37312 25360 37352
rect 28629 37315 28687 37321
rect 28629 37312 28641 37315
rect 24627 37284 24808 37312
rect 25332 37284 28641 37312
rect 24627 37281 24639 37284
rect 24581 37275 24639 37281
rect 24780 37256 24808 37284
rect 28629 37281 28641 37284
rect 28675 37281 28687 37315
rect 28629 37275 28687 37281
rect 29549 37315 29607 37321
rect 29549 37281 29561 37315
rect 29595 37312 29607 37315
rect 29914 37312 29920 37324
rect 29595 37284 29920 37312
rect 29595 37281 29607 37284
rect 29549 37275 29607 37281
rect 29914 37272 29920 37284
rect 29972 37272 29978 37324
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 2041 37247 2099 37253
rect 2041 37244 2053 37247
rect 1820 37216 2053 37244
rect 1820 37204 1826 37216
rect 2041 37213 2053 37216
rect 2087 37213 2099 37247
rect 18322 37244 18328 37256
rect 18283 37216 18328 37244
rect 2041 37207 2099 37213
rect 18322 37204 18328 37216
rect 18380 37204 18386 37256
rect 18417 37247 18475 37253
rect 18417 37213 18429 37247
rect 18463 37213 18475 37247
rect 18690 37244 18696 37256
rect 18651 37216 18696 37244
rect 18417 37207 18475 37213
rect 18432 37176 18460 37207
rect 18690 37204 18696 37216
rect 18748 37204 18754 37256
rect 20901 37247 20959 37253
rect 20901 37213 20913 37247
rect 20947 37244 20959 37247
rect 20990 37244 20996 37256
rect 20947 37216 20996 37244
rect 20947 37213 20959 37216
rect 20901 37207 20959 37213
rect 20990 37204 20996 37216
rect 21048 37204 21054 37256
rect 21085 37247 21143 37253
rect 21085 37213 21097 37247
rect 21131 37213 21143 37247
rect 21085 37207 21143 37213
rect 21453 37247 21511 37253
rect 21453 37213 21465 37247
rect 21499 37244 21511 37247
rect 21910 37244 21916 37256
rect 21499 37216 21916 37244
rect 21499 37213 21511 37216
rect 21453 37207 21511 37213
rect 18598 37176 18604 37188
rect 18432 37148 18604 37176
rect 18598 37136 18604 37148
rect 18656 37136 18662 37188
rect 21100 37176 21128 37207
rect 21910 37204 21916 37216
rect 21968 37204 21974 37256
rect 23014 37244 23020 37256
rect 22975 37216 23020 37244
rect 23014 37204 23020 37216
rect 23072 37204 23078 37256
rect 23385 37247 23443 37253
rect 23385 37213 23397 37247
rect 23431 37213 23443 37247
rect 24670 37244 24676 37256
rect 24631 37216 24676 37244
rect 23385 37207 23443 37213
rect 22554 37176 22560 37188
rect 21100 37148 22560 37176
rect 22554 37136 22560 37148
rect 22612 37136 22618 37188
rect 23400 37176 23428 37207
rect 24670 37204 24676 37216
rect 24728 37204 24734 37256
rect 24762 37204 24768 37256
rect 24820 37204 24826 37256
rect 25961 37247 26019 37253
rect 25961 37213 25973 37247
rect 26007 37213 26019 37247
rect 25961 37207 26019 37213
rect 28353 37247 28411 37253
rect 28353 37213 28365 37247
rect 28399 37213 28411 37247
rect 28353 37207 28411 37213
rect 28445 37247 28503 37253
rect 28445 37213 28457 37247
rect 28491 37244 28503 37247
rect 28534 37244 28540 37256
rect 28491 37216 28540 37244
rect 28491 37213 28503 37216
rect 28445 37207 28503 37213
rect 22756 37148 23428 37176
rect 18141 37111 18199 37117
rect 18141 37077 18153 37111
rect 18187 37108 18199 37111
rect 18506 37108 18512 37120
rect 18187 37080 18512 37108
rect 18187 37077 18199 37080
rect 18141 37071 18199 37077
rect 18506 37068 18512 37080
rect 18564 37068 18570 37120
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 22756 37108 22784 37148
rect 24302 37136 24308 37188
rect 24360 37176 24366 37188
rect 24397 37179 24455 37185
rect 24397 37176 24409 37179
rect 24360 37148 24409 37176
rect 24360 37136 24366 37148
rect 24397 37145 24409 37148
rect 24443 37145 24455 37179
rect 24397 37139 24455 37145
rect 19392 37080 22784 37108
rect 23109 37111 23167 37117
rect 19392 37068 19398 37080
rect 23109 37077 23121 37111
rect 23155 37108 23167 37111
rect 24118 37108 24124 37120
rect 23155 37080 24124 37108
rect 23155 37077 23167 37080
rect 23109 37071 23167 37077
rect 24118 37068 24124 37080
rect 24176 37068 24182 37120
rect 24854 37108 24860 37120
rect 24815 37080 24860 37108
rect 24854 37068 24860 37080
rect 24912 37068 24918 37120
rect 25976 37108 26004 37207
rect 26234 37176 26240 37188
rect 26195 37148 26240 37176
rect 26234 37136 26240 37148
rect 26292 37136 26298 37188
rect 27614 37176 27620 37188
rect 27462 37148 27620 37176
rect 27614 37136 27620 37148
rect 27672 37136 27678 37188
rect 28368 37176 28396 37207
rect 28534 37204 28540 37216
rect 28592 37204 28598 37256
rect 28718 37244 28724 37256
rect 28679 37216 28724 37244
rect 28718 37204 28724 37216
rect 28776 37204 28782 37256
rect 29638 37204 29644 37256
rect 29696 37244 29702 37256
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 29696 37216 29745 37244
rect 29696 37204 29702 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 29917 37179 29975 37185
rect 29917 37176 29929 37179
rect 28368 37148 29929 37176
rect 29917 37145 29929 37148
rect 29963 37145 29975 37179
rect 29917 37139 29975 37145
rect 27522 37108 27528 37120
rect 25976 37080 27528 37108
rect 27522 37068 27528 37080
rect 27580 37068 27586 37120
rect 27706 37108 27712 37120
rect 27667 37080 27712 37108
rect 27706 37068 27712 37080
rect 27764 37068 27770 37120
rect 28169 37111 28227 37117
rect 28169 37077 28181 37111
rect 28215 37108 28227 37111
rect 28442 37108 28448 37120
rect 28215 37080 28448 37108
rect 28215 37077 28227 37080
rect 28169 37071 28227 37077
rect 28442 37068 28448 37080
rect 28500 37068 28506 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 26234 36904 26240 36916
rect 26195 36876 26240 36904
rect 26234 36864 26240 36876
rect 26292 36864 26298 36916
rect 28718 36904 28724 36916
rect 28276 36876 28724 36904
rect 17954 36796 17960 36848
rect 18012 36796 18018 36848
rect 21726 36836 21732 36848
rect 21022 36808 21732 36836
rect 21726 36796 21732 36808
rect 21784 36796 21790 36848
rect 21910 36796 21916 36848
rect 21968 36836 21974 36848
rect 28276 36836 28304 36876
rect 28718 36864 28724 36876
rect 28776 36864 28782 36916
rect 28442 36836 28448 36848
rect 21968 36808 28304 36836
rect 28403 36808 28448 36836
rect 21968 36796 21974 36808
rect 28442 36796 28448 36808
rect 28500 36796 28506 36848
rect 29454 36796 29460 36848
rect 29512 36796 29518 36848
rect 1762 36768 1768 36780
rect 1723 36740 1768 36768
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 24302 36728 24308 36780
rect 24360 36768 24366 36780
rect 25498 36768 25504 36780
rect 24360 36740 25504 36768
rect 24360 36728 24366 36740
rect 25498 36728 25504 36740
rect 25556 36768 25562 36780
rect 25593 36771 25651 36777
rect 25593 36768 25605 36771
rect 25556 36740 25605 36768
rect 25556 36728 25562 36740
rect 25593 36737 25605 36740
rect 25639 36737 25651 36771
rect 25593 36731 25651 36737
rect 26234 36728 26240 36780
rect 26292 36768 26298 36780
rect 26421 36771 26479 36777
rect 26421 36768 26433 36771
rect 26292 36740 26433 36768
rect 26292 36728 26298 36740
rect 26421 36737 26433 36740
rect 26467 36737 26479 36771
rect 26421 36731 26479 36737
rect 27522 36728 27528 36780
rect 27580 36768 27586 36780
rect 28169 36771 28227 36777
rect 28169 36768 28181 36771
rect 27580 36740 28181 36768
rect 27580 36728 27586 36740
rect 28169 36737 28181 36740
rect 28215 36737 28227 36771
rect 30650 36768 30656 36780
rect 30611 36740 30656 36768
rect 28169 36731 28227 36737
rect 30650 36728 30656 36740
rect 30708 36728 30714 36780
rect 1949 36703 2007 36709
rect 1949 36669 1961 36703
rect 1995 36700 2007 36703
rect 2222 36700 2228 36712
rect 1995 36672 2228 36700
rect 1995 36669 2007 36672
rect 1949 36663 2007 36669
rect 2222 36660 2228 36672
rect 2280 36660 2286 36712
rect 2774 36700 2780 36712
rect 2735 36672 2780 36700
rect 2774 36660 2780 36672
rect 2832 36660 2838 36712
rect 16666 36700 16672 36712
rect 16627 36672 16672 36700
rect 16666 36660 16672 36672
rect 16724 36660 16730 36712
rect 16945 36703 17003 36709
rect 16945 36669 16957 36703
rect 16991 36700 17003 36703
rect 18230 36700 18236 36712
rect 16991 36672 18236 36700
rect 16991 36669 17003 36672
rect 16945 36663 17003 36669
rect 18230 36660 18236 36672
rect 18288 36660 18294 36712
rect 19426 36700 19432 36712
rect 18340 36672 19432 36700
rect 16666 36524 16672 36576
rect 16724 36564 16730 36576
rect 18340 36564 18368 36672
rect 19426 36660 19432 36672
rect 19484 36700 19490 36712
rect 19521 36703 19579 36709
rect 19521 36700 19533 36703
rect 19484 36672 19533 36700
rect 19484 36660 19490 36672
rect 19521 36669 19533 36672
rect 19567 36669 19579 36703
rect 19794 36700 19800 36712
rect 19755 36672 19800 36700
rect 19521 36663 19579 36669
rect 19794 36660 19800 36672
rect 19852 36660 19858 36712
rect 16724 36536 18368 36564
rect 18417 36567 18475 36573
rect 16724 36524 16730 36536
rect 18417 36533 18429 36567
rect 18463 36564 18475 36567
rect 18598 36564 18604 36576
rect 18463 36536 18604 36564
rect 18463 36533 18475 36536
rect 18417 36527 18475 36533
rect 18598 36524 18604 36536
rect 18656 36524 18662 36576
rect 21266 36564 21272 36576
rect 21227 36536 21272 36564
rect 21266 36524 21272 36536
rect 21324 36524 21330 36576
rect 25590 36524 25596 36576
rect 25648 36564 25654 36576
rect 25685 36567 25743 36573
rect 25685 36564 25697 36567
rect 25648 36536 25697 36564
rect 25648 36524 25654 36536
rect 25685 36533 25697 36536
rect 25731 36533 25743 36567
rect 29914 36564 29920 36576
rect 29875 36536 29920 36564
rect 25685 36527 25743 36533
rect 29914 36524 29920 36536
rect 29972 36524 29978 36576
rect 30742 36564 30748 36576
rect 30703 36536 30748 36564
rect 30742 36524 30748 36536
rect 30800 36524 30806 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 2222 36360 2228 36372
rect 2183 36332 2228 36360
rect 2222 36320 2228 36332
rect 2280 36320 2286 36372
rect 17681 36363 17739 36369
rect 17681 36329 17693 36363
rect 17727 36360 17739 36363
rect 18601 36363 18659 36369
rect 18601 36360 18613 36363
rect 17727 36332 18613 36360
rect 17727 36329 17739 36332
rect 17681 36323 17739 36329
rect 18601 36329 18613 36332
rect 18647 36329 18659 36363
rect 18601 36323 18659 36329
rect 19794 36320 19800 36372
rect 19852 36360 19858 36372
rect 20717 36363 20775 36369
rect 20717 36360 20729 36363
rect 19852 36332 20729 36360
rect 19852 36320 19858 36332
rect 20717 36329 20729 36332
rect 20763 36329 20775 36363
rect 21726 36360 21732 36372
rect 21687 36332 21732 36360
rect 20717 36323 20775 36329
rect 21726 36320 21732 36332
rect 21784 36320 21790 36372
rect 23014 36320 23020 36372
rect 23072 36360 23078 36372
rect 23753 36363 23811 36369
rect 23753 36360 23765 36363
rect 23072 36332 23765 36360
rect 23072 36320 23078 36332
rect 23753 36329 23765 36332
rect 23799 36329 23811 36363
rect 23753 36323 23811 36329
rect 24946 36320 24952 36372
rect 25004 36360 25010 36372
rect 25225 36363 25283 36369
rect 25225 36360 25237 36363
rect 25004 36332 25237 36360
rect 25004 36320 25010 36332
rect 25225 36329 25237 36332
rect 25271 36329 25283 36363
rect 25225 36323 25283 36329
rect 28353 36363 28411 36369
rect 28353 36329 28365 36363
rect 28399 36360 28411 36363
rect 28534 36360 28540 36372
rect 28399 36332 28540 36360
rect 28399 36329 28411 36332
rect 28353 36323 28411 36329
rect 28534 36320 28540 36332
rect 28592 36320 28598 36372
rect 40678 36292 40684 36304
rect 6886 36264 40684 36292
rect 2133 36159 2191 36165
rect 2133 36125 2145 36159
rect 2179 36156 2191 36159
rect 2406 36156 2412 36168
rect 2179 36128 2412 36156
rect 2179 36125 2191 36128
rect 2133 36119 2191 36125
rect 2406 36116 2412 36128
rect 2464 36156 2470 36168
rect 6886 36156 6914 36264
rect 40678 36252 40684 36264
rect 40736 36252 40742 36304
rect 17494 36224 17500 36236
rect 17455 36196 17500 36224
rect 17494 36184 17500 36196
rect 17552 36184 17558 36236
rect 18230 36224 18236 36236
rect 18191 36196 18236 36224
rect 18230 36184 18236 36196
rect 18288 36184 18294 36236
rect 18598 36224 18604 36236
rect 18340 36196 18604 36224
rect 2464 36128 6914 36156
rect 17405 36159 17463 36165
rect 2464 36116 2470 36128
rect 17405 36125 17417 36159
rect 17451 36156 17463 36159
rect 18340 36156 18368 36196
rect 18598 36184 18604 36196
rect 18656 36184 18662 36236
rect 22646 36224 22652 36236
rect 20916 36196 22652 36224
rect 17451 36128 18368 36156
rect 18417 36159 18475 36165
rect 17451 36125 17463 36128
rect 17405 36119 17463 36125
rect 18417 36125 18429 36159
rect 18463 36156 18475 36159
rect 18506 36156 18512 36168
rect 18463 36128 18512 36156
rect 18463 36125 18475 36128
rect 18417 36119 18475 36125
rect 18506 36116 18512 36128
rect 18564 36116 18570 36168
rect 18693 36159 18751 36165
rect 18693 36125 18705 36159
rect 18739 36156 18751 36159
rect 19426 36156 19432 36168
rect 18739 36128 19432 36156
rect 18739 36125 18751 36128
rect 18693 36119 18751 36125
rect 19426 36116 19432 36128
rect 19484 36116 19490 36168
rect 20916 36165 20944 36196
rect 22646 36184 22652 36196
rect 22704 36184 22710 36236
rect 23845 36227 23903 36233
rect 23845 36193 23857 36227
rect 23891 36224 23903 36227
rect 24394 36224 24400 36236
rect 23891 36196 24400 36224
rect 23891 36193 23903 36196
rect 23845 36187 23903 36193
rect 24394 36184 24400 36196
rect 24452 36184 24458 36236
rect 26421 36227 26479 36233
rect 26421 36224 26433 36227
rect 25240 36196 26433 36224
rect 20901 36159 20959 36165
rect 20901 36125 20913 36159
rect 20947 36125 20959 36159
rect 21082 36156 21088 36168
rect 21043 36128 21088 36156
rect 20901 36119 20959 36125
rect 21082 36116 21088 36128
rect 21140 36116 21146 36168
rect 21177 36159 21235 36165
rect 21177 36125 21189 36159
rect 21223 36125 21235 36159
rect 21177 36119 21235 36125
rect 11974 36048 11980 36100
rect 12032 36088 12038 36100
rect 21192 36088 21220 36119
rect 21450 36116 21456 36168
rect 21508 36156 21514 36168
rect 21637 36159 21695 36165
rect 21637 36156 21649 36159
rect 21508 36128 21649 36156
rect 21508 36116 21514 36128
rect 21637 36125 21649 36128
rect 21683 36125 21695 36159
rect 21637 36119 21695 36125
rect 22373 36159 22431 36165
rect 22373 36125 22385 36159
rect 22419 36125 22431 36159
rect 22373 36119 22431 36125
rect 22388 36088 22416 36119
rect 23474 36116 23480 36168
rect 23532 36156 23538 36168
rect 23569 36159 23627 36165
rect 23569 36156 23581 36159
rect 23532 36128 23581 36156
rect 23532 36116 23538 36128
rect 23569 36125 23581 36128
rect 23615 36125 23627 36159
rect 23569 36119 23627 36125
rect 23661 36159 23719 36165
rect 23661 36125 23673 36159
rect 23707 36156 23719 36159
rect 24578 36156 24584 36168
rect 23707 36128 24584 36156
rect 23707 36125 23719 36128
rect 23661 36119 23719 36125
rect 24578 36116 24584 36128
rect 24636 36116 24642 36168
rect 25240 36088 25268 36196
rect 26421 36193 26433 36196
rect 26467 36224 26479 36227
rect 27338 36224 27344 36236
rect 26467 36196 27344 36224
rect 26467 36193 26479 36196
rect 26421 36187 26479 36193
rect 27338 36184 27344 36196
rect 27396 36184 27402 36236
rect 27430 36184 27436 36236
rect 27488 36224 27494 36236
rect 28905 36227 28963 36233
rect 28905 36224 28917 36227
rect 27488 36196 28917 36224
rect 27488 36184 27494 36196
rect 28905 36193 28917 36196
rect 28951 36193 28963 36227
rect 28905 36187 28963 36193
rect 25314 36116 25320 36168
rect 25372 36156 25378 36168
rect 25409 36159 25467 36165
rect 25409 36156 25421 36159
rect 25372 36128 25421 36156
rect 25372 36116 25378 36128
rect 25409 36125 25421 36128
rect 25455 36125 25467 36159
rect 25409 36119 25467 36125
rect 25498 36116 25504 36168
rect 25556 36156 25562 36168
rect 25593 36159 25651 36165
rect 25593 36156 25605 36159
rect 25556 36128 25605 36156
rect 25556 36116 25562 36128
rect 25593 36125 25605 36128
rect 25639 36125 25651 36159
rect 25593 36119 25651 36125
rect 25685 36159 25743 36165
rect 25685 36125 25697 36159
rect 25731 36125 25743 36159
rect 25685 36119 25743 36125
rect 12032 36060 21220 36088
rect 22066 36060 25268 36088
rect 25700 36088 25728 36119
rect 25958 36116 25964 36168
rect 26016 36156 26022 36168
rect 26145 36159 26203 36165
rect 26145 36156 26157 36159
rect 26016 36128 26157 36156
rect 26016 36116 26022 36128
rect 26145 36125 26157 36128
rect 26191 36125 26203 36159
rect 26145 36119 26203 36125
rect 26237 36159 26295 36165
rect 26237 36125 26249 36159
rect 26283 36156 26295 36159
rect 26694 36156 26700 36168
rect 26283 36128 26700 36156
rect 26283 36125 26295 36128
rect 26237 36119 26295 36125
rect 26694 36116 26700 36128
rect 26752 36116 26758 36168
rect 27890 36116 27896 36168
rect 27948 36156 27954 36168
rect 28478 36159 28536 36165
rect 28478 36156 28490 36159
rect 27948 36128 28490 36156
rect 27948 36116 27954 36128
rect 28478 36125 28490 36128
rect 28524 36125 28536 36159
rect 28478 36119 28536 36125
rect 28994 36116 29000 36168
rect 29052 36156 29058 36168
rect 29733 36159 29791 36165
rect 29733 36156 29745 36159
rect 29052 36128 29745 36156
rect 29052 36116 29058 36128
rect 29733 36125 29745 36128
rect 29779 36156 29791 36159
rect 29914 36156 29920 36168
rect 29779 36128 29920 36156
rect 29779 36125 29791 36128
rect 29733 36119 29791 36125
rect 29914 36116 29920 36128
rect 29972 36116 29978 36168
rect 26421 36091 26479 36097
rect 26421 36088 26433 36091
rect 25700 36060 26433 36088
rect 12032 36048 12038 36060
rect 18322 35980 18328 36032
rect 18380 36020 18386 36032
rect 22066 36020 22094 36060
rect 26421 36057 26433 36060
rect 26467 36057 26479 36091
rect 26421 36051 26479 36057
rect 29086 36048 29092 36100
rect 29144 36088 29150 36100
rect 29549 36091 29607 36097
rect 29549 36088 29561 36091
rect 29144 36060 29561 36088
rect 29144 36048 29150 36060
rect 29549 36057 29561 36060
rect 29595 36088 29607 36091
rect 29638 36088 29644 36100
rect 29595 36060 29644 36088
rect 29595 36057 29607 36060
rect 29549 36051 29607 36057
rect 29638 36048 29644 36060
rect 29696 36048 29702 36100
rect 22554 36020 22560 36032
rect 18380 35992 22094 36020
rect 22515 35992 22560 36020
rect 18380 35980 18386 35992
rect 22554 35980 22560 35992
rect 22612 35980 22618 36032
rect 26602 35980 26608 36032
rect 26660 36020 26666 36032
rect 27706 36020 27712 36032
rect 26660 35992 27712 36020
rect 26660 35980 26666 35992
rect 27706 35980 27712 35992
rect 27764 35980 27770 36032
rect 28537 36023 28595 36029
rect 28537 35989 28549 36023
rect 28583 36020 28595 36023
rect 29454 36020 29460 36032
rect 28583 35992 29460 36020
rect 28583 35989 28595 35992
rect 28537 35983 28595 35989
rect 29454 35980 29460 35992
rect 29512 36020 29518 36032
rect 29917 36023 29975 36029
rect 29917 36020 29929 36023
rect 29512 35992 29929 36020
rect 29512 35980 29518 35992
rect 29917 35989 29929 35992
rect 29963 35989 29975 36023
rect 29917 35983 29975 35989
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 17589 35819 17647 35825
rect 17589 35785 17601 35819
rect 17635 35816 17647 35819
rect 17954 35816 17960 35828
rect 17635 35788 17960 35816
rect 17635 35785 17647 35788
rect 17589 35779 17647 35785
rect 17954 35776 17960 35788
rect 18012 35776 18018 35828
rect 18690 35776 18696 35828
rect 18748 35816 18754 35828
rect 22646 35816 22652 35828
rect 18748 35788 22508 35816
rect 22607 35788 22652 35816
rect 18748 35776 18754 35788
rect 21266 35708 21272 35760
rect 21324 35748 21330 35760
rect 22373 35751 22431 35757
rect 22373 35748 22385 35751
rect 21324 35720 22385 35748
rect 21324 35708 21330 35720
rect 22373 35717 22385 35720
rect 22419 35717 22431 35751
rect 22480 35748 22508 35788
rect 22646 35776 22652 35788
rect 22704 35776 22710 35828
rect 24118 35776 24124 35828
rect 24176 35816 24182 35828
rect 24213 35819 24271 35825
rect 24213 35816 24225 35819
rect 24176 35788 24225 35816
rect 24176 35776 24182 35788
rect 24213 35785 24225 35788
rect 24259 35785 24271 35819
rect 24213 35779 24271 35785
rect 24486 35776 24492 35828
rect 24544 35816 24550 35828
rect 31018 35816 31024 35828
rect 24544 35788 31024 35816
rect 24544 35776 24550 35788
rect 31018 35776 31024 35788
rect 31076 35776 31082 35828
rect 23198 35748 23204 35760
rect 22480 35720 23204 35748
rect 22373 35711 22431 35717
rect 23198 35708 23204 35720
rect 23256 35748 23262 35760
rect 26786 35748 26792 35760
rect 23256 35720 26792 35748
rect 23256 35708 23262 35720
rect 26786 35708 26792 35720
rect 26844 35708 26850 35760
rect 27522 35708 27528 35760
rect 27580 35748 27586 35760
rect 27580 35720 29868 35748
rect 27580 35708 27586 35720
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 15930 35640 15936 35692
rect 15988 35680 15994 35692
rect 17497 35683 17555 35689
rect 17497 35680 17509 35683
rect 15988 35652 17509 35680
rect 15988 35640 15994 35652
rect 17497 35649 17509 35652
rect 17543 35680 17555 35683
rect 19334 35680 19340 35692
rect 17543 35652 19340 35680
rect 17543 35649 17555 35652
rect 17497 35643 17555 35649
rect 19334 35640 19340 35652
rect 19392 35640 19398 35692
rect 21818 35640 21824 35692
rect 21876 35680 21882 35692
rect 22097 35683 22155 35689
rect 22097 35680 22109 35683
rect 21876 35652 22109 35680
rect 21876 35640 21882 35652
rect 22097 35649 22109 35652
rect 22143 35649 22155 35683
rect 22097 35643 22155 35649
rect 22281 35683 22339 35689
rect 22281 35649 22293 35683
rect 22327 35649 22339 35683
rect 22281 35643 22339 35649
rect 22465 35683 22523 35689
rect 22465 35649 22477 35683
rect 22511 35680 22523 35683
rect 23474 35680 23480 35692
rect 22511 35652 23480 35680
rect 22511 35649 22523 35652
rect 22465 35643 22523 35649
rect 22002 35572 22008 35624
rect 22060 35612 22066 35624
rect 22296 35612 22324 35643
rect 23474 35640 23480 35652
rect 23532 35640 23538 35692
rect 24029 35683 24087 35689
rect 24029 35649 24041 35683
rect 24075 35649 24087 35683
rect 24394 35680 24400 35692
rect 24355 35652 24400 35680
rect 24029 35643 24087 35649
rect 22060 35584 22324 35612
rect 24044 35612 24072 35643
rect 24394 35640 24400 35652
rect 24452 35640 24458 35692
rect 24578 35680 24584 35692
rect 24539 35652 24584 35680
rect 24578 35640 24584 35652
rect 24636 35640 24642 35692
rect 26510 35640 26516 35692
rect 26568 35680 26574 35692
rect 27430 35680 27436 35692
rect 26568 35652 27436 35680
rect 26568 35640 26574 35652
rect 27430 35640 27436 35652
rect 27488 35640 27494 35692
rect 28166 35680 28172 35692
rect 28127 35652 28172 35680
rect 28166 35640 28172 35652
rect 28224 35640 28230 35692
rect 28905 35683 28963 35689
rect 28905 35680 28917 35683
rect 28368 35652 28917 35680
rect 24946 35612 24952 35624
rect 24044 35584 24952 35612
rect 22060 35572 22066 35584
rect 20530 35504 20536 35556
rect 20588 35544 20594 35556
rect 22296 35544 22324 35584
rect 24946 35572 24952 35584
rect 25004 35572 25010 35624
rect 25682 35612 25688 35624
rect 25643 35584 25688 35612
rect 25682 35572 25688 35584
rect 25740 35572 25746 35624
rect 26145 35615 26203 35621
rect 26145 35581 26157 35615
rect 26191 35612 26203 35615
rect 26234 35612 26240 35624
rect 26191 35584 26240 35612
rect 26191 35581 26203 35584
rect 26145 35575 26203 35581
rect 26234 35572 26240 35584
rect 26292 35572 26298 35624
rect 25314 35544 25320 35556
rect 20588 35516 22094 35544
rect 22296 35516 25320 35544
rect 20588 35504 20594 35516
rect 1397 35479 1455 35485
rect 1397 35445 1409 35479
rect 1443 35476 1455 35479
rect 2130 35476 2136 35488
rect 1443 35448 2136 35476
rect 1443 35445 1455 35448
rect 1397 35439 1455 35445
rect 2130 35436 2136 35448
rect 2188 35436 2194 35488
rect 22066 35476 22094 35516
rect 25314 35504 25320 35516
rect 25372 35504 25378 35556
rect 26053 35547 26111 35553
rect 26053 35513 26065 35547
rect 26099 35544 26111 35547
rect 26326 35544 26332 35556
rect 26099 35516 26332 35544
rect 26099 35513 26111 35516
rect 26053 35507 26111 35513
rect 26326 35504 26332 35516
rect 26384 35504 26390 35556
rect 27338 35504 27344 35556
rect 27396 35544 27402 35556
rect 28368 35553 28396 35652
rect 28905 35649 28917 35652
rect 28951 35649 28963 35683
rect 29086 35680 29092 35692
rect 29047 35652 29092 35680
rect 28905 35643 28963 35649
rect 29086 35640 29092 35652
rect 29144 35640 29150 35692
rect 29840 35689 29868 35720
rect 30742 35708 30748 35760
rect 30800 35708 30806 35760
rect 29825 35683 29883 35689
rect 29825 35649 29837 35683
rect 29871 35649 29883 35683
rect 48130 35680 48136 35692
rect 48091 35652 48136 35680
rect 29825 35643 29883 35649
rect 48130 35640 48136 35652
rect 48188 35640 48194 35692
rect 28445 35615 28503 35621
rect 28445 35581 28457 35615
rect 28491 35612 28503 35615
rect 28626 35612 28632 35624
rect 28491 35584 28632 35612
rect 28491 35581 28503 35584
rect 28445 35575 28503 35581
rect 28626 35572 28632 35584
rect 28684 35572 28690 35624
rect 30101 35615 30159 35621
rect 30101 35581 30113 35615
rect 30147 35612 30159 35615
rect 30742 35612 30748 35624
rect 30147 35584 30748 35612
rect 30147 35581 30159 35584
rect 30101 35575 30159 35581
rect 30742 35572 30748 35584
rect 30800 35572 30806 35624
rect 27617 35547 27675 35553
rect 27617 35544 27629 35547
rect 27396 35516 27629 35544
rect 27396 35504 27402 35516
rect 27617 35513 27629 35516
rect 27663 35513 27675 35547
rect 27617 35507 27675 35513
rect 28353 35547 28411 35553
rect 28353 35513 28365 35547
rect 28399 35513 28411 35547
rect 28353 35507 28411 35513
rect 24394 35476 24400 35488
rect 22066 35448 24400 35476
rect 24394 35436 24400 35448
rect 24452 35436 24458 35488
rect 24489 35479 24547 35485
rect 24489 35445 24501 35479
rect 24535 35476 24547 35479
rect 26142 35476 26148 35488
rect 24535 35448 26148 35476
rect 24535 35445 24547 35448
rect 24489 35439 24547 35445
rect 26142 35436 26148 35448
rect 26200 35436 26206 35488
rect 28258 35476 28264 35488
rect 28219 35448 28264 35476
rect 28258 35436 28264 35448
rect 28316 35436 28322 35488
rect 28442 35436 28448 35488
rect 28500 35476 28506 35488
rect 28997 35479 29055 35485
rect 28997 35476 29009 35479
rect 28500 35448 29009 35476
rect 28500 35436 28506 35448
rect 28997 35445 29009 35448
rect 29043 35445 29055 35479
rect 28997 35439 29055 35445
rect 30558 35436 30564 35488
rect 30616 35476 30622 35488
rect 31573 35479 31631 35485
rect 31573 35476 31585 35479
rect 30616 35448 31585 35476
rect 30616 35436 30622 35448
rect 31573 35445 31585 35448
rect 31619 35445 31631 35479
rect 31573 35439 31631 35445
rect 47118 35436 47124 35488
rect 47176 35476 47182 35488
rect 47949 35479 48007 35485
rect 47949 35476 47961 35479
rect 47176 35448 47961 35476
rect 47176 35436 47182 35448
rect 47949 35445 47961 35448
rect 47995 35445 48007 35479
rect 47949 35439 48007 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 21818 35272 21824 35284
rect 21779 35244 21824 35272
rect 21818 35232 21824 35244
rect 21876 35232 21882 35284
rect 26326 35272 26332 35284
rect 26287 35244 26332 35272
rect 26326 35232 26332 35244
rect 26384 35232 26390 35284
rect 27893 35275 27951 35281
rect 27893 35241 27905 35275
rect 27939 35272 27951 35275
rect 28442 35272 28448 35284
rect 27939 35244 28448 35272
rect 27939 35241 27951 35244
rect 27893 35235 27951 35241
rect 28442 35232 28448 35244
rect 28500 35232 28506 35284
rect 28813 35275 28871 35281
rect 28813 35241 28825 35275
rect 28859 35272 28871 35275
rect 28994 35272 29000 35284
rect 28859 35244 29000 35272
rect 28859 35241 28871 35244
rect 28813 35235 28871 35241
rect 28994 35232 29000 35244
rect 29052 35232 29058 35284
rect 30742 35232 30748 35284
rect 30800 35272 30806 35284
rect 31021 35275 31079 35281
rect 31021 35272 31033 35275
rect 30800 35244 31033 35272
rect 30800 35232 30806 35244
rect 31021 35241 31033 35244
rect 31067 35241 31079 35275
rect 31021 35235 31079 35241
rect 24762 35164 24768 35216
rect 24820 35204 24826 35216
rect 26602 35204 26608 35216
rect 24820 35176 26608 35204
rect 24820 35164 24826 35176
rect 17129 35139 17187 35145
rect 17129 35105 17141 35139
rect 17175 35136 17187 35139
rect 19426 35136 19432 35148
rect 17175 35108 19432 35136
rect 17175 35105 17187 35108
rect 17129 35099 17187 35105
rect 19426 35096 19432 35108
rect 19484 35136 19490 35148
rect 20162 35136 20168 35148
rect 19484 35108 20168 35136
rect 19484 35096 19490 35108
rect 20162 35096 20168 35108
rect 20220 35096 20226 35148
rect 21637 35139 21695 35145
rect 21637 35105 21649 35139
rect 21683 35136 21695 35139
rect 22094 35136 22100 35148
rect 21683 35108 22100 35136
rect 21683 35105 21695 35108
rect 21637 35099 21695 35105
rect 22094 35096 22100 35108
rect 22152 35096 22158 35148
rect 25240 35145 25268 35176
rect 26602 35164 26608 35176
rect 26660 35164 26666 35216
rect 28258 35164 28264 35216
rect 28316 35204 28322 35216
rect 28902 35204 28908 35216
rect 28316 35176 28908 35204
rect 28316 35164 28322 35176
rect 28902 35164 28908 35176
rect 28960 35164 28966 35216
rect 30009 35207 30067 35213
rect 30009 35173 30021 35207
rect 30055 35204 30067 35207
rect 30055 35176 30696 35204
rect 30055 35173 30067 35176
rect 30009 35167 30067 35173
rect 25225 35139 25283 35145
rect 25225 35105 25237 35139
rect 25271 35105 25283 35139
rect 25590 35136 25596 35148
rect 25551 35108 25596 35136
rect 25225 35099 25283 35105
rect 25590 35096 25596 35108
rect 25648 35096 25654 35148
rect 26789 35139 26847 35145
rect 26789 35105 26801 35139
rect 26835 35136 26847 35139
rect 27246 35136 27252 35148
rect 26835 35108 27252 35136
rect 26835 35105 26847 35108
rect 26789 35099 26847 35105
rect 27246 35096 27252 35108
rect 27304 35096 27310 35148
rect 28626 35136 28632 35148
rect 28587 35108 28632 35136
rect 28626 35096 28632 35108
rect 28684 35096 28690 35148
rect 30558 35136 30564 35148
rect 28828 35108 30564 35136
rect 16850 35068 16856 35080
rect 16811 35040 16856 35068
rect 16850 35028 16856 35040
rect 16908 35028 16914 35080
rect 17034 35068 17040 35080
rect 16995 35040 17040 35068
rect 17034 35028 17040 35040
rect 17092 35028 17098 35080
rect 19334 35068 19340 35080
rect 19247 35040 19340 35068
rect 19334 35028 19340 35040
rect 19392 35028 19398 35080
rect 20346 35028 20352 35080
rect 20404 35068 20410 35080
rect 20533 35071 20591 35077
rect 20533 35068 20545 35071
rect 20404 35040 20545 35068
rect 20404 35028 20410 35040
rect 20533 35037 20545 35040
rect 20579 35037 20591 35071
rect 20533 35031 20591 35037
rect 21266 35028 21272 35080
rect 21324 35068 21330 35080
rect 21545 35071 21603 35077
rect 21545 35068 21557 35071
rect 21324 35040 21557 35068
rect 21324 35028 21330 35040
rect 21545 35037 21557 35040
rect 21591 35037 21603 35071
rect 21545 35031 21603 35037
rect 24397 35071 24455 35077
rect 24397 35037 24409 35071
rect 24443 35068 24455 35071
rect 24854 35068 24860 35080
rect 24443 35040 24860 35068
rect 24443 35037 24455 35040
rect 24397 35031 24455 35037
rect 24854 35028 24860 35040
rect 24912 35028 24918 35080
rect 25130 35028 25136 35080
rect 25188 35068 25194 35080
rect 25685 35071 25743 35077
rect 25685 35068 25697 35071
rect 25188 35040 25697 35068
rect 25188 35028 25194 35040
rect 25685 35037 25697 35040
rect 25731 35068 25743 35071
rect 26326 35068 26332 35080
rect 25731 35040 26332 35068
rect 25731 35037 25743 35040
rect 25685 35031 25743 35037
rect 26326 35028 26332 35040
rect 26384 35028 26390 35080
rect 26510 35068 26516 35080
rect 26471 35040 26516 35068
rect 26510 35028 26516 35040
rect 26568 35028 26574 35080
rect 26602 35028 26608 35080
rect 26660 35068 26666 35080
rect 26878 35068 26884 35080
rect 26660 35040 26705 35068
rect 26839 35040 26884 35068
rect 26660 35028 26666 35040
rect 26878 35028 26884 35040
rect 26936 35028 26942 35080
rect 27706 35068 27712 35080
rect 27667 35040 27712 35068
rect 27706 35028 27712 35040
rect 27764 35028 27770 35080
rect 28828 35077 28856 35108
rect 30558 35096 30564 35108
rect 30616 35096 30622 35148
rect 30668 35145 30696 35176
rect 30653 35139 30711 35145
rect 30653 35105 30665 35139
rect 30699 35136 30711 35139
rect 30926 35136 30932 35148
rect 30699 35108 30932 35136
rect 30699 35105 30711 35108
rect 30653 35099 30711 35105
rect 30926 35096 30932 35108
rect 30984 35096 30990 35148
rect 27985 35071 28043 35077
rect 27985 35037 27997 35071
rect 28031 35068 28043 35071
rect 28813 35071 28871 35077
rect 28031 35040 28672 35068
rect 28031 35037 28043 35040
rect 27985 35031 28043 35037
rect 19352 35000 19380 35028
rect 20806 35000 20812 35012
rect 19352 34972 20812 35000
rect 20806 34960 20812 34972
rect 20864 35000 20870 35012
rect 21450 35000 21456 35012
rect 20864 34972 21456 35000
rect 20864 34960 20870 34972
rect 21450 34960 21456 34972
rect 21508 34960 21514 35012
rect 24026 34960 24032 35012
rect 24084 35000 24090 35012
rect 24581 35003 24639 35009
rect 24581 35000 24593 35003
rect 24084 34972 24593 35000
rect 24084 34960 24090 34972
rect 24581 34969 24593 34972
rect 24627 35000 24639 35003
rect 24627 34972 27660 35000
rect 24627 34969 24639 34972
rect 24581 34963 24639 34969
rect 16669 34935 16727 34941
rect 16669 34901 16681 34935
rect 16715 34932 16727 34935
rect 16758 34932 16764 34944
rect 16715 34904 16764 34932
rect 16715 34901 16727 34904
rect 16669 34895 16727 34901
rect 16758 34892 16764 34904
rect 16816 34892 16822 34944
rect 19426 34932 19432 34944
rect 19387 34904 19432 34932
rect 19426 34892 19432 34904
rect 19484 34892 19490 34944
rect 20530 34892 20536 34944
rect 20588 34932 20594 34944
rect 20717 34935 20775 34941
rect 20717 34932 20729 34935
rect 20588 34904 20729 34932
rect 20588 34892 20594 34904
rect 20717 34901 20729 34904
rect 20763 34901 20775 34935
rect 20717 34895 20775 34901
rect 22370 34892 22376 34944
rect 22428 34932 22434 34944
rect 24765 34935 24823 34941
rect 24765 34932 24777 34935
rect 22428 34904 24777 34932
rect 22428 34892 22434 34904
rect 24765 34901 24777 34904
rect 24811 34901 24823 34935
rect 25866 34932 25872 34944
rect 25827 34904 25872 34932
rect 24765 34895 24823 34901
rect 25866 34892 25872 34904
rect 25924 34892 25930 34944
rect 27430 34892 27436 34944
rect 27488 34932 27494 34944
rect 27525 34935 27583 34941
rect 27525 34932 27537 34935
rect 27488 34904 27537 34932
rect 27488 34892 27494 34904
rect 27525 34901 27537 34904
rect 27571 34901 27583 34935
rect 27632 34932 27660 34972
rect 28166 34960 28172 35012
rect 28224 35000 28230 35012
rect 28534 35000 28540 35012
rect 28224 34972 28540 35000
rect 28224 34960 28230 34972
rect 28534 34960 28540 34972
rect 28592 34960 28598 35012
rect 28644 35000 28672 35040
rect 28813 35037 28825 35071
rect 28859 35037 28871 35071
rect 28813 35031 28871 35037
rect 28994 35028 29000 35080
rect 29052 35028 29058 35080
rect 30282 35068 30288 35080
rect 30243 35040 30288 35068
rect 30282 35028 30288 35040
rect 30340 35028 30346 35080
rect 30469 35071 30527 35077
rect 30469 35037 30481 35071
rect 30515 35037 30527 35071
rect 30469 35031 30527 35037
rect 30837 35071 30895 35077
rect 30837 35037 30849 35071
rect 30883 35068 30895 35071
rect 31018 35068 31024 35080
rect 30883 35040 31024 35068
rect 30883 35037 30895 35040
rect 30837 35031 30895 35037
rect 29012 35000 29040 35028
rect 28644 34972 29040 35000
rect 29822 34960 29828 35012
rect 29880 35000 29886 35012
rect 30484 35000 30512 35031
rect 31018 35028 31024 35040
rect 31076 35028 31082 35080
rect 48133 35071 48191 35077
rect 48133 35037 48145 35071
rect 48179 35068 48191 35071
rect 48222 35068 48228 35080
rect 48179 35040 48228 35068
rect 48179 35037 48191 35040
rect 48133 35031 48191 35037
rect 48222 35028 48228 35040
rect 48280 35028 48286 35080
rect 29880 34972 30512 35000
rect 29880 34960 29886 34972
rect 28718 34932 28724 34944
rect 27632 34904 28724 34932
rect 27525 34895 27583 34901
rect 28718 34892 28724 34904
rect 28776 34932 28782 34944
rect 28997 34935 29055 34941
rect 28997 34932 29009 34935
rect 28776 34904 29009 34932
rect 28776 34892 28782 34904
rect 28997 34901 29009 34904
rect 29043 34901 29055 34935
rect 28997 34895 29055 34901
rect 47854 34892 47860 34944
rect 47912 34932 47918 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47912 34904 47961 34932
rect 47912 34892 47918 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 16850 34688 16856 34740
rect 16908 34728 16914 34740
rect 17221 34731 17279 34737
rect 17221 34728 17233 34731
rect 16908 34700 17233 34728
rect 16908 34688 16914 34700
rect 17221 34697 17233 34700
rect 17267 34697 17279 34731
rect 18322 34728 18328 34740
rect 17221 34691 17279 34697
rect 17420 34700 18328 34728
rect 15930 34592 15936 34604
rect 15891 34564 15936 34592
rect 15930 34552 15936 34564
rect 15988 34552 15994 34604
rect 17420 34601 17448 34700
rect 18322 34688 18328 34700
rect 18380 34688 18386 34740
rect 21082 34688 21088 34740
rect 21140 34728 21146 34740
rect 24394 34728 24400 34740
rect 21140 34700 24400 34728
rect 21140 34688 21146 34700
rect 24394 34688 24400 34700
rect 24452 34688 24458 34740
rect 24489 34731 24547 34737
rect 24489 34697 24501 34731
rect 24535 34728 24547 34731
rect 24578 34728 24584 34740
rect 24535 34700 24584 34728
rect 24535 34697 24547 34700
rect 24489 34691 24547 34697
rect 24578 34688 24584 34700
rect 24636 34688 24642 34740
rect 25041 34731 25099 34737
rect 25041 34697 25053 34731
rect 25087 34728 25099 34731
rect 25222 34728 25228 34740
rect 25087 34700 25228 34728
rect 25087 34697 25099 34700
rect 25041 34691 25099 34697
rect 25222 34688 25228 34700
rect 25280 34688 25286 34740
rect 25590 34688 25596 34740
rect 25648 34688 25654 34740
rect 27706 34728 27712 34740
rect 27667 34700 27712 34728
rect 27706 34688 27712 34700
rect 27764 34688 27770 34740
rect 29365 34731 29423 34737
rect 27816 34700 28856 34728
rect 18690 34660 18696 34672
rect 17788 34632 18696 34660
rect 17788 34601 17816 34632
rect 18690 34620 18696 34632
rect 18748 34620 18754 34672
rect 19426 34620 19432 34672
rect 19484 34620 19490 34672
rect 22094 34660 22100 34672
rect 22066 34620 22100 34660
rect 22152 34660 22158 34672
rect 23109 34663 23167 34669
rect 23109 34660 23121 34663
rect 22152 34632 23121 34660
rect 22152 34620 22158 34632
rect 23109 34629 23121 34632
rect 23155 34660 23167 34663
rect 23382 34660 23388 34672
rect 23155 34632 23388 34660
rect 23155 34629 23167 34632
rect 23109 34623 23167 34629
rect 23382 34620 23388 34632
rect 23440 34620 23446 34672
rect 24026 34660 24032 34672
rect 23987 34632 24032 34660
rect 24026 34620 24032 34632
rect 24084 34620 24090 34672
rect 25130 34620 25136 34672
rect 25188 34660 25194 34672
rect 25409 34663 25467 34669
rect 25188 34632 25268 34660
rect 25188 34620 25194 34632
rect 17405 34595 17463 34601
rect 17405 34561 17417 34595
rect 17451 34561 17463 34595
rect 17405 34555 17463 34561
rect 17497 34595 17555 34601
rect 17497 34561 17509 34595
rect 17543 34561 17555 34595
rect 17497 34555 17555 34561
rect 17773 34595 17831 34601
rect 17773 34561 17785 34595
rect 17819 34561 17831 34595
rect 20898 34592 20904 34604
rect 17773 34555 17831 34561
rect 20180 34564 20904 34592
rect 16025 34527 16083 34533
rect 16025 34493 16037 34527
rect 16071 34524 16083 34527
rect 16574 34524 16580 34536
rect 16071 34496 16580 34524
rect 16071 34493 16083 34496
rect 16025 34487 16083 34493
rect 16574 34484 16580 34496
rect 16632 34484 16638 34536
rect 17310 34484 17316 34536
rect 17368 34524 17374 34536
rect 17512 34524 17540 34555
rect 17368 34496 17540 34524
rect 17368 34484 17374 34496
rect 17586 34484 17592 34536
rect 17644 34524 17650 34536
rect 17681 34527 17739 34533
rect 17681 34524 17693 34527
rect 17644 34496 17693 34524
rect 17644 34484 17650 34496
rect 17681 34493 17693 34496
rect 17727 34493 17739 34527
rect 18414 34524 18420 34536
rect 18375 34496 18420 34524
rect 17681 34487 17739 34493
rect 18414 34484 18420 34496
rect 18472 34484 18478 34536
rect 20180 34533 20208 34564
rect 20898 34552 20904 34564
rect 20956 34552 20962 34604
rect 21085 34595 21143 34601
rect 21085 34561 21097 34595
rect 21131 34592 21143 34595
rect 22066 34592 22094 34620
rect 22186 34592 22192 34604
rect 21131 34564 22094 34592
rect 22147 34564 22192 34592
rect 21131 34561 21143 34564
rect 21085 34555 21143 34561
rect 22186 34552 22192 34564
rect 22244 34552 22250 34604
rect 22370 34592 22376 34604
rect 22331 34564 22376 34592
rect 22370 34552 22376 34564
rect 22428 34552 22434 34604
rect 22922 34592 22928 34604
rect 22883 34564 22928 34592
rect 22922 34552 22928 34564
rect 22980 34552 22986 34604
rect 23658 34592 23664 34604
rect 23216 34564 23664 34592
rect 20165 34527 20223 34533
rect 20165 34493 20177 34527
rect 20211 34493 20223 34527
rect 20165 34487 20223 34493
rect 21177 34527 21235 34533
rect 21177 34493 21189 34527
rect 21223 34524 21235 34527
rect 21266 34524 21272 34536
rect 21223 34496 21272 34524
rect 21223 34493 21235 34496
rect 21177 34487 21235 34493
rect 21266 34484 21272 34496
rect 21324 34484 21330 34536
rect 22465 34527 22523 34533
rect 22465 34493 22477 34527
rect 22511 34524 22523 34527
rect 23216 34524 23244 34564
rect 23658 34552 23664 34564
rect 23716 34552 23722 34604
rect 24305 34595 24363 34601
rect 24305 34561 24317 34595
rect 24351 34592 24363 34595
rect 24762 34592 24768 34604
rect 24351 34564 24768 34592
rect 24351 34561 24363 34564
rect 24305 34555 24363 34561
rect 24762 34552 24768 34564
rect 24820 34552 24826 34604
rect 25240 34601 25268 34632
rect 25409 34629 25421 34663
rect 25455 34660 25467 34663
rect 25608 34660 25636 34688
rect 25455 34632 25636 34660
rect 25455 34629 25467 34632
rect 25409 34623 25467 34629
rect 26326 34620 26332 34672
rect 26384 34660 26390 34672
rect 26694 34660 26700 34672
rect 26384 34632 26700 34660
rect 26384 34620 26390 34632
rect 26694 34620 26700 34632
rect 26752 34660 26758 34672
rect 27816 34660 27844 34700
rect 28626 34660 28632 34672
rect 26752 34632 27844 34660
rect 28000 34632 28632 34660
rect 26752 34620 26758 34632
rect 25225 34595 25283 34601
rect 25225 34561 25237 34595
rect 25271 34561 25283 34595
rect 25225 34555 25283 34561
rect 25314 34552 25320 34604
rect 25372 34592 25378 34604
rect 25372 34564 25465 34592
rect 25372 34552 25378 34564
rect 25498 34552 25504 34604
rect 25556 34601 25562 34604
rect 25556 34595 25585 34601
rect 25573 34592 25585 34595
rect 25958 34592 25964 34604
rect 25573 34564 25964 34592
rect 25573 34561 25585 34564
rect 25556 34555 25585 34561
rect 25556 34552 25562 34555
rect 25958 34552 25964 34564
rect 26016 34552 26022 34604
rect 26237 34595 26295 34601
rect 26237 34561 26249 34595
rect 26283 34592 26295 34595
rect 26878 34592 26884 34604
rect 26283 34564 26884 34592
rect 26283 34561 26295 34564
rect 26237 34555 26295 34561
rect 22511 34496 23244 34524
rect 23293 34527 23351 34533
rect 22511 34493 22523 34496
rect 22465 34487 22523 34493
rect 23293 34493 23305 34527
rect 23339 34524 23351 34527
rect 23566 34524 23572 34536
rect 23339 34496 23572 34524
rect 23339 34493 23351 34496
rect 23293 34487 23351 34493
rect 23566 34484 23572 34496
rect 23624 34524 23630 34536
rect 24121 34527 24179 34533
rect 24121 34524 24133 34527
rect 23624 34496 24133 34524
rect 23624 34484 23630 34496
rect 24121 34493 24133 34496
rect 24167 34493 24179 34527
rect 24121 34487 24179 34493
rect 23474 34416 23480 34468
rect 23532 34456 23538 34468
rect 25332 34456 25360 34552
rect 25685 34527 25743 34533
rect 25685 34493 25697 34527
rect 25731 34524 25743 34527
rect 26050 34524 26056 34536
rect 25731 34496 26056 34524
rect 25731 34493 25743 34496
rect 25685 34487 25743 34493
rect 26050 34484 26056 34496
rect 26108 34484 26114 34536
rect 26252 34524 26280 34555
rect 26878 34552 26884 34564
rect 26936 34552 26942 34604
rect 27338 34552 27344 34604
rect 27396 34592 27402 34604
rect 28000 34601 28028 34632
rect 28626 34620 28632 34632
rect 28684 34620 28690 34672
rect 28828 34669 28856 34700
rect 29365 34697 29377 34731
rect 29411 34728 29423 34731
rect 30282 34728 30288 34740
rect 29411 34700 30288 34728
rect 29411 34697 29423 34700
rect 29365 34691 29423 34697
rect 30282 34688 30288 34700
rect 30340 34688 30346 34740
rect 28813 34663 28871 34669
rect 28813 34629 28825 34663
rect 28859 34660 28871 34663
rect 30558 34660 30564 34672
rect 28859 34632 29040 34660
rect 28859 34629 28871 34632
rect 28813 34623 28871 34629
rect 27893 34595 27951 34601
rect 27893 34592 27905 34595
rect 27396 34564 27905 34592
rect 27396 34552 27402 34564
rect 27893 34561 27905 34564
rect 27939 34561 27951 34595
rect 27893 34555 27951 34561
rect 27985 34595 28043 34601
rect 27985 34561 27997 34595
rect 28031 34561 28043 34595
rect 28261 34595 28319 34601
rect 28261 34592 28273 34595
rect 27985 34555 28043 34561
rect 28092 34564 28273 34592
rect 26326 34524 26332 34536
rect 26252 34496 26332 34524
rect 26326 34484 26332 34496
rect 26384 34484 26390 34536
rect 26421 34527 26479 34533
rect 26421 34493 26433 34527
rect 26467 34524 26479 34527
rect 26786 34524 26792 34536
rect 26467 34496 26792 34524
rect 26467 34493 26479 34496
rect 26421 34487 26479 34493
rect 26786 34484 26792 34496
rect 26844 34524 26850 34536
rect 28092 34524 28120 34564
rect 28261 34561 28273 34564
rect 28307 34561 28319 34595
rect 28718 34592 28724 34604
rect 28679 34564 28724 34592
rect 28261 34555 28319 34561
rect 28718 34552 28724 34564
rect 28776 34552 28782 34604
rect 28902 34592 28908 34604
rect 28863 34564 28908 34592
rect 28902 34552 28908 34564
rect 28960 34552 28966 34604
rect 26844 34496 28120 34524
rect 28169 34527 28227 34533
rect 26844 34484 26850 34496
rect 28169 34493 28181 34527
rect 28215 34524 28227 34527
rect 28810 34524 28816 34536
rect 28215 34496 28816 34524
rect 28215 34493 28227 34496
rect 28169 34487 28227 34493
rect 28810 34484 28816 34496
rect 28868 34484 28874 34536
rect 29012 34524 29040 34632
rect 29656 34632 30564 34660
rect 29454 34552 29460 34604
rect 29512 34592 29518 34604
rect 29656 34601 29684 34632
rect 30558 34620 30564 34632
rect 30616 34620 30622 34672
rect 29549 34595 29607 34601
rect 29549 34592 29561 34595
rect 29512 34564 29561 34592
rect 29512 34552 29518 34564
rect 29549 34561 29561 34564
rect 29595 34561 29607 34595
rect 29549 34555 29607 34561
rect 29641 34595 29699 34601
rect 29641 34561 29653 34595
rect 29687 34561 29699 34595
rect 29641 34555 29699 34561
rect 29825 34595 29883 34601
rect 29825 34561 29837 34595
rect 29871 34561 29883 34595
rect 29825 34555 29883 34561
rect 29840 34524 29868 34555
rect 29914 34552 29920 34604
rect 29972 34592 29978 34604
rect 47762 34592 47768 34604
rect 29972 34564 30017 34592
rect 47723 34564 47768 34592
rect 29972 34552 29978 34564
rect 47762 34552 47768 34564
rect 47820 34552 47826 34604
rect 29012 34496 29868 34524
rect 25958 34456 25964 34468
rect 23532 34428 24440 34456
rect 25332 34428 25964 34456
rect 23532 34416 23538 34428
rect 18680 34391 18738 34397
rect 18680 34357 18692 34391
rect 18726 34388 18738 34391
rect 19978 34388 19984 34400
rect 18726 34360 19984 34388
rect 18726 34357 18738 34360
rect 18680 34351 18738 34357
rect 19978 34348 19984 34360
rect 20036 34348 20042 34400
rect 20714 34388 20720 34400
rect 20675 34360 20720 34388
rect 20714 34348 20720 34360
rect 20772 34348 20778 34400
rect 21450 34348 21456 34400
rect 21508 34388 21514 34400
rect 22005 34391 22063 34397
rect 22005 34388 22017 34391
rect 21508 34360 22017 34388
rect 21508 34348 21514 34360
rect 22005 34357 22017 34360
rect 22051 34357 22063 34391
rect 24302 34388 24308 34400
rect 24263 34360 24308 34388
rect 22005 34351 22063 34357
rect 24302 34348 24308 34360
rect 24360 34348 24366 34400
rect 24412 34388 24440 34428
rect 25958 34416 25964 34428
rect 26016 34416 26022 34468
rect 30374 34388 30380 34400
rect 24412 34360 30380 34388
rect 30374 34348 30380 34360
rect 30432 34348 30438 34400
rect 47210 34348 47216 34400
rect 47268 34388 47274 34400
rect 47581 34391 47639 34397
rect 47581 34388 47593 34391
rect 47268 34360 47593 34388
rect 47268 34348 47274 34360
rect 47581 34357 47593 34360
rect 47627 34357 47639 34391
rect 47581 34351 47639 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 19978 34184 19984 34196
rect 6886 34156 19656 34184
rect 19939 34156 19984 34184
rect 1946 34008 1952 34060
rect 2004 34048 2010 34060
rect 6886 34048 6914 34156
rect 2004 34020 6914 34048
rect 15749 34051 15807 34057
rect 2004 34008 2010 34020
rect 15749 34017 15761 34051
rect 15795 34048 15807 34051
rect 16666 34048 16672 34060
rect 15795 34020 16672 34048
rect 15795 34017 15807 34020
rect 15749 34011 15807 34017
rect 16666 34008 16672 34020
rect 16724 34048 16730 34060
rect 18414 34048 18420 34060
rect 16724 34020 18420 34048
rect 16724 34008 16730 34020
rect 18414 34008 18420 34020
rect 18472 34048 18478 34060
rect 19334 34048 19340 34060
rect 18472 34020 19340 34048
rect 18472 34008 18478 34020
rect 19334 34008 19340 34020
rect 19392 34008 19398 34060
rect 19628 34057 19656 34156
rect 19978 34144 19984 34156
rect 20036 34144 20042 34196
rect 21450 34184 21456 34196
rect 21411 34156 21456 34184
rect 21450 34144 21456 34156
rect 21508 34144 21514 34196
rect 22281 34187 22339 34193
rect 22281 34153 22293 34187
rect 22327 34184 22339 34187
rect 23382 34184 23388 34196
rect 22327 34156 23388 34184
rect 22327 34153 22339 34156
rect 22281 34147 22339 34153
rect 23382 34144 23388 34156
rect 23440 34144 23446 34196
rect 23658 34184 23664 34196
rect 23619 34156 23664 34184
rect 23658 34144 23664 34156
rect 23716 34144 23722 34196
rect 24578 34144 24584 34196
rect 24636 34184 24642 34196
rect 25133 34187 25191 34193
rect 25133 34184 25145 34187
rect 24636 34156 25145 34184
rect 24636 34144 24642 34156
rect 25133 34153 25145 34156
rect 25179 34153 25191 34187
rect 25133 34147 25191 34153
rect 25317 34187 25375 34193
rect 25317 34153 25329 34187
rect 25363 34184 25375 34187
rect 25682 34184 25688 34196
rect 25363 34156 25688 34184
rect 25363 34153 25375 34156
rect 25317 34147 25375 34153
rect 25682 34144 25688 34156
rect 25740 34144 25746 34196
rect 28626 34144 28632 34196
rect 28684 34184 28690 34196
rect 28997 34187 29055 34193
rect 28997 34184 29009 34187
rect 28684 34156 29009 34184
rect 28684 34144 28690 34156
rect 28997 34153 29009 34156
rect 29043 34153 29055 34187
rect 28997 34147 29055 34153
rect 20990 34076 20996 34128
rect 21048 34116 21054 34128
rect 21637 34119 21695 34125
rect 21637 34116 21649 34119
rect 21048 34088 21649 34116
rect 21048 34076 21054 34088
rect 21637 34085 21649 34088
rect 21683 34085 21695 34119
rect 22370 34116 22376 34128
rect 21637 34079 21695 34085
rect 22112 34088 22376 34116
rect 19613 34051 19671 34057
rect 19613 34017 19625 34051
rect 19659 34017 19671 34051
rect 20898 34048 20904 34060
rect 19613 34011 19671 34017
rect 19720 34020 20904 34048
rect 1578 33980 1584 33992
rect 1539 33952 1584 33980
rect 1578 33940 1584 33952
rect 1636 33940 1642 33992
rect 19242 33980 19248 33992
rect 19203 33952 19248 33980
rect 19242 33940 19248 33952
rect 19300 33940 19306 33992
rect 19429 33983 19487 33989
rect 19429 33949 19441 33983
rect 19475 33949 19487 33983
rect 19429 33943 19487 33949
rect 19521 33983 19579 33989
rect 19521 33949 19533 33983
rect 19567 33980 19579 33983
rect 19720 33980 19748 34020
rect 20898 34008 20904 34020
rect 20956 34008 20962 34060
rect 19567 33952 19748 33980
rect 19797 33983 19855 33989
rect 19567 33949 19579 33952
rect 19521 33943 19579 33949
rect 19797 33949 19809 33983
rect 19843 33980 19855 33983
rect 20530 33980 20536 33992
rect 19843 33952 20536 33980
rect 19843 33949 19855 33952
rect 19797 33943 19855 33949
rect 16025 33915 16083 33921
rect 16025 33881 16037 33915
rect 16071 33881 16083 33915
rect 16025 33875 16083 33881
rect 1397 33847 1455 33853
rect 1397 33813 1409 33847
rect 1443 33844 1455 33847
rect 1946 33844 1952 33856
rect 1443 33816 1952 33844
rect 1443 33813 1455 33816
rect 1397 33807 1455 33813
rect 1946 33804 1952 33816
rect 2004 33804 2010 33856
rect 16040 33844 16068 33875
rect 16574 33872 16580 33924
rect 16632 33872 16638 33924
rect 19444 33912 19472 33943
rect 20530 33940 20536 33952
rect 20588 33940 20594 33992
rect 21082 33980 21088 33992
rect 21043 33952 21088 33980
rect 21082 33940 21088 33952
rect 21140 33940 21146 33992
rect 21358 33980 21364 33992
rect 21319 33952 21364 33980
rect 21358 33940 21364 33952
rect 21416 33940 21422 33992
rect 22112 33989 22140 34088
rect 22370 34076 22376 34088
rect 22428 34076 22434 34128
rect 22186 34008 22192 34060
rect 22244 34048 22250 34060
rect 22281 34051 22339 34057
rect 22281 34048 22293 34051
rect 22244 34020 22293 34048
rect 22244 34008 22250 34020
rect 22281 34017 22293 34020
rect 22327 34048 22339 34051
rect 22922 34048 22928 34060
rect 22327 34020 22928 34048
rect 22327 34017 22339 34020
rect 22281 34011 22339 34017
rect 22922 34008 22928 34020
rect 22980 34008 22986 34060
rect 27249 34051 27307 34057
rect 27249 34017 27261 34051
rect 27295 34048 27307 34051
rect 27522 34048 27528 34060
rect 27295 34020 27528 34048
rect 27295 34017 27307 34020
rect 27249 34011 27307 34017
rect 27522 34008 27528 34020
rect 27580 34008 27586 34060
rect 47118 34048 47124 34060
rect 47079 34020 47124 34048
rect 47118 34008 47124 34020
rect 47176 34008 47182 34060
rect 47670 34048 47676 34060
rect 47631 34020 47676 34048
rect 47670 34008 47676 34020
rect 47728 34008 47734 34060
rect 22097 33983 22155 33989
rect 22097 33949 22109 33983
rect 22143 33949 22155 33983
rect 22370 33980 22376 33992
rect 22331 33952 22376 33980
rect 22097 33943 22155 33949
rect 22370 33940 22376 33952
rect 22428 33940 22434 33992
rect 23566 33980 23572 33992
rect 23527 33952 23572 33980
rect 23566 33940 23572 33952
rect 23624 33940 23630 33992
rect 25498 33980 25504 33992
rect 24964 33952 25504 33980
rect 20070 33912 20076 33924
rect 19444 33884 20076 33912
rect 20070 33872 20076 33884
rect 20128 33872 20134 33924
rect 24964 33921 24992 33952
rect 25498 33940 25504 33952
rect 25556 33980 25562 33992
rect 25777 33983 25835 33989
rect 25777 33980 25789 33983
rect 25556 33952 25789 33980
rect 25556 33940 25562 33952
rect 25777 33949 25789 33952
rect 25823 33949 25835 33983
rect 30466 33980 30472 33992
rect 30427 33952 30472 33980
rect 25777 33943 25835 33949
rect 30466 33940 30472 33952
rect 30524 33940 30530 33992
rect 30834 33980 30840 33992
rect 30795 33952 30840 33980
rect 30834 33940 30840 33952
rect 30892 33940 30898 33992
rect 24949 33915 25007 33921
rect 24949 33881 24961 33915
rect 24995 33881 25007 33915
rect 24949 33875 25007 33881
rect 25165 33915 25223 33921
rect 25165 33881 25177 33915
rect 25211 33912 25223 33915
rect 25866 33912 25872 33924
rect 25211 33884 25872 33912
rect 25211 33881 25223 33884
rect 25165 33875 25223 33881
rect 25866 33872 25872 33884
rect 25924 33872 25930 33924
rect 27430 33872 27436 33924
rect 27488 33912 27494 33924
rect 27525 33915 27583 33921
rect 27525 33912 27537 33915
rect 27488 33884 27537 33912
rect 27488 33872 27494 33884
rect 27525 33881 27537 33884
rect 27571 33881 27583 33915
rect 29638 33912 29644 33924
rect 28750 33884 29644 33912
rect 27525 33875 27583 33881
rect 29638 33872 29644 33884
rect 29696 33872 29702 33924
rect 30374 33872 30380 33924
rect 30432 33912 30438 33924
rect 30653 33915 30711 33921
rect 30653 33912 30665 33915
rect 30432 33884 30665 33912
rect 30432 33872 30438 33884
rect 30653 33881 30665 33884
rect 30699 33881 30711 33915
rect 30653 33875 30711 33881
rect 30745 33915 30803 33921
rect 30745 33881 30757 33915
rect 30791 33881 30803 33915
rect 30745 33875 30803 33881
rect 16758 33844 16764 33856
rect 16040 33816 16764 33844
rect 16758 33804 16764 33816
rect 16816 33804 16822 33856
rect 17310 33804 17316 33856
rect 17368 33844 17374 33856
rect 17497 33847 17555 33853
rect 17497 33844 17509 33847
rect 17368 33816 17509 33844
rect 17368 33804 17374 33816
rect 17497 33813 17509 33816
rect 17543 33813 17555 33847
rect 17497 33807 17555 33813
rect 22278 33804 22284 33856
rect 22336 33844 22342 33856
rect 22557 33847 22615 33853
rect 22557 33844 22569 33847
rect 22336 33816 22569 33844
rect 22336 33804 22342 33816
rect 22557 33813 22569 33816
rect 22603 33813 22615 33847
rect 25958 33844 25964 33856
rect 25871 33816 25964 33844
rect 22557 33807 22615 33813
rect 25958 33804 25964 33816
rect 26016 33844 26022 33856
rect 27890 33844 27896 33856
rect 26016 33816 27896 33844
rect 26016 33804 26022 33816
rect 27890 33804 27896 33816
rect 27948 33804 27954 33856
rect 29730 33804 29736 33856
rect 29788 33844 29794 33856
rect 30760 33844 30788 33875
rect 47210 33872 47216 33924
rect 47268 33912 47274 33924
rect 47268 33884 47313 33912
rect 47268 33872 47274 33884
rect 29788 33816 30788 33844
rect 31021 33847 31079 33853
rect 29788 33804 29794 33816
rect 31021 33813 31033 33847
rect 31067 33844 31079 33847
rect 31294 33844 31300 33856
rect 31067 33816 31300 33844
rect 31067 33813 31079 33816
rect 31021 33807 31079 33813
rect 31294 33804 31300 33816
rect 31352 33804 31358 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 17034 33600 17040 33652
rect 17092 33640 17098 33652
rect 17497 33643 17555 33649
rect 17497 33640 17509 33643
rect 17092 33612 17509 33640
rect 17092 33600 17098 33612
rect 17497 33609 17509 33612
rect 17543 33609 17555 33643
rect 17497 33603 17555 33609
rect 19242 33600 19248 33652
rect 19300 33640 19306 33652
rect 20073 33643 20131 33649
rect 20073 33640 20085 33643
rect 19300 33612 20085 33640
rect 19300 33600 19306 33612
rect 20073 33609 20085 33612
rect 20119 33609 20131 33643
rect 28442 33640 28448 33652
rect 20073 33603 20131 33609
rect 24964 33612 28448 33640
rect 16945 33575 17003 33581
rect 16945 33541 16957 33575
rect 16991 33541 17003 33575
rect 16945 33535 17003 33541
rect 16666 33504 16672 33516
rect 16627 33476 16672 33504
rect 16666 33464 16672 33476
rect 16724 33464 16730 33516
rect 16960 33504 16988 33535
rect 17218 33532 17224 33584
rect 17276 33572 17282 33584
rect 17276 33544 19334 33572
rect 17276 33532 17282 33544
rect 17405 33507 17463 33513
rect 17405 33504 17417 33507
rect 16960 33476 17417 33504
rect 17405 33473 17417 33476
rect 17451 33473 17463 33507
rect 17405 33467 17463 33473
rect 17494 33464 17500 33516
rect 17552 33504 17558 33516
rect 17589 33507 17647 33513
rect 17589 33504 17601 33507
rect 17552 33476 17601 33504
rect 17552 33464 17558 33476
rect 17589 33473 17601 33476
rect 17635 33473 17647 33507
rect 19306 33504 19334 33544
rect 20898 33532 20904 33584
rect 20956 33572 20962 33584
rect 22005 33575 22063 33581
rect 22005 33572 22017 33575
rect 20956 33544 22017 33572
rect 20956 33532 20962 33544
rect 22005 33541 22017 33544
rect 22051 33541 22063 33575
rect 22005 33535 22063 33541
rect 24670 33532 24676 33584
rect 24728 33572 24734 33584
rect 24964 33572 24992 33612
rect 28442 33600 28448 33612
rect 28500 33600 28506 33652
rect 28813 33643 28871 33649
rect 28813 33609 28825 33643
rect 28859 33640 28871 33643
rect 29086 33640 29092 33652
rect 28859 33612 29092 33640
rect 28859 33609 28871 33612
rect 28813 33603 28871 33609
rect 29086 33600 29092 33612
rect 29144 33600 29150 33652
rect 47762 33600 47768 33652
rect 47820 33640 47826 33652
rect 48041 33643 48099 33649
rect 48041 33640 48053 33643
rect 47820 33612 48053 33640
rect 47820 33600 47826 33612
rect 48041 33609 48053 33612
rect 48087 33609 48099 33643
rect 48041 33603 48099 33609
rect 28902 33572 28908 33584
rect 24728 33544 24992 33572
rect 24728 33532 24734 33544
rect 19518 33504 19524 33516
rect 19306 33476 19524 33504
rect 17589 33467 17647 33473
rect 19518 33464 19524 33476
rect 19576 33464 19582 33516
rect 19889 33507 19947 33513
rect 19889 33473 19901 33507
rect 19935 33504 19947 33507
rect 20714 33504 20720 33516
rect 19935 33476 20720 33504
rect 19935 33473 19947 33476
rect 19889 33467 19947 33473
rect 20714 33464 20720 33476
rect 20772 33464 20778 33516
rect 21266 33464 21272 33516
rect 21324 33504 21330 33516
rect 21821 33507 21879 33513
rect 21821 33504 21833 33507
rect 21324 33476 21833 33504
rect 21324 33464 21330 33476
rect 21821 33473 21833 33476
rect 21867 33473 21879 33507
rect 22738 33504 22744 33516
rect 22699 33476 22744 33504
rect 21821 33467 21879 33473
rect 22738 33464 22744 33476
rect 22796 33464 22802 33516
rect 24489 33507 24547 33513
rect 24489 33473 24501 33507
rect 24535 33504 24547 33507
rect 24854 33504 24860 33516
rect 24535 33476 24860 33504
rect 24535 33473 24547 33476
rect 24489 33467 24547 33473
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 24964 33513 24992 33544
rect 28460 33544 28908 33572
rect 28460 33513 28488 33544
rect 28902 33532 28908 33544
rect 28960 33532 28966 33584
rect 24949 33507 25007 33513
rect 24949 33473 24961 33507
rect 24995 33473 25007 33507
rect 28445 33507 28503 33513
rect 28445 33504 28457 33507
rect 24949 33467 25007 33473
rect 27632 33476 28457 33504
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 1673 33439 1731 33445
rect 1673 33405 1685 33439
rect 1719 33436 1731 33439
rect 1854 33436 1860 33448
rect 1719 33408 1860 33436
rect 1719 33405 1731 33408
rect 1673 33399 1731 33405
rect 1854 33396 1860 33408
rect 1912 33396 1918 33448
rect 16945 33439 17003 33445
rect 16945 33405 16957 33439
rect 16991 33436 17003 33439
rect 17034 33436 17040 33448
rect 16991 33408 17040 33436
rect 16991 33405 17003 33408
rect 16945 33399 17003 33405
rect 17034 33396 17040 33408
rect 17092 33436 17098 33448
rect 17310 33436 17316 33448
rect 17092 33408 17316 33436
rect 17092 33396 17098 33408
rect 17310 33396 17316 33408
rect 17368 33396 17374 33448
rect 27632 33380 27660 33476
rect 28445 33473 28457 33476
rect 28491 33473 28503 33507
rect 28626 33504 28632 33516
rect 28587 33476 28632 33504
rect 28445 33467 28503 33473
rect 28626 33464 28632 33476
rect 28684 33464 28690 33516
rect 30466 33464 30472 33516
rect 30524 33504 30530 33516
rect 30929 33507 30987 33513
rect 30929 33504 30941 33507
rect 30524 33476 30941 33504
rect 30524 33464 30530 33476
rect 30929 33473 30941 33476
rect 30975 33504 30987 33507
rect 31018 33504 31024 33516
rect 30975 33476 31024 33504
rect 30975 33473 30987 33476
rect 30929 33467 30987 33473
rect 31018 33464 31024 33476
rect 31076 33464 31082 33516
rect 46842 33504 46848 33516
rect 46803 33476 46848 33504
rect 46842 33464 46848 33476
rect 46900 33464 46906 33516
rect 47581 33507 47639 33513
rect 47581 33473 47593 33507
rect 47627 33504 47639 33507
rect 47762 33504 47768 33516
rect 47627 33476 47768 33504
rect 47627 33473 47639 33476
rect 47581 33467 47639 33473
rect 47762 33464 47768 33476
rect 47820 33464 47826 33516
rect 30834 33436 30840 33448
rect 30795 33408 30840 33436
rect 30834 33396 30840 33408
rect 30892 33396 30898 33448
rect 19334 33328 19340 33380
rect 19392 33368 19398 33380
rect 22925 33371 22983 33377
rect 22925 33368 22937 33371
rect 19392 33340 22937 33368
rect 19392 33328 19398 33340
rect 22925 33337 22937 33340
rect 22971 33368 22983 33371
rect 23566 33368 23572 33380
rect 22971 33340 23572 33368
rect 22971 33337 22983 33340
rect 22925 33331 22983 33337
rect 23566 33328 23572 33340
rect 23624 33328 23630 33380
rect 23658 33328 23664 33380
rect 23716 33368 23722 33380
rect 27614 33368 27620 33380
rect 23716 33340 27620 33368
rect 23716 33328 23722 33340
rect 27614 33328 27620 33340
rect 27672 33328 27678 33380
rect 31297 33371 31355 33377
rect 31297 33337 31309 33371
rect 31343 33368 31355 33371
rect 31570 33368 31576 33380
rect 31343 33340 31576 33368
rect 31343 33337 31355 33340
rect 31297 33331 31355 33337
rect 31570 33328 31576 33340
rect 31628 33328 31634 33380
rect 16761 33303 16819 33309
rect 16761 33269 16773 33303
rect 16807 33300 16819 33303
rect 17218 33300 17224 33312
rect 16807 33272 17224 33300
rect 16807 33269 16819 33272
rect 16761 33263 16819 33269
rect 17218 33260 17224 33272
rect 17276 33260 17282 33312
rect 19889 33303 19947 33309
rect 19889 33269 19901 33303
rect 19935 33300 19947 33303
rect 20714 33300 20720 33312
rect 19935 33272 20720 33300
rect 19935 33269 19947 33272
rect 19889 33263 19947 33269
rect 20714 33260 20720 33272
rect 20772 33300 20778 33312
rect 21358 33300 21364 33312
rect 20772 33272 21364 33300
rect 20772 33260 20778 33272
rect 21358 33260 21364 33272
rect 21416 33260 21422 33312
rect 22189 33303 22247 33309
rect 22189 33269 22201 33303
rect 22235 33300 22247 33303
rect 22370 33300 22376 33312
rect 22235 33272 22376 33300
rect 22235 33269 22247 33272
rect 22189 33263 22247 33269
rect 22370 33260 22376 33272
rect 22428 33300 22434 33312
rect 23106 33300 23112 33312
rect 22428 33272 23112 33300
rect 22428 33260 22434 33272
rect 23106 33260 23112 33272
rect 23164 33260 23170 33312
rect 23842 33260 23848 33312
rect 23900 33300 23906 33312
rect 24305 33303 24363 33309
rect 24305 33300 24317 33303
rect 23900 33272 24317 33300
rect 23900 33260 23906 33272
rect 24305 33269 24317 33272
rect 24351 33269 24363 33303
rect 24305 33263 24363 33269
rect 24946 33260 24952 33312
rect 25004 33300 25010 33312
rect 25041 33303 25099 33309
rect 25041 33300 25053 33303
rect 25004 33272 25053 33300
rect 25004 33260 25010 33272
rect 25041 33269 25053 33272
rect 25087 33269 25099 33303
rect 25041 33263 25099 33269
rect 27338 33260 27344 33312
rect 27396 33300 27402 33312
rect 28445 33303 28503 33309
rect 28445 33300 28457 33303
rect 27396 33272 28457 33300
rect 27396 33260 27402 33272
rect 28445 33269 28457 33272
rect 28491 33300 28503 33303
rect 28534 33300 28540 33312
rect 28491 33272 28540 33300
rect 28491 33269 28503 33272
rect 28445 33263 28503 33269
rect 28534 33260 28540 33272
rect 28592 33300 28598 33312
rect 28718 33300 28724 33312
rect 28592 33272 28724 33300
rect 28592 33260 28598 33272
rect 28718 33260 28724 33272
rect 28776 33260 28782 33312
rect 41414 33260 41420 33312
rect 41472 33300 41478 33312
rect 46937 33303 46995 33309
rect 46937 33300 46949 33303
rect 41472 33272 46949 33300
rect 41472 33260 41478 33272
rect 46937 33269 46949 33272
rect 46983 33269 46995 33303
rect 47854 33300 47860 33312
rect 47815 33272 47860 33300
rect 46937 33263 46995 33269
rect 47854 33260 47860 33272
rect 47912 33260 47918 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1946 33096 1952 33108
rect 1907 33068 1952 33096
rect 1946 33056 1952 33068
rect 2004 33056 2010 33108
rect 16666 33056 16672 33108
rect 16724 33096 16730 33108
rect 17221 33099 17279 33105
rect 17221 33096 17233 33099
rect 16724 33068 17233 33096
rect 16724 33056 16730 33068
rect 17221 33065 17233 33068
rect 17267 33065 17279 33099
rect 17221 33059 17279 33065
rect 17494 33056 17500 33108
rect 17552 33096 17558 33108
rect 17589 33099 17647 33105
rect 17589 33096 17601 33099
rect 17552 33068 17601 33096
rect 17552 33056 17558 33068
rect 17589 33065 17601 33068
rect 17635 33065 17647 33099
rect 17589 33059 17647 33065
rect 17604 33028 17632 33059
rect 17770 33056 17776 33108
rect 17828 33096 17834 33108
rect 21177 33099 21235 33105
rect 21177 33096 21189 33099
rect 17828 33068 21189 33096
rect 17828 33056 17834 33068
rect 21177 33065 21189 33068
rect 21223 33065 21235 33099
rect 21177 33059 21235 33065
rect 21637 33099 21695 33105
rect 21637 33065 21649 33099
rect 21683 33096 21695 33099
rect 22186 33096 22192 33108
rect 21683 33068 22192 33096
rect 21683 33065 21695 33068
rect 21637 33059 21695 33065
rect 22186 33056 22192 33068
rect 22244 33056 22250 33108
rect 24854 33056 24860 33108
rect 24912 33096 24918 33108
rect 24949 33099 25007 33105
rect 24949 33096 24961 33099
rect 24912 33068 24961 33096
rect 24912 33056 24918 33068
rect 24949 33065 24961 33068
rect 24995 33065 25007 33099
rect 24949 33059 25007 33065
rect 25682 33056 25688 33108
rect 25740 33096 25746 33108
rect 26142 33096 26148 33108
rect 25740 33068 26148 33096
rect 25740 33056 25746 33068
rect 26142 33056 26148 33068
rect 26200 33096 26206 33108
rect 26237 33099 26295 33105
rect 26237 33096 26249 33099
rect 26200 33068 26249 33096
rect 26200 33056 26206 33068
rect 26237 33065 26249 33068
rect 26283 33065 26295 33099
rect 26237 33059 26295 33065
rect 27522 33056 27528 33108
rect 27580 33096 27586 33108
rect 28629 33099 28687 33105
rect 28629 33096 28641 33099
rect 27580 33068 28641 33096
rect 27580 33056 27586 33068
rect 28629 33065 28641 33068
rect 28675 33065 28687 33099
rect 29638 33096 29644 33108
rect 29599 33068 29644 33096
rect 28629 33059 28687 33065
rect 19613 33031 19671 33037
rect 19613 33028 19625 33031
rect 17604 33000 19625 33028
rect 19613 32997 19625 33000
rect 19659 32997 19671 33031
rect 19613 32991 19671 32997
rect 25516 33000 27752 33028
rect 2317 32963 2375 32969
rect 2317 32929 2329 32963
rect 2363 32929 2375 32963
rect 2317 32923 2375 32929
rect 1854 32892 1860 32904
rect 1815 32864 1860 32892
rect 1854 32852 1860 32864
rect 1912 32852 1918 32904
rect 2332 32892 2360 32923
rect 17034 32920 17040 32972
rect 17092 32960 17098 32972
rect 17313 32963 17371 32969
rect 17313 32960 17325 32963
rect 17092 32932 17325 32960
rect 17092 32920 17098 32932
rect 17313 32929 17325 32932
rect 17359 32960 17371 32963
rect 18414 32960 18420 32972
rect 17359 32932 18420 32960
rect 17359 32929 17371 32932
rect 17313 32923 17371 32929
rect 18414 32920 18420 32932
rect 18472 32960 18478 32972
rect 21361 32963 21419 32969
rect 18472 32932 20116 32960
rect 18472 32920 18478 32932
rect 2961 32895 3019 32901
rect 2961 32892 2973 32895
rect 2332 32864 2973 32892
rect 2961 32861 2973 32864
rect 3007 32861 3019 32895
rect 17218 32892 17224 32904
rect 17179 32864 17224 32892
rect 2961 32855 3019 32861
rect 17218 32852 17224 32864
rect 17276 32852 17282 32904
rect 18509 32895 18567 32901
rect 18509 32861 18521 32895
rect 18555 32892 18567 32895
rect 19242 32892 19248 32904
rect 18555 32864 19248 32892
rect 18555 32861 18567 32864
rect 18509 32855 18567 32861
rect 19242 32852 19248 32864
rect 19300 32892 19306 32904
rect 19429 32895 19487 32901
rect 19429 32892 19441 32895
rect 19300 32864 19441 32892
rect 19300 32852 19306 32864
rect 19429 32861 19441 32864
rect 19475 32861 19487 32895
rect 19429 32855 19487 32861
rect 19705 32895 19763 32901
rect 19705 32861 19717 32895
rect 19751 32892 19763 32895
rect 19978 32892 19984 32904
rect 19751 32864 19984 32892
rect 19751 32861 19763 32864
rect 19705 32855 19763 32861
rect 18325 32827 18383 32833
rect 18325 32793 18337 32827
rect 18371 32824 18383 32827
rect 18598 32824 18604 32836
rect 18371 32796 18604 32824
rect 18371 32793 18383 32796
rect 18325 32787 18383 32793
rect 18598 32784 18604 32796
rect 18656 32824 18662 32836
rect 19720 32824 19748 32855
rect 19978 32852 19984 32864
rect 20036 32852 20042 32904
rect 20088 32892 20116 32932
rect 21361 32929 21373 32963
rect 21407 32960 21419 32963
rect 22370 32960 22376 32972
rect 21407 32932 22376 32960
rect 21407 32929 21419 32932
rect 21361 32923 21419 32929
rect 22370 32920 22376 32932
rect 22428 32920 22434 32972
rect 21453 32895 21511 32901
rect 21453 32892 21465 32895
rect 20088 32864 21465 32892
rect 21453 32861 21465 32864
rect 21499 32861 21511 32895
rect 21453 32855 21511 32861
rect 22097 32895 22155 32901
rect 22097 32861 22109 32895
rect 22143 32892 22155 32895
rect 24486 32892 24492 32904
rect 22143 32864 24492 32892
rect 22143 32861 22155 32864
rect 22097 32855 22155 32861
rect 24486 32852 24492 32864
rect 24544 32852 24550 32904
rect 24673 32895 24731 32901
rect 24673 32861 24685 32895
rect 24719 32892 24731 32895
rect 25317 32895 25375 32901
rect 25317 32892 25329 32895
rect 24719 32864 25329 32892
rect 24719 32861 24731 32864
rect 24673 32855 24731 32861
rect 25317 32861 25329 32864
rect 25363 32892 25375 32895
rect 25516 32892 25544 33000
rect 25593 32963 25651 32969
rect 25593 32929 25605 32963
rect 25639 32960 25651 32963
rect 26326 32960 26332 32972
rect 25639 32932 26332 32960
rect 25639 32929 25651 32932
rect 25593 32923 25651 32929
rect 26326 32920 26332 32932
rect 26384 32920 26390 32972
rect 27433 32963 27491 32969
rect 27433 32929 27445 32963
rect 27479 32960 27491 32963
rect 27614 32960 27620 32972
rect 27479 32932 27620 32960
rect 27479 32929 27491 32932
rect 27433 32923 27491 32929
rect 27614 32920 27620 32932
rect 27672 32920 27678 32972
rect 25363 32864 25544 32892
rect 26145 32895 26203 32901
rect 25363 32861 25375 32864
rect 25317 32855 25375 32861
rect 26145 32861 26157 32895
rect 26191 32861 26203 32895
rect 26145 32855 26203 32861
rect 18656 32796 19748 32824
rect 21177 32827 21235 32833
rect 18656 32784 18662 32796
rect 21177 32793 21189 32827
rect 21223 32824 21235 32827
rect 21266 32824 21272 32836
rect 21223 32796 21272 32824
rect 21223 32793 21235 32796
rect 21177 32787 21235 32793
rect 21266 32784 21272 32796
rect 21324 32784 21330 32836
rect 26160 32824 26188 32855
rect 27338 32852 27344 32904
rect 27396 32892 27402 32904
rect 27525 32895 27583 32901
rect 27525 32892 27537 32895
rect 27396 32864 27537 32892
rect 27396 32852 27402 32864
rect 27525 32861 27537 32864
rect 27571 32861 27583 32895
rect 27724 32892 27752 33000
rect 27893 32963 27951 32969
rect 27893 32929 27905 32963
rect 27939 32960 27951 32963
rect 28534 32960 28540 32972
rect 27939 32932 28540 32960
rect 27939 32929 27951 32932
rect 27893 32923 27951 32929
rect 28534 32920 28540 32932
rect 28592 32920 28598 32972
rect 28644 32960 28672 33059
rect 29638 33056 29644 33068
rect 29696 33056 29702 33108
rect 28810 32988 28816 33040
rect 28868 33028 28874 33040
rect 28868 33000 31248 33028
rect 28868 32988 28874 33000
rect 31110 32960 31116 32972
rect 28644 32932 31116 32960
rect 31110 32920 31116 32932
rect 31168 32920 31174 32972
rect 31220 32960 31248 33000
rect 47026 32960 47032 32972
rect 31220 32932 47032 32960
rect 47026 32920 47032 32932
rect 47084 32920 47090 32972
rect 29546 32892 29552 32904
rect 27724 32864 28672 32892
rect 29507 32864 29552 32892
rect 27525 32855 27583 32861
rect 26234 32824 26240 32836
rect 26160 32796 26240 32824
rect 26234 32784 26240 32796
rect 26292 32784 26298 32836
rect 28258 32784 28264 32836
rect 28316 32824 28322 32836
rect 28537 32827 28595 32833
rect 28537 32824 28549 32827
rect 28316 32796 28549 32824
rect 28316 32784 28322 32796
rect 28537 32793 28549 32796
rect 28583 32793 28595 32827
rect 28644 32824 28672 32864
rect 29546 32852 29552 32864
rect 29604 32852 29610 32904
rect 46290 32892 46296 32904
rect 46251 32864 46296 32892
rect 46290 32852 46296 32864
rect 46348 32852 46354 32904
rect 30558 32824 30564 32836
rect 28644 32796 30564 32824
rect 28537 32787 28595 32793
rect 30558 32784 30564 32796
rect 30616 32784 30622 32836
rect 31386 32824 31392 32836
rect 31347 32796 31392 32824
rect 31386 32784 31392 32796
rect 31444 32784 31450 32836
rect 33686 32824 33692 32836
rect 32614 32796 33692 32824
rect 33686 32784 33692 32796
rect 33744 32784 33750 32836
rect 46477 32827 46535 32833
rect 46477 32793 46489 32827
rect 46523 32824 46535 32827
rect 46934 32824 46940 32836
rect 46523 32796 46940 32824
rect 46523 32793 46535 32796
rect 46477 32787 46535 32793
rect 46934 32784 46940 32796
rect 46992 32784 46998 32836
rect 48130 32824 48136 32836
rect 48091 32796 48136 32824
rect 48130 32784 48136 32796
rect 48188 32784 48194 32836
rect 2314 32716 2320 32768
rect 2372 32756 2378 32768
rect 2777 32759 2835 32765
rect 2777 32756 2789 32759
rect 2372 32728 2789 32756
rect 2372 32716 2378 32728
rect 2777 32725 2789 32728
rect 2823 32725 2835 32759
rect 2777 32719 2835 32725
rect 18230 32716 18236 32768
rect 18288 32756 18294 32768
rect 18693 32759 18751 32765
rect 18693 32756 18705 32759
rect 18288 32728 18705 32756
rect 18288 32716 18294 32728
rect 18693 32725 18705 32728
rect 18739 32725 18751 32759
rect 18693 32719 18751 32725
rect 19245 32759 19303 32765
rect 19245 32725 19257 32759
rect 19291 32756 19303 32759
rect 19334 32756 19340 32768
rect 19291 32728 19340 32756
rect 19291 32725 19303 32728
rect 19245 32719 19303 32725
rect 19334 32716 19340 32728
rect 19392 32716 19398 32768
rect 20806 32716 20812 32768
rect 20864 32756 20870 32768
rect 22189 32759 22247 32765
rect 22189 32756 22201 32759
rect 20864 32728 22201 32756
rect 20864 32716 20870 32728
rect 22189 32725 22201 32728
rect 22235 32725 22247 32759
rect 22189 32719 22247 32725
rect 25406 32716 25412 32768
rect 25464 32756 25470 32768
rect 25464 32728 25509 32756
rect 25464 32716 25470 32728
rect 28442 32716 28448 32768
rect 28500 32756 28506 32768
rect 29546 32756 29552 32768
rect 28500 32728 29552 32756
rect 28500 32716 28506 32728
rect 29546 32716 29552 32728
rect 29604 32716 29610 32768
rect 30650 32716 30656 32768
rect 30708 32756 30714 32768
rect 31018 32756 31024 32768
rect 30708 32728 31024 32756
rect 30708 32716 30714 32728
rect 31018 32716 31024 32728
rect 31076 32756 31082 32768
rect 31662 32756 31668 32768
rect 31076 32728 31668 32756
rect 31076 32716 31082 32728
rect 31662 32716 31668 32728
rect 31720 32756 31726 32768
rect 32861 32759 32919 32765
rect 32861 32756 32873 32759
rect 31720 32728 32873 32756
rect 31720 32716 31726 32728
rect 32861 32725 32873 32728
rect 32907 32725 32919 32759
rect 32861 32719 32919 32725
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 21266 32552 21272 32564
rect 21227 32524 21272 32552
rect 21266 32512 21272 32524
rect 21324 32512 21330 32564
rect 22738 32512 22744 32564
rect 22796 32552 22802 32564
rect 23017 32555 23075 32561
rect 23017 32552 23029 32555
rect 22796 32524 23029 32552
rect 22796 32512 22802 32524
rect 23017 32521 23029 32524
rect 23063 32521 23075 32555
rect 23017 32515 23075 32521
rect 23106 32512 23112 32564
rect 23164 32552 23170 32564
rect 27525 32555 27583 32561
rect 27525 32552 27537 32555
rect 23164 32524 25176 32552
rect 23164 32512 23170 32524
rect 2314 32484 2320 32496
rect 2275 32456 2320 32484
rect 2314 32444 2320 32456
rect 2372 32444 2378 32496
rect 23842 32484 23848 32496
rect 19076 32456 22232 32484
rect 23803 32456 23848 32484
rect 2130 32416 2136 32428
rect 2091 32388 2136 32416
rect 2130 32376 2136 32388
rect 2188 32376 2194 32428
rect 16666 32376 16672 32428
rect 16724 32416 16730 32428
rect 16853 32419 16911 32425
rect 16853 32416 16865 32419
rect 16724 32388 16865 32416
rect 16724 32376 16730 32388
rect 16853 32385 16865 32388
rect 16899 32416 16911 32419
rect 17770 32416 17776 32428
rect 16899 32388 17356 32416
rect 17731 32388 17776 32416
rect 16899 32385 16911 32388
rect 16853 32379 16911 32385
rect 3973 32351 4031 32357
rect 3973 32317 3985 32351
rect 4019 32348 4031 32351
rect 4614 32348 4620 32360
rect 4019 32320 4620 32348
rect 4019 32317 4031 32320
rect 3973 32311 4031 32317
rect 4614 32308 4620 32320
rect 4672 32308 4678 32360
rect 16945 32351 17003 32357
rect 16945 32317 16957 32351
rect 16991 32348 17003 32351
rect 17218 32348 17224 32360
rect 16991 32320 17224 32348
rect 16991 32317 17003 32320
rect 16945 32311 17003 32317
rect 17218 32308 17224 32320
rect 17276 32308 17282 32360
rect 17328 32348 17356 32388
rect 17770 32376 17776 32388
rect 17828 32376 17834 32428
rect 18966 32376 18972 32428
rect 19024 32416 19030 32428
rect 19076 32425 19104 32456
rect 19061 32419 19119 32425
rect 19061 32416 19073 32419
rect 19024 32388 19073 32416
rect 19024 32376 19030 32388
rect 19061 32385 19073 32388
rect 19107 32385 19119 32419
rect 19334 32416 19340 32428
rect 19295 32388 19340 32416
rect 19061 32379 19119 32385
rect 19334 32376 19340 32388
rect 19392 32376 19398 32428
rect 19978 32376 19984 32428
rect 20036 32416 20042 32428
rect 22204 32425 22232 32456
rect 23842 32444 23848 32456
rect 23900 32444 23906 32496
rect 20809 32419 20867 32425
rect 20809 32416 20821 32419
rect 20036 32388 20821 32416
rect 20036 32376 20042 32388
rect 20809 32385 20821 32388
rect 20855 32385 20867 32419
rect 20809 32379 20867 32385
rect 21085 32419 21143 32425
rect 21085 32385 21097 32419
rect 21131 32416 21143 32419
rect 22189 32419 22247 32425
rect 21131 32388 22140 32416
rect 21131 32385 21143 32388
rect 21085 32379 21143 32385
rect 18046 32348 18052 32360
rect 17328 32320 18052 32348
rect 18046 32308 18052 32320
rect 18104 32308 18110 32360
rect 19242 32308 19248 32360
rect 19300 32348 19306 32360
rect 20901 32351 20959 32357
rect 20901 32348 20913 32351
rect 19300 32320 20913 32348
rect 19300 32308 19306 32320
rect 20901 32317 20913 32320
rect 20947 32348 20959 32351
rect 21174 32348 21180 32360
rect 20947 32320 21180 32348
rect 20947 32317 20959 32320
rect 20901 32311 20959 32317
rect 21174 32308 21180 32320
rect 21232 32308 21238 32360
rect 22005 32351 22063 32357
rect 22005 32317 22017 32351
rect 22051 32317 22063 32351
rect 22112 32348 22140 32388
rect 22189 32385 22201 32419
rect 22235 32416 22247 32419
rect 22554 32416 22560 32428
rect 22235 32388 22560 32416
rect 22235 32385 22247 32388
rect 22189 32379 22247 32385
rect 22554 32376 22560 32388
rect 22612 32376 22618 32428
rect 22922 32416 22928 32428
rect 22883 32388 22928 32416
rect 22922 32376 22928 32388
rect 22980 32376 22986 32428
rect 23566 32416 23572 32428
rect 23527 32388 23572 32416
rect 23566 32376 23572 32388
rect 23624 32376 23630 32428
rect 24946 32376 24952 32428
rect 25004 32376 25010 32428
rect 25148 32416 25176 32524
rect 25792 32524 27537 32552
rect 25590 32444 25596 32496
rect 25648 32484 25654 32496
rect 25792 32493 25820 32524
rect 27525 32521 27537 32524
rect 27571 32521 27583 32555
rect 27525 32515 27583 32521
rect 28626 32512 28632 32564
rect 28684 32552 28690 32564
rect 30561 32555 30619 32561
rect 30561 32552 30573 32555
rect 28684 32524 30573 32552
rect 28684 32512 28690 32524
rect 30561 32521 30573 32524
rect 30607 32521 30619 32555
rect 30561 32515 30619 32521
rect 31113 32555 31171 32561
rect 31113 32521 31125 32555
rect 31159 32552 31171 32555
rect 31386 32552 31392 32564
rect 31159 32524 31392 32552
rect 31159 32521 31171 32524
rect 31113 32515 31171 32521
rect 31386 32512 31392 32524
rect 31444 32512 31450 32564
rect 33686 32552 33692 32564
rect 33647 32524 33692 32552
rect 33686 32512 33692 32524
rect 33744 32512 33750 32564
rect 46934 32552 46940 32564
rect 46895 32524 46940 32552
rect 46934 32512 46940 32524
rect 46992 32512 46998 32564
rect 47026 32512 47032 32564
rect 47084 32552 47090 32564
rect 48041 32555 48099 32561
rect 48041 32552 48053 32555
rect 47084 32524 48053 32552
rect 47084 32512 47090 32524
rect 48041 32521 48053 32524
rect 48087 32521 48099 32555
rect 48041 32515 48099 32521
rect 25777 32487 25835 32493
rect 25777 32484 25789 32487
rect 25648 32456 25789 32484
rect 25648 32444 25654 32456
rect 25777 32453 25789 32456
rect 25823 32453 25835 32487
rect 25777 32447 25835 32453
rect 25866 32444 25872 32496
rect 25924 32484 25930 32496
rect 25977 32487 26035 32493
rect 25977 32484 25989 32487
rect 25924 32456 25989 32484
rect 25924 32444 25930 32456
rect 25977 32453 25989 32456
rect 26023 32453 26035 32487
rect 25977 32447 26035 32453
rect 26234 32444 26240 32496
rect 26292 32484 26298 32496
rect 27433 32487 27491 32493
rect 27433 32484 27445 32487
rect 26292 32456 27445 32484
rect 26292 32444 26298 32456
rect 27433 32453 27445 32456
rect 27479 32484 27491 32487
rect 41414 32484 41420 32496
rect 27479 32456 41420 32484
rect 27479 32453 27491 32456
rect 27433 32447 27491 32453
rect 41414 32444 41420 32456
rect 41472 32444 41478 32496
rect 25148 32388 28120 32416
rect 24578 32348 24584 32360
rect 22112 32320 24584 32348
rect 22005 32311 22063 32317
rect 17236 32280 17264 32308
rect 17678 32280 17684 32292
rect 17236 32252 17684 32280
rect 17678 32240 17684 32252
rect 17736 32240 17742 32292
rect 20714 32280 20720 32292
rect 19260 32252 20720 32280
rect 1394 32172 1400 32224
rect 1452 32212 1458 32224
rect 1673 32215 1731 32221
rect 1673 32212 1685 32215
rect 1452 32184 1685 32212
rect 1452 32172 1458 32184
rect 1673 32181 1685 32184
rect 1719 32181 1731 32215
rect 17218 32212 17224 32224
rect 17179 32184 17224 32212
rect 1673 32175 1731 32181
rect 17218 32172 17224 32184
rect 17276 32172 17282 32224
rect 17310 32172 17316 32224
rect 17368 32212 17374 32224
rect 18690 32212 18696 32224
rect 17368 32184 18696 32212
rect 17368 32172 17374 32184
rect 18690 32172 18696 32184
rect 18748 32172 18754 32224
rect 19260 32221 19288 32252
rect 20714 32240 20720 32252
rect 20772 32240 20778 32292
rect 19245 32215 19303 32221
rect 19245 32181 19257 32215
rect 19291 32181 19303 32215
rect 19245 32175 19303 32181
rect 19334 32172 19340 32224
rect 19392 32212 19398 32224
rect 19613 32215 19671 32221
rect 19613 32212 19625 32215
rect 19392 32184 19625 32212
rect 19392 32172 19398 32184
rect 19613 32181 19625 32184
rect 19659 32181 19671 32215
rect 19613 32175 19671 32181
rect 21085 32215 21143 32221
rect 21085 32181 21097 32215
rect 21131 32212 21143 32215
rect 21358 32212 21364 32224
rect 21131 32184 21364 32212
rect 21131 32181 21143 32184
rect 21085 32175 21143 32181
rect 21358 32172 21364 32184
rect 21416 32212 21422 32224
rect 22020 32212 22048 32311
rect 24578 32308 24584 32320
rect 24636 32348 24642 32360
rect 25317 32351 25375 32357
rect 25317 32348 25329 32351
rect 24636 32320 25329 32348
rect 24636 32308 24642 32320
rect 25317 32317 25329 32320
rect 25363 32317 25375 32351
rect 25317 32311 25375 32317
rect 25958 32308 25964 32360
rect 26016 32348 26022 32360
rect 28092 32348 28120 32388
rect 28166 32376 28172 32428
rect 28224 32416 28230 32428
rect 28353 32419 28411 32425
rect 28224 32388 28269 32416
rect 28224 32376 28230 32388
rect 28353 32385 28365 32419
rect 28399 32416 28411 32419
rect 28442 32416 28448 32428
rect 28399 32388 28448 32416
rect 28399 32385 28411 32388
rect 28353 32379 28411 32385
rect 28442 32376 28448 32388
rect 28500 32376 28506 32428
rect 28534 32376 28540 32428
rect 28592 32416 28598 32428
rect 28813 32419 28871 32425
rect 28813 32416 28825 32419
rect 28592 32388 28825 32416
rect 28592 32376 28598 32388
rect 28813 32385 28825 32388
rect 28859 32385 28871 32419
rect 28994 32416 29000 32428
rect 28955 32388 29000 32416
rect 28813 32379 28871 32385
rect 28994 32376 29000 32388
rect 29052 32376 29058 32428
rect 29917 32419 29975 32425
rect 29917 32385 29929 32419
rect 29963 32385 29975 32419
rect 29917 32379 29975 32385
rect 30064 32419 30122 32425
rect 30064 32385 30076 32419
rect 30110 32416 30122 32419
rect 31294 32416 31300 32428
rect 30110 32388 30972 32416
rect 31255 32388 31300 32416
rect 30110 32385 30122 32388
rect 30064 32379 30122 32385
rect 29932 32348 29960 32379
rect 26016 32320 26832 32348
rect 28092 32320 29960 32348
rect 30285 32351 30343 32357
rect 26016 32308 26022 32320
rect 24854 32240 24860 32292
rect 24912 32280 24918 32292
rect 26145 32283 26203 32289
rect 26145 32280 26157 32283
rect 24912 32252 26157 32280
rect 24912 32240 24918 32252
rect 26145 32249 26157 32252
rect 26191 32249 26203 32283
rect 26145 32243 26203 32249
rect 22370 32212 22376 32224
rect 21416 32184 22048 32212
rect 22331 32184 22376 32212
rect 21416 32172 21422 32184
rect 22370 32172 22376 32184
rect 22428 32172 22434 32224
rect 22462 32172 22468 32224
rect 22520 32212 22526 32224
rect 23934 32212 23940 32224
rect 22520 32184 23940 32212
rect 22520 32172 22526 32184
rect 23934 32172 23940 32184
rect 23992 32172 23998 32224
rect 25130 32172 25136 32224
rect 25188 32212 25194 32224
rect 25314 32212 25320 32224
rect 25188 32184 25320 32212
rect 25188 32172 25194 32184
rect 25314 32172 25320 32184
rect 25372 32212 25378 32224
rect 25961 32215 26019 32221
rect 25961 32212 25973 32215
rect 25372 32184 25973 32212
rect 25372 32172 25378 32184
rect 25961 32181 25973 32184
rect 26007 32181 26019 32215
rect 26804 32212 26832 32320
rect 30285 32317 30297 32351
rect 30331 32348 30343 32351
rect 30834 32348 30840 32360
rect 30331 32320 30840 32348
rect 30331 32317 30343 32320
rect 30285 32311 30343 32317
rect 30834 32308 30840 32320
rect 30892 32308 30898 32360
rect 30944 32348 30972 32388
rect 31294 32376 31300 32388
rect 31352 32376 31358 32428
rect 31478 32416 31484 32428
rect 31439 32388 31484 32416
rect 31478 32376 31484 32388
rect 31536 32376 31542 32428
rect 31570 32376 31576 32428
rect 31628 32416 31634 32428
rect 31628 32388 31673 32416
rect 31628 32376 31634 32388
rect 31754 32376 31760 32428
rect 31812 32416 31818 32428
rect 32125 32419 32183 32425
rect 32125 32416 32137 32419
rect 31812 32388 32137 32416
rect 31812 32376 31818 32388
rect 32125 32385 32137 32388
rect 32171 32385 32183 32419
rect 32125 32379 32183 32385
rect 32309 32419 32367 32425
rect 32309 32385 32321 32419
rect 32355 32416 32367 32419
rect 32953 32419 33011 32425
rect 32355 32388 32720 32416
rect 32355 32385 32367 32388
rect 32309 32379 32367 32385
rect 32692 32360 32720 32388
rect 32953 32385 32965 32419
rect 32999 32385 33011 32419
rect 32953 32379 33011 32385
rect 33597 32419 33655 32425
rect 33597 32385 33609 32419
rect 33643 32416 33655 32419
rect 33686 32416 33692 32428
rect 33643 32388 33692 32416
rect 33643 32385 33655 32388
rect 33597 32379 33655 32385
rect 31018 32348 31024 32360
rect 30944 32320 31024 32348
rect 31018 32308 31024 32320
rect 31076 32348 31082 32360
rect 32493 32351 32551 32357
rect 32493 32348 32505 32351
rect 31076 32320 32505 32348
rect 31076 32308 31082 32320
rect 32493 32317 32505 32320
rect 32539 32317 32551 32351
rect 32493 32311 32551 32317
rect 32674 32308 32680 32360
rect 32732 32348 32738 32360
rect 32968 32348 32996 32379
rect 33686 32376 33692 32388
rect 33744 32376 33750 32428
rect 46198 32376 46204 32428
rect 46256 32416 46262 32428
rect 46845 32419 46903 32425
rect 46845 32416 46857 32419
rect 46256 32388 46857 32416
rect 46256 32376 46262 32388
rect 46845 32385 46857 32388
rect 46891 32385 46903 32419
rect 47946 32416 47952 32428
rect 47907 32388 47952 32416
rect 46845 32379 46903 32385
rect 47946 32376 47952 32388
rect 48004 32376 48010 32428
rect 34146 32348 34152 32360
rect 32732 32320 34152 32348
rect 32732 32308 32738 32320
rect 34146 32308 34152 32320
rect 34204 32308 34210 32360
rect 47394 32348 47400 32360
rect 35866 32320 47400 32348
rect 26878 32240 26884 32292
rect 26936 32280 26942 32292
rect 30466 32280 30472 32292
rect 26936 32252 30472 32280
rect 26936 32240 26942 32252
rect 30466 32240 30472 32252
rect 30524 32240 30530 32292
rect 31294 32240 31300 32292
rect 31352 32280 31358 32292
rect 33045 32283 33103 32289
rect 33045 32280 33057 32283
rect 31352 32252 33057 32280
rect 31352 32240 31358 32252
rect 33045 32249 33057 32252
rect 33091 32249 33103 32283
rect 33045 32243 33103 32249
rect 28074 32212 28080 32224
rect 26804 32184 28080 32212
rect 25961 32175 26019 32181
rect 28074 32172 28080 32184
rect 28132 32172 28138 32224
rect 28258 32172 28264 32224
rect 28316 32212 28322 32224
rect 28813 32215 28871 32221
rect 28813 32212 28825 32215
rect 28316 32184 28825 32212
rect 28316 32172 28322 32184
rect 28813 32181 28825 32184
rect 28859 32181 28871 32215
rect 28813 32175 28871 32181
rect 30190 32172 30196 32224
rect 30248 32212 30254 32224
rect 30248 32184 30293 32212
rect 30248 32172 30254 32184
rect 30558 32172 30564 32224
rect 30616 32212 30622 32224
rect 35866 32212 35894 32320
rect 47394 32308 47400 32320
rect 47452 32308 47458 32360
rect 30616 32184 35894 32212
rect 30616 32172 30622 32184
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 17310 32008 17316 32020
rect 7484 31980 17316 32008
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 1581 31875 1639 31881
rect 1581 31841 1593 31875
rect 1627 31872 1639 31875
rect 3881 31875 3939 31881
rect 3881 31872 3893 31875
rect 1627 31844 3893 31872
rect 1627 31841 1639 31844
rect 1581 31835 1639 31841
rect 3881 31841 3893 31844
rect 3927 31841 3939 31875
rect 3881 31835 3939 31841
rect 3234 31804 3240 31816
rect 3195 31776 3240 31804
rect 3234 31764 3240 31776
rect 3292 31764 3298 31816
rect 3786 31804 3792 31816
rect 3699 31776 3792 31804
rect 3786 31764 3792 31776
rect 3844 31804 3850 31816
rect 3970 31804 3976 31816
rect 3844 31776 3976 31804
rect 3844 31764 3850 31776
rect 3970 31764 3976 31776
rect 4028 31764 4034 31816
rect 7484 31813 7512 31980
rect 17310 31968 17316 31980
rect 17368 31968 17374 32020
rect 18233 32011 18291 32017
rect 18233 31977 18245 32011
rect 18279 31977 18291 32011
rect 18233 31971 18291 31977
rect 17589 31943 17647 31949
rect 17589 31909 17601 31943
rect 17635 31940 17647 31943
rect 17770 31940 17776 31952
rect 17635 31912 17776 31940
rect 17635 31909 17647 31912
rect 17589 31903 17647 31909
rect 17770 31900 17776 31912
rect 17828 31900 17834 31952
rect 18046 31900 18052 31952
rect 18104 31940 18110 31952
rect 18248 31940 18276 31971
rect 18690 31968 18696 32020
rect 18748 32008 18754 32020
rect 18748 31980 22324 32008
rect 18748 31968 18754 31980
rect 21174 31940 21180 31952
rect 18104 31912 18276 31940
rect 21135 31912 21180 31940
rect 18104 31900 18110 31912
rect 21174 31900 21180 31912
rect 21232 31900 21238 31952
rect 22296 31940 22324 31980
rect 22922 31968 22928 32020
rect 22980 32008 22986 32020
rect 26237 32011 26295 32017
rect 26237 32008 26249 32011
rect 22980 31980 26249 32008
rect 22980 31968 22986 31980
rect 26237 31977 26249 31980
rect 26283 32008 26295 32011
rect 28166 32008 28172 32020
rect 26283 31980 28172 32008
rect 26283 31977 26295 31980
rect 26237 31971 26295 31977
rect 28166 31968 28172 31980
rect 28224 31968 28230 32020
rect 28902 31968 28908 32020
rect 28960 32008 28966 32020
rect 29362 32008 29368 32020
rect 28960 31980 29368 32008
rect 28960 31968 28966 31980
rect 29362 31968 29368 31980
rect 29420 31968 29426 32020
rect 30190 31968 30196 32020
rect 30248 32008 30254 32020
rect 30377 32011 30435 32017
rect 30377 32008 30389 32011
rect 30248 31980 30389 32008
rect 30248 31968 30254 31980
rect 30377 31977 30389 31980
rect 30423 31977 30435 32011
rect 30377 31971 30435 31977
rect 30466 31968 30472 32020
rect 30524 32008 30530 32020
rect 39850 32008 39856 32020
rect 30524 31980 39856 32008
rect 30524 31968 30530 31980
rect 39850 31968 39856 31980
rect 39908 31968 39914 32020
rect 46290 31968 46296 32020
rect 46348 32008 46354 32020
rect 47673 32011 47731 32017
rect 47673 32008 47685 32011
rect 46348 31980 47685 32008
rect 46348 31968 46354 31980
rect 47673 31977 47685 31980
rect 47719 31977 47731 32011
rect 47673 31971 47731 31977
rect 26878 31940 26884 31952
rect 22296 31912 26884 31940
rect 26878 31900 26884 31912
rect 26936 31900 26942 31952
rect 30006 31940 30012 31952
rect 28460 31912 30012 31940
rect 15841 31875 15899 31881
rect 15841 31841 15853 31875
rect 15887 31872 15899 31875
rect 16850 31872 16856 31884
rect 15887 31844 16856 31872
rect 15887 31841 15899 31844
rect 15841 31835 15899 31841
rect 16850 31832 16856 31844
rect 16908 31872 16914 31884
rect 16908 31844 17356 31872
rect 16908 31832 16914 31844
rect 7469 31807 7527 31813
rect 7469 31773 7481 31807
rect 7515 31773 7527 31807
rect 17328 31804 17356 31844
rect 17678 31832 17684 31884
rect 17736 31872 17742 31884
rect 17736 31844 18276 31872
rect 17736 31832 17742 31844
rect 17328 31776 18000 31804
rect 7469 31767 7527 31773
rect 16117 31739 16175 31745
rect 16117 31705 16129 31739
rect 16163 31705 16175 31739
rect 17862 31736 17868 31748
rect 17342 31708 17868 31736
rect 16117 31699 16175 31705
rect 7558 31668 7564 31680
rect 7519 31640 7564 31668
rect 7558 31628 7564 31640
rect 7616 31628 7622 31680
rect 16132 31668 16160 31699
rect 17862 31696 17868 31708
rect 17920 31696 17926 31748
rect 17126 31668 17132 31680
rect 16132 31640 17132 31668
rect 17126 31628 17132 31640
rect 17184 31628 17190 31680
rect 17972 31668 18000 31776
rect 18248 31745 18276 31844
rect 18322 31832 18328 31884
rect 18380 31872 18386 31884
rect 18380 31844 18425 31872
rect 18380 31832 18386 31844
rect 18690 31832 18696 31884
rect 18748 31872 18754 31884
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 18748 31844 19441 31872
rect 18748 31832 18754 31844
rect 19429 31841 19441 31844
rect 19475 31872 19487 31875
rect 22462 31872 22468 31884
rect 19475 31844 22140 31872
rect 22423 31844 22468 31872
rect 19475 31841 19487 31844
rect 19429 31835 19487 31841
rect 22112 31816 22140 31844
rect 22462 31832 22468 31844
rect 22520 31832 22526 31884
rect 22554 31832 22560 31884
rect 22612 31872 22618 31884
rect 23753 31875 23811 31881
rect 22612 31844 23704 31872
rect 22612 31832 22618 31844
rect 18509 31807 18567 31813
rect 18509 31773 18521 31807
rect 18555 31804 18567 31807
rect 18598 31804 18604 31816
rect 18555 31776 18604 31804
rect 18555 31773 18567 31776
rect 18509 31767 18567 31773
rect 18598 31764 18604 31776
rect 18656 31764 18662 31816
rect 18966 31804 18972 31816
rect 18708 31776 18972 31804
rect 18233 31739 18291 31745
rect 18233 31705 18245 31739
rect 18279 31705 18291 31739
rect 18233 31699 18291 31705
rect 18598 31668 18604 31680
rect 17972 31640 18604 31668
rect 18598 31628 18604 31640
rect 18656 31628 18662 31680
rect 18708 31677 18736 31776
rect 18966 31764 18972 31776
rect 19024 31764 19030 31816
rect 20806 31764 20812 31816
rect 20864 31764 20870 31816
rect 22002 31764 22008 31816
rect 22060 31764 22066 31816
rect 22094 31764 22100 31816
rect 22152 31764 22158 31816
rect 22249 31807 22307 31813
rect 22249 31773 22261 31807
rect 22295 31804 22307 31807
rect 22295 31773 22324 31804
rect 22249 31767 22324 31773
rect 19426 31696 19432 31748
rect 19484 31736 19490 31748
rect 19705 31739 19763 31745
rect 19705 31736 19717 31739
rect 19484 31708 19717 31736
rect 19484 31696 19490 31708
rect 19705 31705 19717 31708
rect 19751 31705 19763 31739
rect 22020 31736 22048 31764
rect 22296 31736 22324 31767
rect 22370 31764 22376 31816
rect 22428 31804 22434 31816
rect 22428 31776 22473 31804
rect 22428 31764 22434 31776
rect 22738 31764 22744 31816
rect 22796 31804 22802 31816
rect 23676 31813 23704 31844
rect 23753 31841 23765 31875
rect 23799 31872 23811 31875
rect 23934 31872 23940 31884
rect 23799 31844 23940 31872
rect 23799 31841 23811 31844
rect 23753 31835 23811 31841
rect 23934 31832 23940 31844
rect 23992 31872 23998 31884
rect 25866 31872 25872 31884
rect 23992 31844 25872 31872
rect 23992 31832 23998 31844
rect 25866 31832 25872 31844
rect 25924 31832 25930 31884
rect 27157 31875 27215 31881
rect 27157 31841 27169 31875
rect 27203 31872 27215 31875
rect 27430 31872 27436 31884
rect 27203 31844 27436 31872
rect 27203 31841 27215 31844
rect 27157 31835 27215 31841
rect 27430 31832 27436 31844
rect 27488 31832 27494 31884
rect 28074 31832 28080 31884
rect 28132 31872 28138 31884
rect 28460 31872 28488 31912
rect 30006 31900 30012 31912
rect 30064 31900 30070 31952
rect 30742 31940 30748 31952
rect 30703 31912 30748 31940
rect 30742 31900 30748 31912
rect 30800 31900 30806 31952
rect 34146 31940 34152 31952
rect 31404 31912 31754 31940
rect 34107 31912 34152 31940
rect 28132 31844 28488 31872
rect 28132 31832 28138 31844
rect 28718 31832 28724 31884
rect 28776 31872 28782 31884
rect 28905 31875 28963 31881
rect 28905 31872 28917 31875
rect 28776 31844 28917 31872
rect 28776 31832 28782 31844
rect 28905 31841 28917 31844
rect 28951 31841 28963 31875
rect 29641 31875 29699 31881
rect 29641 31872 29653 31875
rect 28905 31835 28963 31841
rect 29104 31844 29653 31872
rect 23017 31807 23075 31813
rect 23017 31804 23029 31807
rect 22796 31776 23029 31804
rect 22796 31764 22802 31776
rect 23017 31773 23029 31776
rect 23063 31773 23075 31807
rect 23017 31767 23075 31773
rect 23661 31807 23719 31813
rect 23661 31773 23673 31807
rect 23707 31773 23719 31807
rect 23661 31767 23719 31773
rect 23842 31764 23848 31816
rect 23900 31804 23906 31816
rect 24949 31807 25007 31813
rect 23900 31776 23945 31804
rect 23900 31764 23906 31776
rect 24949 31773 24961 31807
rect 24995 31804 25007 31807
rect 25038 31804 25044 31816
rect 24995 31776 25044 31804
rect 24995 31773 25007 31776
rect 24949 31767 25007 31773
rect 25038 31764 25044 31776
rect 25096 31764 25102 31816
rect 29104 31804 29132 31844
rect 29641 31841 29653 31844
rect 29687 31841 29699 31875
rect 31018 31872 31024 31884
rect 29641 31835 29699 31841
rect 30380 31844 31024 31872
rect 28566 31776 29132 31804
rect 29362 31764 29368 31816
rect 29420 31764 29426 31816
rect 29546 31804 29552 31816
rect 29507 31776 29552 31804
rect 29546 31764 29552 31776
rect 29604 31764 29610 31816
rect 30380 31813 30408 31844
rect 31018 31832 31024 31844
rect 31076 31832 31082 31884
rect 31110 31832 31116 31884
rect 31168 31872 31174 31884
rect 31404 31872 31432 31912
rect 31168 31844 31432 31872
rect 31726 31872 31754 31912
rect 34146 31900 34152 31912
rect 34204 31900 34210 31952
rect 32401 31875 32459 31881
rect 32401 31872 32413 31875
rect 31726 31844 32413 31872
rect 31168 31832 31174 31844
rect 32401 31841 32413 31844
rect 32447 31841 32459 31875
rect 32401 31835 32459 31841
rect 32677 31875 32735 31881
rect 32677 31841 32689 31875
rect 32723 31872 32735 31875
rect 33134 31872 33140 31884
rect 32723 31844 33140 31872
rect 32723 31841 32735 31844
rect 32677 31835 32735 31841
rect 33134 31832 33140 31844
rect 33192 31832 33198 31884
rect 30377 31807 30435 31813
rect 29656 31776 30328 31804
rect 22020 31708 22324 31736
rect 27433 31739 27491 31745
rect 19705 31699 19763 31705
rect 27433 31705 27445 31739
rect 27479 31736 27491 31739
rect 27706 31736 27712 31748
rect 27479 31708 27712 31736
rect 27479 31705 27491 31708
rect 27433 31699 27491 31705
rect 27706 31696 27712 31708
rect 27764 31696 27770 31748
rect 29380 31736 29408 31764
rect 29656 31736 29684 31776
rect 29380 31708 29684 31736
rect 30300 31736 30328 31776
rect 30377 31773 30389 31807
rect 30423 31773 30435 31807
rect 30377 31767 30435 31773
rect 30466 31764 30472 31816
rect 30524 31804 30530 31816
rect 31294 31804 31300 31816
rect 30524 31776 30569 31804
rect 30668 31776 31156 31804
rect 31255 31776 31300 31804
rect 30524 31764 30530 31776
rect 30668 31736 30696 31776
rect 30300 31708 30696 31736
rect 31128 31736 31156 31776
rect 31294 31764 31300 31776
rect 31352 31764 31358 31816
rect 31570 31813 31576 31816
rect 31389 31807 31447 31813
rect 31389 31773 31401 31807
rect 31435 31804 31447 31807
rect 31527 31807 31576 31813
rect 31435 31776 31469 31804
rect 31435 31773 31447 31776
rect 31389 31767 31447 31773
rect 31527 31773 31539 31807
rect 31573 31773 31576 31807
rect 31527 31767 31576 31773
rect 31404 31736 31432 31767
rect 31570 31764 31576 31767
rect 31628 31764 31634 31816
rect 31665 31807 31723 31813
rect 31665 31773 31677 31807
rect 31711 31773 31723 31807
rect 31665 31767 31723 31773
rect 31128 31708 31432 31736
rect 18693 31671 18751 31677
rect 18693 31637 18705 31671
rect 18739 31637 18751 31671
rect 18693 31631 18751 31637
rect 21266 31628 21272 31680
rect 21324 31668 21330 31680
rect 22005 31671 22063 31677
rect 22005 31668 22017 31671
rect 21324 31640 22017 31668
rect 21324 31628 21330 31640
rect 22005 31637 22017 31640
rect 22051 31637 22063 31671
rect 22005 31631 22063 31637
rect 22094 31628 22100 31680
rect 22152 31668 22158 31680
rect 23109 31671 23167 31677
rect 23109 31668 23121 31671
rect 22152 31640 23121 31668
rect 22152 31628 22158 31640
rect 23109 31637 23121 31640
rect 23155 31637 23167 31671
rect 23109 31631 23167 31637
rect 25222 31628 25228 31680
rect 25280 31668 25286 31680
rect 29730 31668 29736 31680
rect 25280 31640 29736 31668
rect 25280 31628 25286 31640
rect 29730 31628 29736 31640
rect 29788 31628 29794 31680
rect 30742 31628 30748 31680
rect 30800 31668 30806 31680
rect 31680 31668 31708 31767
rect 33778 31764 33784 31816
rect 33836 31764 33842 31816
rect 30800 31640 31708 31668
rect 31757 31671 31815 31677
rect 30800 31628 30806 31640
rect 31757 31637 31769 31671
rect 31803 31668 31815 31671
rect 32398 31668 32404 31680
rect 31803 31640 32404 31668
rect 31803 31637 31815 31640
rect 31757 31631 31815 31637
rect 32398 31628 32404 31640
rect 32456 31628 32462 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 17126 31424 17132 31476
rect 17184 31464 17190 31476
rect 17313 31467 17371 31473
rect 17313 31464 17325 31467
rect 17184 31436 17325 31464
rect 17184 31424 17190 31436
rect 17313 31433 17325 31436
rect 17359 31433 17371 31467
rect 17862 31464 17868 31476
rect 17823 31436 17868 31464
rect 17313 31427 17371 31433
rect 17862 31424 17868 31436
rect 17920 31424 17926 31476
rect 19426 31424 19432 31476
rect 19484 31464 19490 31476
rect 19705 31467 19763 31473
rect 19705 31464 19717 31467
rect 19484 31436 19717 31464
rect 19484 31424 19490 31436
rect 19705 31433 19717 31436
rect 19751 31433 19763 31467
rect 19705 31427 19763 31433
rect 21450 31424 21456 31476
rect 21508 31464 21514 31476
rect 23569 31467 23627 31473
rect 23569 31464 23581 31467
rect 21508 31436 23581 31464
rect 21508 31424 21514 31436
rect 23569 31433 23581 31436
rect 23615 31464 23627 31467
rect 23842 31464 23848 31476
rect 23615 31436 23848 31464
rect 23615 31433 23627 31436
rect 23569 31427 23627 31433
rect 23842 31424 23848 31436
rect 23900 31424 23906 31476
rect 24394 31424 24400 31476
rect 24452 31464 24458 31476
rect 27154 31464 27160 31476
rect 24452 31436 27160 31464
rect 24452 31424 24458 31436
rect 27154 31424 27160 31436
rect 27212 31464 27218 31476
rect 27212 31436 27660 31464
rect 27212 31424 27218 31436
rect 1854 31356 1860 31408
rect 1912 31396 1918 31408
rect 2777 31399 2835 31405
rect 2777 31396 2789 31399
rect 1912 31368 2789 31396
rect 1912 31356 1918 31368
rect 2777 31365 2789 31368
rect 2823 31365 2835 31399
rect 2777 31359 2835 31365
rect 17037 31399 17095 31405
rect 17037 31365 17049 31399
rect 17083 31396 17095 31399
rect 18874 31396 18880 31408
rect 17083 31368 18880 31396
rect 17083 31365 17095 31368
rect 17037 31359 17095 31365
rect 18874 31356 18880 31368
rect 18932 31356 18938 31408
rect 19334 31396 19340 31408
rect 18984 31368 19340 31396
rect 15933 31331 15991 31337
rect 15933 31297 15945 31331
rect 15979 31297 15991 31331
rect 15933 31291 15991 31297
rect 16117 31331 16175 31337
rect 16117 31297 16129 31331
rect 16163 31328 16175 31331
rect 16574 31328 16580 31340
rect 16163 31300 16580 31328
rect 16163 31297 16175 31300
rect 16117 31291 16175 31297
rect 2590 31260 2596 31272
rect 2551 31232 2596 31260
rect 2590 31220 2596 31232
rect 2648 31220 2654 31272
rect 4433 31263 4491 31269
rect 4433 31229 4445 31263
rect 4479 31260 4491 31263
rect 4614 31260 4620 31272
rect 4479 31232 4620 31260
rect 4479 31229 4491 31232
rect 4433 31223 4491 31229
rect 4614 31220 4620 31232
rect 4672 31220 4678 31272
rect 6546 31084 6552 31136
rect 6604 31124 6610 31136
rect 6917 31127 6975 31133
rect 6917 31124 6929 31127
rect 6604 31096 6929 31124
rect 6604 31084 6610 31096
rect 6917 31093 6929 31096
rect 6963 31093 6975 31127
rect 15948 31124 15976 31291
rect 16574 31288 16580 31300
rect 16632 31288 16638 31340
rect 16669 31331 16727 31337
rect 16669 31297 16681 31331
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 16025 31263 16083 31269
rect 16025 31229 16037 31263
rect 16071 31260 16083 31263
rect 16684 31260 16712 31291
rect 16758 31288 16764 31340
rect 16816 31337 16822 31340
rect 16816 31331 16847 31337
rect 16835 31297 16847 31331
rect 16816 31291 16847 31297
rect 16945 31331 17003 31337
rect 16945 31297 16957 31331
rect 16991 31297 17003 31331
rect 16945 31291 17003 31297
rect 16816 31288 16822 31291
rect 16071 31232 16712 31260
rect 16960 31260 16988 31291
rect 17126 31288 17132 31340
rect 17184 31337 17190 31340
rect 18984 31337 19012 31368
rect 19334 31356 19340 31368
rect 19392 31356 19398 31408
rect 20901 31399 20959 31405
rect 20901 31365 20913 31399
rect 20947 31396 20959 31399
rect 22370 31396 22376 31408
rect 20947 31368 22376 31396
rect 20947 31365 20959 31368
rect 20901 31359 20959 31365
rect 22370 31356 22376 31368
rect 22428 31356 22434 31408
rect 22554 31356 22560 31408
rect 22612 31356 22618 31408
rect 27338 31356 27344 31408
rect 27396 31396 27402 31408
rect 27632 31396 27660 31436
rect 27706 31424 27712 31476
rect 27764 31464 27770 31476
rect 28077 31467 28135 31473
rect 28077 31464 28089 31467
rect 27764 31436 28089 31464
rect 27764 31424 27770 31436
rect 28077 31433 28089 31436
rect 28123 31433 28135 31467
rect 28902 31464 28908 31476
rect 28863 31436 28908 31464
rect 28077 31427 28135 31433
rect 28902 31424 28908 31436
rect 28960 31424 28966 31476
rect 33134 31464 33140 31476
rect 33095 31436 33140 31464
rect 33134 31424 33140 31436
rect 33192 31424 33198 31476
rect 33778 31464 33784 31476
rect 33739 31436 33784 31464
rect 33778 31424 33784 31436
rect 33836 31424 33842 31476
rect 46474 31424 46480 31476
rect 46532 31464 46538 31476
rect 46842 31464 46848 31476
rect 46532 31436 46848 31464
rect 46532 31424 46538 31436
rect 46842 31424 46848 31436
rect 46900 31424 46906 31476
rect 27801 31399 27859 31405
rect 27801 31396 27813 31399
rect 27396 31368 27568 31396
rect 27632 31368 27813 31396
rect 27396 31356 27402 31368
rect 17184 31328 17192 31337
rect 17773 31331 17831 31337
rect 17184 31300 17229 31328
rect 17184 31291 17192 31300
rect 17773 31297 17785 31331
rect 17819 31297 17831 31331
rect 17773 31291 17831 31297
rect 18969 31331 19027 31337
rect 18969 31297 18981 31331
rect 19015 31297 19027 31331
rect 18969 31291 19027 31297
rect 19153 31331 19211 31337
rect 19153 31297 19165 31331
rect 19199 31330 19211 31331
rect 19199 31328 19288 31330
rect 19426 31328 19432 31340
rect 19199 31302 19432 31328
rect 19199 31297 19211 31302
rect 19260 31300 19432 31302
rect 19153 31291 19211 31297
rect 17184 31288 17190 31291
rect 16960 31232 17724 31260
rect 16071 31229 16083 31232
rect 16025 31223 16083 31229
rect 17218 31124 17224 31136
rect 15948 31096 17224 31124
rect 6917 31087 6975 31093
rect 17218 31084 17224 31096
rect 17276 31084 17282 31136
rect 17696 31124 17724 31232
rect 17788 31192 17816 31291
rect 19426 31288 19432 31300
rect 19484 31288 19490 31340
rect 19521 31331 19579 31337
rect 19521 31297 19533 31331
rect 19567 31328 19579 31331
rect 20530 31328 20536 31340
rect 19567 31300 20536 31328
rect 19567 31297 19579 31300
rect 19521 31291 19579 31297
rect 20530 31288 20536 31300
rect 20588 31288 20594 31340
rect 24578 31288 24584 31340
rect 24636 31328 24642 31340
rect 24673 31331 24731 31337
rect 24673 31328 24685 31331
rect 24636 31300 24685 31328
rect 24636 31288 24642 31300
rect 24673 31297 24685 31300
rect 24719 31297 24731 31331
rect 25498 31328 25504 31340
rect 25459 31300 25504 31328
rect 24673 31291 24731 31297
rect 25498 31288 25504 31300
rect 25556 31288 25562 31340
rect 27540 31337 27568 31368
rect 27801 31365 27813 31368
rect 27847 31365 27859 31399
rect 27801 31359 27859 31365
rect 31202 31356 31208 31408
rect 31260 31396 31266 31408
rect 31260 31368 32996 31396
rect 31260 31356 31266 31368
rect 32968 31340 32996 31368
rect 27433 31331 27491 31337
rect 27433 31297 27445 31331
rect 27479 31297 27491 31331
rect 27433 31291 27491 31297
rect 27526 31331 27584 31337
rect 27526 31297 27538 31331
rect 27572 31297 27584 31331
rect 27526 31291 27584 31297
rect 19242 31260 19248 31272
rect 19203 31232 19248 31260
rect 19242 31220 19248 31232
rect 19300 31220 19306 31272
rect 19337 31263 19395 31269
rect 19337 31229 19349 31263
rect 19383 31260 19395 31263
rect 19978 31260 19984 31272
rect 19383 31232 19984 31260
rect 19383 31229 19395 31232
rect 19337 31223 19395 31229
rect 19978 31220 19984 31232
rect 20036 31220 20042 31272
rect 21821 31263 21879 31269
rect 21821 31229 21833 31263
rect 21867 31229 21879 31263
rect 21821 31223 21879 31229
rect 22097 31263 22155 31269
rect 22097 31229 22109 31263
rect 22143 31260 22155 31263
rect 22186 31260 22192 31272
rect 22143 31232 22192 31260
rect 22143 31229 22155 31232
rect 22097 31223 22155 31229
rect 20898 31192 20904 31204
rect 17788 31164 20904 31192
rect 20898 31152 20904 31164
rect 20956 31192 20962 31204
rect 21085 31195 21143 31201
rect 21085 31192 21097 31195
rect 20956 31164 21097 31192
rect 20956 31152 20962 31164
rect 21085 31161 21097 31164
rect 21131 31161 21143 31195
rect 21085 31155 21143 31161
rect 20990 31124 20996 31136
rect 17696 31096 20996 31124
rect 20990 31084 20996 31096
rect 21048 31084 21054 31136
rect 21836 31124 21864 31223
rect 22186 31220 22192 31232
rect 22244 31220 22250 31272
rect 24765 31263 24823 31269
rect 24765 31229 24777 31263
rect 24811 31260 24823 31263
rect 24854 31260 24860 31272
rect 24811 31232 24860 31260
rect 24811 31229 24823 31232
rect 24765 31223 24823 31229
rect 24854 31220 24860 31232
rect 24912 31220 24918 31272
rect 25041 31263 25099 31269
rect 25041 31229 25053 31263
rect 25087 31260 25099 31263
rect 25406 31260 25412 31272
rect 25087 31232 25412 31260
rect 25087 31229 25099 31232
rect 25041 31223 25099 31229
rect 25406 31220 25412 31232
rect 25464 31220 25470 31272
rect 27448 31260 27476 31291
rect 27614 31288 27620 31340
rect 27672 31328 27678 31340
rect 27709 31331 27767 31337
rect 27709 31328 27721 31331
rect 27672 31300 27721 31328
rect 27672 31288 27678 31300
rect 27709 31297 27721 31300
rect 27755 31297 27767 31331
rect 27709 31291 27767 31297
rect 27939 31331 27997 31337
rect 27939 31297 27951 31331
rect 27985 31328 27997 31331
rect 28626 31328 28632 31340
rect 27985 31300 28632 31328
rect 27985 31297 27997 31300
rect 27939 31291 27997 31297
rect 28626 31288 28632 31300
rect 28684 31288 28690 31340
rect 28810 31328 28816 31340
rect 28771 31300 28816 31328
rect 28810 31288 28816 31300
rect 28868 31288 28874 31340
rect 28994 31328 29000 31340
rect 28955 31300 29000 31328
rect 28994 31288 29000 31300
rect 29052 31288 29058 31340
rect 30834 31288 30840 31340
rect 30892 31328 30898 31340
rect 31021 31331 31079 31337
rect 31021 31328 31033 31331
rect 30892 31300 31033 31328
rect 30892 31288 30898 31300
rect 31021 31297 31033 31300
rect 31067 31297 31079 31331
rect 32398 31328 32404 31340
rect 32359 31300 32404 31328
rect 31021 31291 31079 31297
rect 32398 31288 32404 31300
rect 32456 31288 32462 31340
rect 32582 31328 32588 31340
rect 32543 31300 32588 31328
rect 32582 31288 32588 31300
rect 32640 31288 32646 31340
rect 32674 31288 32680 31340
rect 32732 31328 32738 31340
rect 32950 31328 32956 31340
rect 32732 31300 32777 31328
rect 32863 31300 32956 31328
rect 32732 31288 32738 31300
rect 32950 31288 32956 31300
rect 33008 31288 33014 31340
rect 33686 31328 33692 31340
rect 33647 31300 33692 31328
rect 33686 31288 33692 31300
rect 33744 31288 33750 31340
rect 28258 31260 28264 31272
rect 27448 31232 28264 31260
rect 28258 31220 28264 31232
rect 28316 31220 28322 31272
rect 30466 31220 30472 31272
rect 30524 31260 30530 31272
rect 30745 31263 30803 31269
rect 30745 31260 30757 31263
rect 30524 31232 30757 31260
rect 30524 31220 30530 31232
rect 30745 31229 30757 31232
rect 30791 31260 30803 31263
rect 31110 31260 31116 31272
rect 30791 31232 31116 31260
rect 30791 31229 30803 31232
rect 30745 31223 30803 31229
rect 31110 31220 31116 31232
rect 31168 31220 31174 31272
rect 32490 31220 32496 31272
rect 32548 31260 32554 31272
rect 32769 31263 32827 31269
rect 32769 31260 32781 31263
rect 32548 31232 32781 31260
rect 32548 31220 32554 31232
rect 32769 31229 32781 31232
rect 32815 31229 32827 31263
rect 32769 31223 32827 31229
rect 22094 31124 22100 31136
rect 21836 31096 22100 31124
rect 22094 31084 22100 31096
rect 22152 31084 22158 31136
rect 25685 31127 25743 31133
rect 25685 31093 25697 31127
rect 25731 31124 25743 31127
rect 25866 31124 25872 31136
rect 25731 31096 25872 31124
rect 25731 31093 25743 31096
rect 25685 31087 25743 31093
rect 25866 31084 25872 31096
rect 25924 31084 25930 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 16574 30880 16580 30932
rect 16632 30920 16638 30932
rect 20898 30920 20904 30932
rect 16632 30892 20904 30920
rect 16632 30880 16638 30892
rect 20898 30880 20904 30892
rect 20956 30880 20962 30932
rect 21913 30923 21971 30929
rect 21913 30889 21925 30923
rect 21959 30920 21971 30923
rect 22186 30920 22192 30932
rect 21959 30892 22192 30920
rect 21959 30889 21971 30892
rect 21913 30883 21971 30889
rect 22186 30880 22192 30892
rect 22244 30880 22250 30932
rect 22465 30923 22523 30929
rect 22465 30889 22477 30923
rect 22511 30920 22523 30923
rect 22554 30920 22560 30932
rect 22511 30892 22560 30920
rect 22511 30889 22523 30892
rect 22465 30883 22523 30889
rect 22554 30880 22560 30892
rect 22612 30880 22618 30932
rect 24581 30923 24639 30929
rect 24581 30889 24593 30923
rect 24627 30920 24639 30923
rect 24670 30920 24676 30932
rect 24627 30892 24676 30920
rect 24627 30889 24639 30892
rect 24581 30883 24639 30889
rect 21634 30812 21640 30864
rect 21692 30852 21698 30864
rect 22002 30852 22008 30864
rect 21692 30824 22008 30852
rect 21692 30812 21698 30824
rect 22002 30812 22008 30824
rect 22060 30812 22066 30864
rect 6546 30784 6552 30796
rect 6507 30756 6552 30784
rect 6546 30744 6552 30756
rect 6604 30744 6610 30796
rect 6733 30787 6791 30793
rect 6733 30753 6745 30787
rect 6779 30784 6791 30787
rect 7558 30784 7564 30796
rect 6779 30756 7564 30784
rect 6779 30753 6791 30756
rect 6733 30747 6791 30753
rect 7558 30744 7564 30756
rect 7616 30744 7622 30796
rect 8202 30784 8208 30796
rect 8163 30756 8208 30784
rect 8202 30744 8208 30756
rect 8260 30744 8266 30796
rect 20990 30744 20996 30796
rect 21048 30784 21054 30796
rect 24596 30784 24624 30883
rect 24670 30880 24676 30892
rect 24728 30880 24734 30932
rect 25317 30923 25375 30929
rect 25317 30889 25329 30923
rect 25363 30889 25375 30923
rect 25498 30920 25504 30932
rect 25459 30892 25504 30920
rect 25317 30883 25375 30889
rect 25332 30852 25360 30883
rect 25498 30880 25504 30892
rect 25556 30880 25562 30932
rect 30190 30920 30196 30932
rect 30151 30892 30196 30920
rect 30190 30880 30196 30892
rect 30248 30880 30254 30932
rect 30745 30923 30803 30929
rect 30745 30889 30757 30923
rect 30791 30920 30803 30923
rect 30834 30920 30840 30932
rect 30791 30892 30840 30920
rect 30791 30889 30803 30892
rect 30745 30883 30803 30889
rect 30834 30880 30840 30892
rect 30892 30880 30898 30932
rect 26237 30855 26295 30861
rect 25332 30824 26096 30852
rect 26068 30784 26096 30824
rect 26237 30821 26249 30855
rect 26283 30852 26295 30855
rect 26326 30852 26332 30864
rect 26283 30824 26332 30852
rect 26283 30821 26295 30824
rect 26237 30815 26295 30821
rect 26326 30812 26332 30824
rect 26384 30812 26390 30864
rect 26970 30852 26976 30864
rect 26883 30824 26976 30852
rect 26970 30812 26976 30824
rect 27028 30852 27034 30864
rect 32582 30852 32588 30864
rect 27028 30824 32588 30852
rect 27028 30812 27034 30824
rect 28813 30787 28871 30793
rect 28813 30784 28825 30787
rect 21048 30756 21588 30784
rect 21048 30744 21054 30756
rect 21266 30716 21272 30728
rect 21227 30688 21272 30716
rect 21266 30676 21272 30688
rect 21324 30676 21330 30728
rect 21450 30725 21456 30728
rect 21417 30719 21456 30725
rect 21417 30685 21429 30719
rect 21417 30679 21456 30685
rect 21450 30676 21456 30679
rect 21508 30676 21514 30728
rect 21560 30725 21588 30756
rect 22388 30756 24624 30784
rect 24964 30756 25360 30784
rect 21545 30719 21603 30725
rect 21545 30685 21557 30719
rect 21591 30685 21603 30719
rect 21545 30679 21603 30685
rect 21726 30676 21732 30728
rect 21784 30725 21790 30728
rect 22388 30725 22416 30756
rect 21784 30716 21792 30725
rect 22373 30719 22431 30725
rect 21784 30688 21829 30716
rect 21784 30679 21792 30688
rect 22373 30685 22385 30719
rect 22419 30685 22431 30719
rect 22373 30679 22431 30685
rect 21784 30676 21790 30679
rect 22554 30676 22560 30728
rect 22612 30716 22618 30728
rect 24397 30719 24455 30725
rect 24397 30716 24409 30719
rect 22612 30688 24409 30716
rect 22612 30676 22618 30688
rect 24397 30685 24409 30688
rect 24443 30716 24455 30719
rect 24964 30716 24992 30756
rect 25222 30716 25228 30728
rect 24443 30688 24992 30716
rect 25056 30688 25228 30716
rect 24443 30685 24455 30688
rect 24397 30679 24455 30685
rect 18874 30608 18880 30660
rect 18932 30648 18938 30660
rect 21637 30651 21695 30657
rect 21637 30648 21649 30651
rect 18932 30620 21649 30648
rect 18932 30608 18938 30620
rect 21637 30617 21649 30620
rect 21683 30648 21695 30651
rect 25056 30648 25084 30688
rect 25222 30676 25228 30688
rect 25280 30676 25286 30728
rect 25332 30716 25360 30756
rect 26068 30756 28825 30784
rect 26068 30725 26096 30756
rect 28813 30753 28825 30756
rect 28859 30753 28871 30787
rect 28813 30747 28871 30753
rect 30282 30744 30288 30796
rect 30340 30784 30346 30796
rect 30929 30787 30987 30793
rect 30929 30784 30941 30787
rect 30340 30756 30941 30784
rect 30340 30744 30346 30756
rect 30929 30753 30941 30756
rect 30975 30753 30987 30787
rect 30929 30747 30987 30753
rect 26053 30719 26111 30725
rect 25332 30688 26004 30716
rect 21683 30620 25084 30648
rect 25133 30651 25191 30657
rect 21683 30617 21695 30620
rect 21637 30611 21695 30617
rect 25133 30617 25145 30651
rect 25179 30617 25191 30651
rect 25133 30611 25191 30617
rect 25148 30580 25176 30611
rect 25314 30608 25320 30660
rect 25372 30657 25378 30660
rect 25372 30651 25391 30657
rect 25379 30617 25391 30651
rect 25976 30648 26004 30688
rect 26053 30685 26065 30719
rect 26099 30685 26111 30719
rect 27985 30719 28043 30725
rect 27985 30716 27997 30719
rect 26053 30679 26111 30685
rect 26160 30688 27997 30716
rect 26160 30648 26188 30688
rect 27985 30685 27997 30688
rect 28031 30685 28043 30719
rect 27985 30679 28043 30685
rect 28534 30676 28540 30728
rect 28592 30716 28598 30728
rect 28721 30719 28779 30725
rect 28721 30716 28733 30719
rect 28592 30688 28733 30716
rect 28592 30676 28598 30688
rect 28721 30685 28733 30688
rect 28767 30685 28779 30719
rect 28721 30679 28779 30685
rect 28994 30676 29000 30728
rect 29052 30716 29058 30728
rect 30009 30719 30067 30725
rect 30009 30716 30021 30719
rect 29052 30688 30021 30716
rect 29052 30676 29058 30688
rect 30009 30685 30021 30688
rect 30055 30685 30067 30719
rect 30650 30716 30656 30728
rect 30611 30688 30656 30716
rect 30009 30679 30067 30685
rect 30650 30676 30656 30688
rect 30708 30676 30714 30728
rect 32398 30716 32404 30728
rect 32359 30688 32404 30716
rect 32398 30676 32404 30688
rect 32456 30676 32462 30728
rect 32508 30716 32536 30824
rect 32582 30812 32588 30824
rect 32640 30812 32646 30864
rect 32769 30787 32827 30793
rect 32769 30753 32781 30787
rect 32815 30784 32827 30787
rect 40402 30784 40408 30796
rect 32815 30756 40408 30784
rect 32815 30753 32827 30756
rect 32769 30747 32827 30753
rect 40402 30744 40408 30756
rect 40460 30744 40466 30796
rect 47026 30744 47032 30796
rect 47084 30784 47090 30796
rect 47121 30787 47179 30793
rect 47121 30784 47133 30787
rect 47084 30756 47133 30784
rect 47084 30744 47090 30756
rect 47121 30753 47133 30756
rect 47167 30784 47179 30787
rect 47670 30784 47676 30796
rect 47167 30756 47676 30784
rect 47167 30753 47179 30756
rect 47121 30747 47179 30753
rect 47670 30744 47676 30756
rect 47728 30744 47734 30796
rect 32585 30719 32643 30725
rect 32585 30716 32597 30719
rect 32508 30688 32597 30716
rect 32585 30685 32597 30688
rect 32631 30685 32643 30719
rect 32585 30679 32643 30685
rect 32674 30676 32680 30728
rect 32732 30716 32738 30728
rect 32950 30716 32956 30728
rect 32732 30688 32777 30716
rect 32911 30688 32956 30716
rect 32732 30676 32738 30688
rect 32950 30676 32956 30688
rect 33008 30676 33014 30728
rect 25976 30620 26188 30648
rect 25372 30611 25391 30617
rect 25372 30608 25378 30611
rect 26510 30608 26516 30660
rect 26568 30648 26574 30660
rect 26786 30648 26792 30660
rect 26568 30620 26792 30648
rect 26568 30608 26574 30620
rect 26786 30608 26792 30620
rect 26844 30608 26850 30660
rect 29825 30651 29883 30657
rect 29825 30617 29837 30651
rect 29871 30648 29883 30651
rect 30282 30648 30288 30660
rect 29871 30620 30288 30648
rect 29871 30617 29883 30620
rect 29825 30611 29883 30617
rect 30282 30608 30288 30620
rect 30340 30608 30346 30660
rect 46014 30608 46020 30660
rect 46072 30648 46078 30660
rect 46845 30651 46903 30657
rect 46845 30648 46857 30651
rect 46072 30620 46857 30648
rect 46072 30608 46078 30620
rect 46845 30617 46857 30620
rect 46891 30617 46903 30651
rect 46845 30611 46903 30617
rect 46937 30651 46995 30657
rect 46937 30617 46949 30651
rect 46983 30648 46995 30651
rect 47762 30648 47768 30660
rect 46983 30620 47768 30648
rect 46983 30617 46995 30620
rect 46937 30611 46995 30617
rect 47762 30608 47768 30620
rect 47820 30608 47826 30660
rect 25590 30580 25596 30592
rect 25148 30552 25596 30580
rect 25590 30540 25596 30552
rect 25648 30580 25654 30592
rect 25958 30580 25964 30592
rect 25648 30552 25964 30580
rect 25648 30540 25654 30552
rect 25958 30540 25964 30552
rect 26016 30540 26022 30592
rect 28169 30583 28227 30589
rect 28169 30549 28181 30583
rect 28215 30580 28227 30583
rect 28258 30580 28264 30592
rect 28215 30552 28264 30580
rect 28215 30549 28227 30552
rect 28169 30543 28227 30549
rect 28258 30540 28264 30552
rect 28316 30540 28322 30592
rect 30374 30540 30380 30592
rect 30432 30580 30438 30592
rect 30929 30583 30987 30589
rect 30929 30580 30941 30583
rect 30432 30552 30941 30580
rect 30432 30540 30438 30552
rect 30929 30549 30941 30552
rect 30975 30549 30987 30583
rect 33134 30580 33140 30592
rect 33095 30552 33140 30580
rect 30929 30543 30987 30549
rect 33134 30540 33140 30552
rect 33192 30540 33198 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 20162 30376 20168 30388
rect 19484 30348 20168 30376
rect 19484 30336 19490 30348
rect 20162 30336 20168 30348
rect 20220 30376 20226 30388
rect 28442 30376 28448 30388
rect 20220 30348 22324 30376
rect 20220 30336 20226 30348
rect 17954 30268 17960 30320
rect 18012 30268 18018 30320
rect 16850 30200 16856 30252
rect 16908 30240 16914 30252
rect 16945 30243 17003 30249
rect 16945 30240 16957 30243
rect 16908 30212 16957 30240
rect 16908 30200 16914 30212
rect 16945 30209 16957 30212
rect 16991 30209 17003 30243
rect 16945 30203 17003 30209
rect 19058 30200 19064 30252
rect 19116 30240 19122 30252
rect 19245 30243 19303 30249
rect 19245 30240 19257 30243
rect 19116 30212 19257 30240
rect 19116 30200 19122 30212
rect 19245 30209 19257 30212
rect 19291 30209 19303 30243
rect 19426 30240 19432 30252
rect 19387 30212 19432 30240
rect 19245 30203 19303 30209
rect 19426 30200 19432 30212
rect 19484 30200 19490 30252
rect 19613 30243 19671 30249
rect 19613 30209 19625 30243
rect 19659 30209 19671 30243
rect 19613 30203 19671 30209
rect 17221 30175 17279 30181
rect 17221 30141 17233 30175
rect 17267 30172 17279 30175
rect 19518 30172 19524 30184
rect 17267 30144 18644 30172
rect 19479 30144 19524 30172
rect 17267 30141 17279 30144
rect 17221 30135 17279 30141
rect 18616 30104 18644 30144
rect 19518 30132 19524 30144
rect 19576 30132 19582 30184
rect 19628 30172 19656 30203
rect 19794 30200 19800 30252
rect 19852 30240 19858 30252
rect 19852 30212 19897 30240
rect 19852 30200 19858 30212
rect 20070 30172 20076 30184
rect 19628 30144 20076 30172
rect 20070 30132 20076 30144
rect 20128 30132 20134 30184
rect 19981 30107 20039 30113
rect 19981 30104 19993 30107
rect 18616 30076 19993 30104
rect 19981 30073 19993 30076
rect 20027 30073 20039 30107
rect 22296 30104 22324 30348
rect 27540 30348 28448 30376
rect 27540 30317 27568 30348
rect 28442 30336 28448 30348
rect 28500 30336 28506 30388
rect 28810 30336 28816 30388
rect 28868 30376 28874 30388
rect 29641 30379 29699 30385
rect 28868 30348 29040 30376
rect 28868 30336 28874 30348
rect 27525 30311 27583 30317
rect 25332 30280 26096 30308
rect 25332 30252 25360 30280
rect 24121 30243 24179 30249
rect 24121 30209 24133 30243
rect 24167 30209 24179 30243
rect 24854 30240 24860 30252
rect 24767 30212 24860 30240
rect 24121 30203 24179 30209
rect 24136 30172 24164 30203
rect 24854 30200 24860 30212
rect 24912 30240 24918 30252
rect 25314 30240 25320 30252
rect 24912 30212 25320 30240
rect 24912 30200 24918 30212
rect 25314 30200 25320 30212
rect 25372 30200 25378 30252
rect 25498 30200 25504 30252
rect 25556 30240 25562 30252
rect 25777 30243 25835 30249
rect 25777 30240 25789 30243
rect 25556 30212 25789 30240
rect 25556 30200 25562 30212
rect 25777 30209 25789 30212
rect 25823 30209 25835 30243
rect 25958 30240 25964 30252
rect 25919 30212 25964 30240
rect 25777 30203 25835 30209
rect 25958 30200 25964 30212
rect 26016 30200 26022 30252
rect 26068 30249 26096 30280
rect 27525 30277 27537 30311
rect 27571 30277 27583 30311
rect 28902 30308 28908 30320
rect 27525 30271 27583 30277
rect 28460 30280 28908 30308
rect 26053 30243 26111 30249
rect 26053 30209 26065 30243
rect 26099 30209 26111 30243
rect 26053 30203 26111 30209
rect 27798 30200 27804 30252
rect 27856 30240 27862 30252
rect 28460 30249 28488 30280
rect 28902 30268 28908 30280
rect 28960 30268 28966 30320
rect 29012 30308 29040 30348
rect 29641 30345 29653 30379
rect 29687 30376 29699 30379
rect 29730 30376 29736 30388
rect 29687 30348 29736 30376
rect 29687 30345 29699 30348
rect 29641 30339 29699 30345
rect 29730 30336 29736 30348
rect 29788 30336 29794 30388
rect 30561 30379 30619 30385
rect 30561 30345 30573 30379
rect 30607 30345 30619 30379
rect 30561 30339 30619 30345
rect 30576 30308 30604 30339
rect 47762 30336 47768 30388
rect 47820 30376 47826 30388
rect 48222 30376 48228 30388
rect 47820 30348 48228 30376
rect 47820 30336 47826 30348
rect 48222 30336 48228 30348
rect 48280 30336 48286 30388
rect 33134 30308 33140 30320
rect 29012 30280 30604 30308
rect 33095 30280 33140 30308
rect 33134 30268 33140 30280
rect 33192 30268 33198 30320
rect 33778 30268 33784 30320
rect 33836 30268 33842 30320
rect 28353 30243 28411 30249
rect 28353 30240 28365 30243
rect 27856 30212 28365 30240
rect 27856 30200 27862 30212
rect 28353 30209 28365 30212
rect 28399 30209 28411 30243
rect 28353 30203 28411 30209
rect 28445 30243 28503 30249
rect 28445 30209 28457 30243
rect 28491 30209 28503 30243
rect 28445 30203 28503 30209
rect 28721 30243 28779 30249
rect 28721 30209 28733 30243
rect 28767 30240 28779 30243
rect 28994 30240 29000 30252
rect 28767 30212 29000 30240
rect 28767 30209 28779 30212
rect 28721 30203 28779 30209
rect 28994 30200 29000 30212
rect 29052 30200 29058 30252
rect 29454 30240 29460 30252
rect 29415 30212 29460 30240
rect 29454 30200 29460 30212
rect 29512 30200 29518 30252
rect 29638 30200 29644 30252
rect 29696 30240 29702 30252
rect 29914 30240 29920 30252
rect 29696 30212 29920 30240
rect 29696 30200 29702 30212
rect 29914 30200 29920 30212
rect 29972 30200 29978 30252
rect 30193 30243 30251 30249
rect 30193 30209 30205 30243
rect 30239 30240 30251 30243
rect 30834 30240 30840 30252
rect 30239 30212 30840 30240
rect 30239 30209 30251 30212
rect 30193 30203 30251 30209
rect 30834 30200 30840 30212
rect 30892 30240 30898 30252
rect 31021 30243 31079 30249
rect 31021 30240 31033 30243
rect 30892 30212 31033 30240
rect 30892 30200 30898 30212
rect 31021 30209 31033 30212
rect 31067 30209 31079 30243
rect 31021 30203 31079 30209
rect 25406 30172 25412 30184
rect 24136 30144 25412 30172
rect 25406 30132 25412 30144
rect 25464 30132 25470 30184
rect 25593 30175 25651 30181
rect 25593 30141 25605 30175
rect 25639 30172 25651 30175
rect 26786 30172 26792 30184
rect 25639 30144 26792 30172
rect 25639 30141 25651 30144
rect 25593 30135 25651 30141
rect 26786 30132 26792 30144
rect 26844 30172 26850 30184
rect 28629 30175 28687 30181
rect 28629 30172 28641 30175
rect 26844 30144 28641 30172
rect 26844 30132 26850 30144
rect 28629 30141 28641 30144
rect 28675 30141 28687 30175
rect 28629 30135 28687 30141
rect 30006 30132 30012 30184
rect 30064 30172 30070 30184
rect 30282 30172 30288 30184
rect 30064 30144 30288 30172
rect 30064 30132 30070 30144
rect 30282 30132 30288 30144
rect 30340 30132 30346 30184
rect 31294 30172 31300 30184
rect 31255 30144 31300 30172
rect 31294 30132 31300 30144
rect 31352 30132 31358 30184
rect 32858 30172 32864 30184
rect 32819 30144 32864 30172
rect 32858 30132 32864 30144
rect 32916 30132 32922 30184
rect 24305 30107 24363 30113
rect 24305 30104 24317 30107
rect 22296 30076 24317 30104
rect 19981 30067 20039 30073
rect 24305 30073 24317 30076
rect 24351 30104 24363 30107
rect 29086 30104 29092 30116
rect 24351 30076 29092 30104
rect 24351 30073 24363 30076
rect 24305 30067 24363 30073
rect 29086 30064 29092 30076
rect 29144 30064 29150 30116
rect 31573 30107 31631 30113
rect 31573 30073 31585 30107
rect 31619 30104 31631 30107
rect 32398 30104 32404 30116
rect 31619 30076 32404 30104
rect 31619 30073 31631 30076
rect 31573 30067 31631 30073
rect 32398 30064 32404 30076
rect 32456 30064 32462 30116
rect 18693 30039 18751 30045
rect 18693 30005 18705 30039
rect 18739 30036 18751 30039
rect 19794 30036 19800 30048
rect 18739 30008 19800 30036
rect 18739 30005 18751 30008
rect 18693 29999 18751 30005
rect 19794 29996 19800 30008
rect 19852 29996 19858 30048
rect 25041 30039 25099 30045
rect 25041 30005 25053 30039
rect 25087 30036 25099 30039
rect 25314 30036 25320 30048
rect 25087 30008 25320 30036
rect 25087 30005 25099 30008
rect 25041 29999 25099 30005
rect 25314 29996 25320 30008
rect 25372 30036 25378 30048
rect 25774 30036 25780 30048
rect 25372 30008 25780 30036
rect 25372 29996 25378 30008
rect 25774 29996 25780 30008
rect 25832 29996 25838 30048
rect 27430 29996 27436 30048
rect 27488 30036 27494 30048
rect 27617 30039 27675 30045
rect 27617 30036 27629 30039
rect 27488 30008 27629 30036
rect 27488 29996 27494 30008
rect 27617 30005 27629 30008
rect 27663 30005 27675 30039
rect 27617 29999 27675 30005
rect 27706 29996 27712 30048
rect 27764 30036 27770 30048
rect 28169 30039 28227 30045
rect 28169 30036 28181 30039
rect 27764 30008 28181 30036
rect 27764 29996 27770 30008
rect 28169 30005 28181 30008
rect 28215 30005 28227 30039
rect 28169 29999 28227 30005
rect 30377 30039 30435 30045
rect 30377 30005 30389 30039
rect 30423 30036 30435 30039
rect 30650 30036 30656 30048
rect 30423 30008 30656 30036
rect 30423 30005 30435 30008
rect 30377 29999 30435 30005
rect 30650 29996 30656 30008
rect 30708 29996 30714 30048
rect 31386 30036 31392 30048
rect 31347 30008 31392 30036
rect 31386 29996 31392 30008
rect 31444 29996 31450 30048
rect 31754 29996 31760 30048
rect 31812 30036 31818 30048
rect 32674 30036 32680 30048
rect 31812 30008 32680 30036
rect 31812 29996 31818 30008
rect 32674 29996 32680 30008
rect 32732 30036 32738 30048
rect 34609 30039 34667 30045
rect 34609 30036 34621 30039
rect 32732 30008 34621 30036
rect 32732 29996 32738 30008
rect 34609 30005 34621 30008
rect 34655 30005 34667 30039
rect 34609 29999 34667 30005
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 17954 29792 17960 29844
rect 18012 29832 18018 29844
rect 18049 29835 18107 29841
rect 18049 29832 18061 29835
rect 18012 29804 18061 29832
rect 18012 29792 18018 29804
rect 18049 29801 18061 29804
rect 18095 29801 18107 29835
rect 18049 29795 18107 29801
rect 19518 29792 19524 29844
rect 19576 29832 19582 29844
rect 19705 29835 19763 29841
rect 19705 29832 19717 29835
rect 19576 29804 19717 29832
rect 19576 29792 19582 29804
rect 19705 29801 19717 29804
rect 19751 29801 19763 29835
rect 19705 29795 19763 29801
rect 19978 29792 19984 29844
rect 20036 29832 20042 29844
rect 20533 29835 20591 29841
rect 20533 29832 20545 29835
rect 20036 29804 20545 29832
rect 20036 29792 20042 29804
rect 20533 29801 20545 29804
rect 20579 29801 20591 29835
rect 20533 29795 20591 29801
rect 22646 29792 22652 29844
rect 22704 29832 22710 29844
rect 28813 29835 28871 29841
rect 22704 29804 28396 29832
rect 22704 29792 22710 29804
rect 28368 29764 28396 29804
rect 28813 29801 28825 29835
rect 28859 29832 28871 29835
rect 28994 29832 29000 29844
rect 28859 29804 29000 29832
rect 28859 29801 28871 29804
rect 28813 29795 28871 29801
rect 28994 29792 29000 29804
rect 29052 29792 29058 29844
rect 29914 29832 29920 29844
rect 29875 29804 29920 29832
rect 29914 29792 29920 29804
rect 29972 29792 29978 29844
rect 30190 29792 30196 29844
rect 30248 29832 30254 29844
rect 31294 29832 31300 29844
rect 30248 29804 31300 29832
rect 30248 29792 30254 29804
rect 31294 29792 31300 29804
rect 31352 29792 31358 29844
rect 33778 29832 33784 29844
rect 33739 29804 33784 29832
rect 33778 29792 33784 29804
rect 33836 29792 33842 29844
rect 29932 29764 29960 29792
rect 28368 29736 29960 29764
rect 19518 29696 19524 29708
rect 19479 29668 19524 29696
rect 19518 29656 19524 29668
rect 19576 29656 19582 29708
rect 20346 29656 20352 29708
rect 20404 29696 20410 29708
rect 24765 29699 24823 29705
rect 20404 29668 24716 29696
rect 20404 29656 20410 29668
rect 17957 29631 18015 29637
rect 17957 29597 17969 29631
rect 18003 29628 18015 29631
rect 18138 29628 18144 29640
rect 18003 29600 18144 29628
rect 18003 29597 18015 29600
rect 17957 29591 18015 29597
rect 18138 29588 18144 29600
rect 18196 29588 18202 29640
rect 19429 29631 19487 29637
rect 19429 29597 19441 29631
rect 19475 29628 19487 29631
rect 19794 29628 19800 29640
rect 19475 29600 19800 29628
rect 19475 29597 19487 29600
rect 19429 29591 19487 29597
rect 19794 29588 19800 29600
rect 19852 29628 19858 29640
rect 20070 29628 20076 29640
rect 19852 29600 20076 29628
rect 19852 29588 19858 29600
rect 20070 29588 20076 29600
rect 20128 29588 20134 29640
rect 20441 29631 20499 29637
rect 20441 29597 20453 29631
rect 20487 29597 20499 29631
rect 20714 29628 20720 29640
rect 20675 29600 20720 29628
rect 20441 29591 20499 29597
rect 20456 29560 20484 29591
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 24489 29631 24547 29637
rect 24489 29597 24501 29631
rect 24535 29628 24547 29631
rect 24578 29628 24584 29640
rect 24535 29600 24584 29628
rect 24535 29597 24547 29600
rect 24489 29591 24547 29597
rect 24578 29588 24584 29600
rect 24636 29588 24642 29640
rect 24688 29628 24716 29668
rect 24765 29665 24777 29699
rect 24811 29696 24823 29699
rect 24854 29696 24860 29708
rect 24811 29668 24860 29696
rect 24811 29665 24823 29668
rect 24765 29659 24823 29665
rect 24854 29656 24860 29668
rect 24912 29656 24918 29708
rect 27430 29696 27436 29708
rect 27080 29668 27436 29696
rect 27080 29640 27108 29668
rect 27430 29656 27436 29668
rect 27488 29696 27494 29708
rect 30469 29699 30527 29705
rect 30469 29696 30481 29699
rect 27488 29668 30481 29696
rect 27488 29656 27494 29668
rect 30469 29665 30481 29668
rect 30515 29696 30527 29699
rect 32858 29696 32864 29708
rect 30515 29668 32864 29696
rect 30515 29665 30527 29668
rect 30469 29659 30527 29665
rect 32858 29656 32864 29668
rect 32916 29656 32922 29708
rect 25590 29628 25596 29640
rect 24688 29600 25596 29628
rect 25590 29588 25596 29600
rect 25648 29628 25654 29640
rect 25777 29631 25835 29637
rect 25777 29628 25789 29631
rect 25648 29600 25789 29628
rect 25648 29588 25654 29600
rect 25777 29597 25789 29600
rect 25823 29597 25835 29631
rect 27062 29628 27068 29640
rect 27023 29600 27068 29628
rect 25777 29591 25835 29597
rect 27062 29588 27068 29600
rect 27120 29588 27126 29640
rect 29730 29628 29736 29640
rect 29691 29600 29736 29628
rect 29730 29588 29736 29600
rect 29788 29588 29794 29640
rect 30006 29588 30012 29640
rect 30064 29628 30070 29640
rect 33686 29628 33692 29640
rect 30064 29600 30109 29628
rect 33647 29600 33692 29628
rect 30064 29588 30070 29600
rect 33686 29588 33692 29600
rect 33744 29588 33750 29640
rect 48130 29628 48136 29640
rect 48091 29600 48136 29628
rect 48130 29588 48136 29600
rect 48188 29588 48194 29640
rect 20806 29560 20812 29572
rect 20456 29532 20812 29560
rect 20806 29520 20812 29532
rect 20864 29520 20870 29572
rect 27341 29563 27399 29569
rect 27341 29529 27353 29563
rect 27387 29560 27399 29563
rect 27430 29560 27436 29572
rect 27387 29532 27436 29560
rect 27387 29529 27399 29532
rect 27341 29523 27399 29529
rect 27430 29520 27436 29532
rect 27488 29520 27494 29572
rect 28350 29520 28356 29572
rect 28408 29520 28414 29572
rect 29549 29563 29607 29569
rect 29549 29529 29561 29563
rect 29595 29560 29607 29563
rect 30745 29563 30803 29569
rect 30745 29560 30757 29563
rect 29595 29532 30757 29560
rect 29595 29529 29607 29532
rect 29549 29523 29607 29529
rect 30745 29529 30757 29532
rect 30791 29529 30803 29563
rect 32122 29560 32128 29572
rect 31970 29532 32128 29560
rect 30745 29523 30803 29529
rect 32122 29520 32128 29532
rect 32180 29520 32186 29572
rect 20530 29452 20536 29504
rect 20588 29492 20594 29504
rect 20993 29495 21051 29501
rect 20993 29492 21005 29495
rect 20588 29464 21005 29492
rect 20588 29452 20594 29464
rect 20993 29461 21005 29464
rect 21039 29461 21051 29495
rect 20993 29455 21051 29461
rect 23106 29452 23112 29504
rect 23164 29492 23170 29504
rect 25961 29495 26019 29501
rect 25961 29492 25973 29495
rect 23164 29464 25973 29492
rect 23164 29452 23170 29464
rect 25961 29461 25973 29464
rect 26007 29492 26019 29495
rect 27982 29492 27988 29504
rect 26007 29464 27988 29492
rect 26007 29461 26019 29464
rect 25961 29455 26019 29461
rect 27982 29452 27988 29464
rect 28040 29452 28046 29504
rect 30006 29452 30012 29504
rect 30064 29492 30070 29504
rect 32217 29495 32275 29501
rect 32217 29492 32229 29495
rect 30064 29464 32229 29492
rect 30064 29452 30070 29464
rect 32217 29461 32229 29464
rect 32263 29461 32275 29495
rect 47946 29492 47952 29504
rect 47907 29464 47952 29492
rect 32217 29455 32275 29461
rect 47946 29452 47952 29464
rect 48004 29452 48010 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 19521 29291 19579 29297
rect 19521 29257 19533 29291
rect 19567 29288 19579 29291
rect 19978 29288 19984 29300
rect 19567 29260 19984 29288
rect 19567 29257 19579 29260
rect 19521 29251 19579 29257
rect 19978 29248 19984 29260
rect 20036 29248 20042 29300
rect 20898 29248 20904 29300
rect 20956 29288 20962 29300
rect 21726 29288 21732 29300
rect 20956 29260 21732 29288
rect 20956 29248 20962 29260
rect 21726 29248 21732 29260
rect 21784 29288 21790 29300
rect 25406 29288 25412 29300
rect 21784 29260 24992 29288
rect 25367 29260 25412 29288
rect 21784 29248 21790 29260
rect 16850 29220 16856 29232
rect 16684 29192 16856 29220
rect 16684 29164 16712 29192
rect 16850 29180 16856 29192
rect 16908 29180 16914 29232
rect 18969 29223 19027 29229
rect 18969 29220 18981 29223
rect 18170 29192 18981 29220
rect 18969 29189 18981 29192
rect 19015 29189 19027 29223
rect 21910 29220 21916 29232
rect 18969 29183 19027 29189
rect 19904 29192 20852 29220
rect 19904 29164 19932 29192
rect 16666 29152 16672 29164
rect 16579 29124 16672 29152
rect 16666 29112 16672 29124
rect 16724 29112 16730 29164
rect 18230 29112 18236 29164
rect 18288 29152 18294 29164
rect 18877 29155 18935 29161
rect 18877 29152 18889 29155
rect 18288 29124 18889 29152
rect 18288 29112 18294 29124
rect 18877 29121 18889 29124
rect 18923 29121 18935 29155
rect 19705 29155 19763 29161
rect 19705 29152 19717 29155
rect 18877 29115 18935 29121
rect 19628 29124 19717 29152
rect 18417 29087 18475 29093
rect 18417 29053 18429 29087
rect 18463 29084 18475 29087
rect 19628 29084 19656 29124
rect 19705 29121 19717 29124
rect 19751 29152 19763 29155
rect 19886 29152 19892 29164
rect 19751 29124 19892 29152
rect 19751 29121 19763 29124
rect 19705 29115 19763 29121
rect 19886 29112 19892 29124
rect 19944 29112 19950 29164
rect 19981 29155 20039 29161
rect 19981 29121 19993 29155
rect 20027 29152 20039 29155
rect 20070 29152 20076 29164
rect 20027 29124 20076 29152
rect 20027 29121 20039 29124
rect 19981 29115 20039 29121
rect 20070 29112 20076 29124
rect 20128 29112 20134 29164
rect 20530 29152 20536 29164
rect 20491 29124 20536 29152
rect 20530 29112 20536 29124
rect 20588 29112 20594 29164
rect 20824 29161 20852 29192
rect 21100 29192 21916 29220
rect 21100 29161 21128 29192
rect 21910 29180 21916 29192
rect 21968 29220 21974 29232
rect 23014 29220 23020 29232
rect 21968 29192 23020 29220
rect 21968 29180 21974 29192
rect 23014 29180 23020 29192
rect 23072 29180 23078 29232
rect 20717 29155 20775 29161
rect 20717 29121 20729 29155
rect 20763 29121 20775 29155
rect 20717 29115 20775 29121
rect 20809 29155 20867 29161
rect 20809 29121 20821 29155
rect 20855 29121 20867 29155
rect 20809 29115 20867 29121
rect 21085 29155 21143 29161
rect 21085 29121 21097 29155
rect 21131 29121 21143 29155
rect 21085 29115 21143 29121
rect 18463 29056 19656 29084
rect 18463 29053 18475 29056
rect 18417 29047 18475 29053
rect 19426 28976 19432 29028
rect 19484 29016 19490 29028
rect 19889 29019 19947 29025
rect 19889 29016 19901 29019
rect 19484 28988 19901 29016
rect 19484 28976 19490 28988
rect 19889 28985 19901 28988
rect 19935 28985 19947 29019
rect 20732 29016 20760 29115
rect 21818 29112 21824 29164
rect 21876 29152 21882 29164
rect 21876 29124 22048 29152
rect 21876 29112 21882 29124
rect 20901 29087 20959 29093
rect 20901 29053 20913 29087
rect 20947 29084 20959 29087
rect 21174 29084 21180 29096
rect 20947 29056 21180 29084
rect 20947 29053 20959 29056
rect 20901 29047 20959 29053
rect 21174 29044 21180 29056
rect 21232 29044 21238 29096
rect 22020 29084 22048 29124
rect 22094 29112 22100 29164
rect 22152 29152 22158 29164
rect 22649 29155 22707 29161
rect 22649 29152 22661 29155
rect 22152 29124 22661 29152
rect 22152 29112 22158 29124
rect 22649 29121 22661 29124
rect 22695 29121 22707 29155
rect 22649 29115 22707 29121
rect 24026 29112 24032 29164
rect 24084 29112 24090 29164
rect 24578 29112 24584 29164
rect 24636 29152 24642 29164
rect 24857 29155 24915 29161
rect 24857 29152 24869 29155
rect 24636 29124 24869 29152
rect 24636 29112 24642 29124
rect 24857 29121 24869 29124
rect 24903 29121 24915 29155
rect 24857 29115 24915 29121
rect 22112 29084 22140 29112
rect 22922 29084 22928 29096
rect 22020 29056 22140 29084
rect 22883 29056 22928 29084
rect 22922 29044 22928 29056
rect 22980 29044 22986 29096
rect 22646 29016 22652 29028
rect 20732 28988 22652 29016
rect 19889 28979 19947 28985
rect 22646 28976 22652 28988
rect 22704 28976 22710 29028
rect 24964 29016 24992 29260
rect 25406 29248 25412 29260
rect 25464 29248 25470 29300
rect 27430 29288 27436 29300
rect 27391 29260 27436 29288
rect 27430 29248 27436 29260
rect 27488 29248 27494 29300
rect 29730 29248 29736 29300
rect 29788 29288 29794 29300
rect 30193 29291 30251 29297
rect 30193 29288 30205 29291
rect 29788 29260 30205 29288
rect 29788 29248 29794 29260
rect 30193 29257 30205 29260
rect 30239 29257 30251 29291
rect 30193 29251 30251 29257
rect 32122 29248 32128 29300
rect 32180 29288 32186 29300
rect 32217 29291 32275 29297
rect 32217 29288 32229 29291
rect 32180 29260 32229 29288
rect 32180 29248 32186 29260
rect 32217 29257 32229 29260
rect 32263 29257 32275 29291
rect 32217 29251 32275 29257
rect 25424 29152 25452 29248
rect 28997 29223 29055 29229
rect 28997 29220 29009 29223
rect 27632 29192 29009 29220
rect 27632 29161 27660 29192
rect 28997 29189 29009 29192
rect 29043 29189 29055 29223
rect 43346 29220 43352 29232
rect 28997 29183 29055 29189
rect 30392 29192 43352 29220
rect 25869 29155 25927 29161
rect 25869 29152 25881 29155
rect 25424 29124 25881 29152
rect 25869 29121 25881 29124
rect 25915 29121 25927 29155
rect 25869 29115 25927 29121
rect 27617 29155 27675 29161
rect 27617 29121 27629 29155
rect 27663 29121 27675 29155
rect 27617 29115 27675 29121
rect 27706 29112 27712 29164
rect 27764 29152 27770 29164
rect 27982 29152 27988 29164
rect 27764 29124 27809 29152
rect 27943 29124 27988 29152
rect 27764 29112 27770 29124
rect 27982 29112 27988 29124
rect 28040 29112 28046 29164
rect 28810 29152 28816 29164
rect 28771 29124 28816 29152
rect 28810 29112 28816 29124
rect 28868 29152 28874 29164
rect 30282 29152 30288 29164
rect 28868 29124 30288 29152
rect 28868 29112 28874 29124
rect 30282 29112 30288 29124
rect 30340 29112 30346 29164
rect 30392 29161 30420 29192
rect 43346 29180 43352 29192
rect 43404 29180 43410 29232
rect 30377 29155 30435 29161
rect 30377 29121 30389 29155
rect 30423 29121 30435 29155
rect 30377 29115 30435 29121
rect 30469 29155 30527 29161
rect 30469 29121 30481 29155
rect 30515 29121 30527 29155
rect 30469 29115 30527 29121
rect 25130 29084 25136 29096
rect 25043 29056 25136 29084
rect 25130 29044 25136 29056
rect 25188 29084 25194 29096
rect 25682 29084 25688 29096
rect 25188 29056 25688 29084
rect 25188 29044 25194 29056
rect 25682 29044 25688 29056
rect 25740 29044 25746 29096
rect 28629 29087 28687 29093
rect 27816 29056 28580 29084
rect 27816 29028 27844 29056
rect 26053 29019 26111 29025
rect 26053 29016 26065 29019
rect 24964 28988 26065 29016
rect 26053 28985 26065 28988
rect 26099 29016 26111 29019
rect 27798 29016 27804 29028
rect 26099 28988 27804 29016
rect 26099 28985 26111 28988
rect 26053 28979 26111 28985
rect 27798 28976 27804 28988
rect 27856 28976 27862 29028
rect 27893 29019 27951 29025
rect 27893 28985 27905 29019
rect 27939 29016 27951 29019
rect 27982 29016 27988 29028
rect 27939 28988 27988 29016
rect 27939 28985 27951 28988
rect 27893 28979 27951 28985
rect 27982 28976 27988 28988
rect 28040 28976 28046 29028
rect 28552 29016 28580 29056
rect 28629 29053 28641 29087
rect 28675 29084 28687 29087
rect 28994 29084 29000 29096
rect 28675 29056 29000 29084
rect 28675 29053 28687 29056
rect 28629 29047 28687 29053
rect 28994 29044 29000 29056
rect 29052 29044 29058 29096
rect 30484 29084 30512 29115
rect 30558 29112 30564 29164
rect 30616 29152 30622 29164
rect 30653 29155 30711 29161
rect 30653 29152 30665 29155
rect 30616 29124 30665 29152
rect 30616 29112 30622 29124
rect 30653 29121 30665 29124
rect 30699 29121 30711 29155
rect 30653 29115 30711 29121
rect 30742 29112 30748 29164
rect 30800 29152 30806 29164
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 30800 29124 30845 29152
rect 31726 29124 32137 29152
rect 30800 29112 30806 29124
rect 30484 29056 30696 29084
rect 30668 29028 30696 29056
rect 29638 29016 29644 29028
rect 28552 28988 29644 29016
rect 29638 28976 29644 28988
rect 29696 29016 29702 29028
rect 30006 29016 30012 29028
rect 29696 28988 30012 29016
rect 29696 28976 29702 28988
rect 30006 28976 30012 28988
rect 30064 28976 30070 29028
rect 30650 28976 30656 29028
rect 30708 28976 30714 29028
rect 16932 28951 16990 28957
rect 16932 28917 16944 28951
rect 16978 28948 16990 28951
rect 21269 28951 21327 28957
rect 21269 28948 21281 28951
rect 16978 28920 21281 28948
rect 16978 28917 16990 28920
rect 16932 28911 16990 28917
rect 21269 28917 21281 28920
rect 21315 28917 21327 28951
rect 24394 28948 24400 28960
rect 24355 28920 24400 28948
rect 21269 28911 21327 28917
rect 24394 28908 24400 28920
rect 24452 28908 24458 28960
rect 25225 28951 25283 28957
rect 25225 28917 25237 28951
rect 25271 28948 25283 28951
rect 25498 28948 25504 28960
rect 25271 28920 25504 28948
rect 25271 28917 25283 28920
rect 25225 28911 25283 28917
rect 25498 28908 25504 28920
rect 25556 28908 25562 28960
rect 28258 28908 28264 28960
rect 28316 28948 28322 28960
rect 31726 28948 31754 29124
rect 32125 29121 32137 29124
rect 32171 29152 32183 29155
rect 33686 29152 33692 29164
rect 32171 29124 33692 29152
rect 32171 29121 32183 29124
rect 32125 29115 32183 29121
rect 33686 29112 33692 29124
rect 33744 29112 33750 29164
rect 28316 28920 31754 28948
rect 28316 28908 28322 28920
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 19981 28747 20039 28753
rect 19981 28713 19993 28747
rect 20027 28744 20039 28747
rect 20070 28744 20076 28756
rect 20027 28716 20076 28744
rect 20027 28713 20039 28716
rect 19981 28707 20039 28713
rect 20070 28704 20076 28716
rect 20128 28704 20134 28756
rect 22922 28704 22928 28756
rect 22980 28744 22986 28756
rect 23293 28747 23351 28753
rect 23293 28744 23305 28747
rect 22980 28716 23305 28744
rect 22980 28704 22986 28716
rect 23293 28713 23305 28716
rect 23339 28713 23351 28747
rect 23293 28707 23351 28713
rect 26970 28704 26976 28756
rect 27028 28744 27034 28756
rect 27065 28747 27123 28753
rect 27065 28744 27077 28747
rect 27028 28716 27077 28744
rect 27028 28704 27034 28716
rect 27065 28713 27077 28716
rect 27111 28744 27123 28747
rect 27154 28744 27160 28756
rect 27111 28716 27160 28744
rect 27111 28713 27123 28716
rect 27065 28707 27123 28713
rect 27154 28704 27160 28716
rect 27212 28704 27218 28756
rect 28350 28744 28356 28756
rect 28311 28716 28356 28744
rect 28350 28704 28356 28716
rect 28408 28704 28414 28756
rect 30101 28747 30159 28753
rect 30101 28713 30113 28747
rect 30147 28744 30159 28747
rect 30742 28744 30748 28756
rect 30147 28716 30748 28744
rect 30147 28713 30159 28716
rect 30101 28707 30159 28713
rect 30742 28704 30748 28716
rect 30800 28704 30806 28756
rect 20714 28636 20720 28688
rect 20772 28676 20778 28688
rect 25409 28679 25467 28685
rect 25409 28676 25421 28679
rect 20772 28648 25421 28676
rect 20772 28636 20778 28648
rect 25409 28645 25421 28648
rect 25455 28676 25467 28679
rect 30190 28676 30196 28688
rect 25455 28648 30196 28676
rect 25455 28645 25467 28648
rect 25409 28639 25467 28645
rect 30190 28636 30196 28648
rect 30248 28636 30254 28688
rect 7466 28568 7472 28620
rect 7524 28608 7530 28620
rect 19886 28608 19892 28620
rect 7524 28580 18644 28608
rect 19847 28580 19892 28608
rect 7524 28568 7530 28580
rect 17681 28543 17739 28549
rect 17681 28509 17693 28543
rect 17727 28540 17739 28543
rect 18138 28540 18144 28552
rect 17727 28512 18144 28540
rect 17727 28509 17739 28512
rect 17681 28503 17739 28509
rect 18138 28500 18144 28512
rect 18196 28500 18202 28552
rect 18322 28472 18328 28484
rect 18283 28444 18328 28472
rect 18322 28432 18328 28444
rect 18380 28432 18386 28484
rect 18506 28472 18512 28484
rect 18467 28444 18512 28472
rect 18506 28432 18512 28444
rect 18564 28432 18570 28484
rect 18616 28472 18644 28580
rect 19886 28568 19892 28580
rect 19944 28568 19950 28620
rect 21177 28611 21235 28617
rect 21177 28577 21189 28611
rect 21223 28608 21235 28611
rect 22278 28608 22284 28620
rect 21223 28580 22284 28608
rect 21223 28577 21235 28580
rect 21177 28571 21235 28577
rect 22278 28568 22284 28580
rect 22336 28568 22342 28620
rect 22833 28611 22891 28617
rect 22833 28577 22845 28611
rect 22879 28608 22891 28611
rect 23474 28608 23480 28620
rect 22879 28580 23480 28608
rect 22879 28577 22891 28580
rect 22833 28571 22891 28577
rect 23474 28568 23480 28580
rect 23532 28568 23538 28620
rect 25498 28568 25504 28620
rect 25556 28608 25562 28620
rect 28534 28608 28540 28620
rect 25556 28580 28540 28608
rect 25556 28568 25562 28580
rect 28534 28568 28540 28580
rect 28592 28568 28598 28620
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 19797 28543 19855 28549
rect 19797 28540 19809 28543
rect 19392 28512 19809 28540
rect 19392 28500 19398 28512
rect 19797 28509 19809 28512
rect 19843 28509 19855 28543
rect 19797 28503 19855 28509
rect 21082 28500 21088 28552
rect 21140 28540 21146 28552
rect 21453 28543 21511 28549
rect 21453 28540 21465 28543
rect 21140 28512 21465 28540
rect 21140 28500 21146 28512
rect 21453 28509 21465 28512
rect 21499 28509 21511 28543
rect 21453 28503 21511 28509
rect 22186 28500 22192 28552
rect 22244 28540 22250 28552
rect 22557 28543 22615 28549
rect 22557 28540 22569 28543
rect 22244 28512 22569 28540
rect 22244 28500 22250 28512
rect 22557 28509 22569 28512
rect 22603 28509 22615 28543
rect 22557 28503 22615 28509
rect 22646 28500 22652 28552
rect 22704 28540 22710 28552
rect 22741 28543 22799 28549
rect 22741 28540 22753 28543
rect 22704 28512 22753 28540
rect 22704 28500 22710 28512
rect 22741 28509 22753 28512
rect 22787 28509 22799 28543
rect 22741 28503 22799 28509
rect 22925 28543 22983 28549
rect 22925 28509 22937 28543
rect 22971 28509 22983 28543
rect 23106 28540 23112 28552
rect 23067 28512 23112 28540
rect 22925 28503 22983 28509
rect 22940 28472 22968 28503
rect 23106 28500 23112 28512
rect 23164 28500 23170 28552
rect 25225 28543 25283 28549
rect 25225 28509 25237 28543
rect 25271 28540 25283 28543
rect 25406 28540 25412 28552
rect 25271 28512 25412 28540
rect 25271 28509 25283 28512
rect 25225 28503 25283 28509
rect 25406 28500 25412 28512
rect 25464 28500 25470 28552
rect 26881 28543 26939 28549
rect 26881 28509 26893 28543
rect 26927 28509 26939 28543
rect 28258 28540 28264 28552
rect 28219 28512 28264 28540
rect 26881 28503 26939 28509
rect 18616 28444 22968 28472
rect 24486 28432 24492 28484
rect 24544 28472 24550 28484
rect 26896 28472 26924 28503
rect 28258 28500 28264 28512
rect 28316 28500 28322 28552
rect 30374 28540 30380 28552
rect 30335 28512 30380 28540
rect 30374 28500 30380 28512
rect 30432 28500 30438 28552
rect 24544 28444 26924 28472
rect 24544 28432 24550 28444
rect 17770 28404 17776 28416
rect 17731 28376 17776 28404
rect 17770 28364 17776 28376
rect 17828 28364 17834 28416
rect 18693 28407 18751 28413
rect 18693 28373 18705 28407
rect 18739 28404 18751 28407
rect 19426 28404 19432 28416
rect 18739 28376 19432 28404
rect 18739 28373 18751 28376
rect 18693 28367 18751 28373
rect 19426 28364 19432 28376
rect 19484 28404 19490 28416
rect 19978 28404 19984 28416
rect 19484 28376 19984 28404
rect 19484 28364 19490 28376
rect 19978 28364 19984 28376
rect 20036 28364 20042 28416
rect 20165 28407 20223 28413
rect 20165 28373 20177 28407
rect 20211 28404 20223 28407
rect 20714 28404 20720 28416
rect 20211 28376 20720 28404
rect 20211 28373 20223 28376
rect 20165 28367 20223 28373
rect 20714 28364 20720 28376
rect 20772 28364 20778 28416
rect 21450 28364 21456 28416
rect 21508 28404 21514 28416
rect 24578 28404 24584 28416
rect 21508 28376 24584 28404
rect 21508 28364 21514 28376
rect 24578 28364 24584 28376
rect 24636 28364 24642 28416
rect 26896 28404 26924 28444
rect 29454 28432 29460 28484
rect 29512 28472 29518 28484
rect 30101 28475 30159 28481
rect 30101 28472 30113 28475
rect 29512 28444 30113 28472
rect 29512 28432 29518 28444
rect 30101 28441 30113 28444
rect 30147 28441 30159 28475
rect 30282 28472 30288 28484
rect 30243 28444 30288 28472
rect 30101 28435 30159 28441
rect 30282 28432 30288 28444
rect 30340 28432 30346 28484
rect 29546 28404 29552 28416
rect 26896 28376 29552 28404
rect 29546 28364 29552 28376
rect 29604 28364 29610 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 18506 28160 18512 28212
rect 18564 28200 18570 28212
rect 18601 28203 18659 28209
rect 18601 28200 18613 28203
rect 18564 28172 18613 28200
rect 18564 28160 18570 28172
rect 18601 28169 18613 28172
rect 18647 28200 18659 28203
rect 19334 28200 19340 28212
rect 18647 28172 19340 28200
rect 18647 28169 18659 28172
rect 18601 28163 18659 28169
rect 19334 28160 19340 28172
rect 19392 28200 19398 28212
rect 22186 28200 22192 28212
rect 19392 28172 19748 28200
rect 22147 28172 22192 28200
rect 19392 28160 19398 28172
rect 17770 28092 17776 28144
rect 17828 28092 17834 28144
rect 19426 28092 19432 28144
rect 19484 28132 19490 28144
rect 19484 28104 19656 28132
rect 19484 28092 19490 28104
rect 16666 28024 16672 28076
rect 16724 28064 16730 28076
rect 16853 28067 16911 28073
rect 16853 28064 16865 28067
rect 16724 28036 16865 28064
rect 16724 28024 16730 28036
rect 16853 28033 16865 28036
rect 16899 28033 16911 28067
rect 19518 28064 19524 28076
rect 19479 28036 19524 28064
rect 16853 28027 16911 28033
rect 19518 28024 19524 28036
rect 19576 28024 19582 28076
rect 19628 28073 19656 28104
rect 19614 28067 19672 28073
rect 19614 28033 19626 28067
rect 19660 28033 19672 28067
rect 19720 28064 19748 28172
rect 22186 28160 22192 28172
rect 22244 28160 22250 28212
rect 25590 28160 25596 28212
rect 25648 28200 25654 28212
rect 25685 28203 25743 28209
rect 25685 28200 25697 28203
rect 25648 28172 25697 28200
rect 25648 28160 25654 28172
rect 25685 28169 25697 28172
rect 25731 28169 25743 28203
rect 25685 28163 25743 28169
rect 19797 28135 19855 28141
rect 19797 28101 19809 28135
rect 19843 28132 19855 28135
rect 20625 28135 20683 28141
rect 19843 28104 20576 28132
rect 19843 28101 19855 28104
rect 19797 28095 19855 28101
rect 19897 28067 19955 28073
rect 19720 28054 19840 28064
rect 19897 28054 19909 28067
rect 19720 28036 19909 28054
rect 19614 28027 19672 28033
rect 19812 28033 19909 28036
rect 19943 28033 19955 28067
rect 19812 28027 19955 28033
rect 20027 28067 20085 28073
rect 20027 28033 20039 28067
rect 20073 28064 20085 28067
rect 20548 28064 20576 28104
rect 20625 28101 20637 28135
rect 20671 28132 20683 28135
rect 20714 28132 20720 28144
rect 20671 28104 20720 28132
rect 20671 28101 20683 28104
rect 20625 28095 20683 28101
rect 20714 28092 20720 28104
rect 20772 28092 20778 28144
rect 20809 28135 20867 28141
rect 20809 28101 20821 28135
rect 20855 28132 20867 28135
rect 21082 28132 21088 28144
rect 20855 28104 21088 28132
rect 20855 28101 20867 28104
rect 20809 28095 20867 28101
rect 21082 28092 21088 28104
rect 21140 28132 21146 28144
rect 21266 28132 21272 28144
rect 21140 28104 21272 28132
rect 21140 28092 21146 28104
rect 21266 28092 21272 28104
rect 21324 28092 21330 28144
rect 22094 28132 22100 28144
rect 21652 28104 22100 28132
rect 21652 28064 21680 28104
rect 22094 28092 22100 28104
rect 22152 28092 22158 28144
rect 23474 28132 23480 28144
rect 22848 28104 23480 28132
rect 20073 28036 20484 28064
rect 20548 28036 21680 28064
rect 20073 28033 20085 28036
rect 20027 28027 20085 28033
rect 19812 28026 19932 28027
rect 17129 27999 17187 28005
rect 17129 27965 17141 27999
rect 17175 27996 17187 27999
rect 20456 27996 20484 28036
rect 21726 28024 21732 28076
rect 21784 28064 21790 28076
rect 22848 28073 22876 28104
rect 23474 28092 23480 28104
rect 23532 28132 23538 28144
rect 23753 28135 23811 28141
rect 23753 28132 23765 28135
rect 23532 28104 23765 28132
rect 23532 28092 23538 28104
rect 23753 28101 23765 28104
rect 23799 28132 23811 28135
rect 24394 28132 24400 28144
rect 23799 28104 24400 28132
rect 23799 28101 23811 28104
rect 23753 28095 23811 28101
rect 24394 28092 24400 28104
rect 24452 28092 24458 28144
rect 29365 28135 29423 28141
rect 29365 28101 29377 28135
rect 29411 28132 29423 28135
rect 29454 28132 29460 28144
rect 29411 28104 29460 28132
rect 29411 28101 29423 28104
rect 29365 28095 29423 28101
rect 29454 28092 29460 28104
rect 29512 28092 29518 28144
rect 29546 28092 29552 28144
rect 29604 28132 29610 28144
rect 30650 28132 30656 28144
rect 29604 28104 30656 28132
rect 29604 28092 29610 28104
rect 30650 28092 30656 28104
rect 30708 28092 30714 28144
rect 21821 28067 21879 28073
rect 21821 28064 21833 28067
rect 21784 28036 21833 28064
rect 21784 28024 21790 28036
rect 21821 28033 21833 28036
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 22833 28067 22891 28073
rect 22833 28033 22845 28067
rect 22879 28033 22891 28067
rect 22833 28027 22891 28033
rect 23569 28067 23627 28073
rect 23569 28033 23581 28067
rect 23615 28033 23627 28067
rect 24670 28064 24676 28076
rect 24631 28036 24676 28064
rect 23569 28027 23627 28033
rect 20990 27996 20996 28008
rect 17175 27968 20208 27996
rect 20456 27968 20996 27996
rect 17175 27965 17187 27968
rect 17129 27959 17187 27965
rect 20180 27937 20208 27968
rect 20990 27956 20996 27968
rect 21048 27956 21054 28008
rect 21913 27999 21971 28005
rect 21913 27965 21925 27999
rect 21959 27996 21971 27999
rect 22922 27996 22928 28008
rect 21959 27968 22928 27996
rect 21959 27965 21971 27968
rect 21913 27959 21971 27965
rect 22922 27956 22928 27968
rect 22980 27956 22986 28008
rect 23109 27999 23167 28005
rect 23109 27965 23121 27999
rect 23155 27996 23167 27999
rect 23584 27996 23612 28027
rect 24670 28024 24676 28036
rect 24728 28024 24734 28076
rect 25501 28067 25559 28073
rect 25501 28033 25513 28067
rect 25547 28064 25559 28067
rect 26326 28064 26332 28076
rect 25547 28036 26332 28064
rect 25547 28033 25559 28036
rect 25501 28027 25559 28033
rect 26326 28024 26332 28036
rect 26384 28024 26390 28076
rect 30006 28064 30012 28076
rect 29967 28036 30012 28064
rect 30006 28024 30012 28036
rect 30064 28024 30070 28076
rect 30190 28064 30196 28076
rect 30151 28036 30196 28064
rect 30190 28024 30196 28036
rect 30248 28024 30254 28076
rect 30285 28067 30343 28073
rect 30285 28033 30297 28067
rect 30331 28064 30343 28067
rect 31478 28064 31484 28076
rect 30331 28036 31484 28064
rect 30331 28033 30343 28036
rect 30285 28027 30343 28033
rect 31478 28024 31484 28036
rect 31536 28024 31542 28076
rect 46290 28064 46296 28076
rect 41386 28036 46296 28064
rect 24762 27996 24768 28008
rect 23155 27968 23612 27996
rect 24723 27968 24768 27996
rect 23155 27965 23167 27968
rect 23109 27959 23167 27965
rect 20165 27931 20223 27937
rect 20165 27897 20177 27931
rect 20211 27897 20223 27931
rect 21266 27928 21272 27940
rect 20165 27891 20223 27897
rect 20272 27900 21272 27928
rect 18322 27820 18328 27872
rect 18380 27860 18386 27872
rect 19242 27860 19248 27872
rect 18380 27832 19248 27860
rect 18380 27820 18386 27832
rect 19242 27820 19248 27832
rect 19300 27860 19306 27872
rect 20272 27860 20300 27900
rect 21266 27888 21272 27900
rect 21324 27888 21330 27940
rect 22186 27888 22192 27940
rect 22244 27928 22250 27940
rect 23124 27928 23152 27959
rect 24762 27956 24768 27968
rect 24820 27956 24826 28008
rect 24946 27928 24952 27940
rect 22244 27900 23152 27928
rect 24780 27900 24952 27928
rect 22244 27888 22250 27900
rect 19300 27832 20300 27860
rect 19300 27820 19306 27832
rect 20806 27820 20812 27872
rect 20864 27860 20870 27872
rect 20901 27863 20959 27869
rect 20901 27860 20913 27863
rect 20864 27832 20913 27860
rect 20864 27820 20870 27832
rect 20901 27829 20913 27832
rect 20947 27860 20959 27863
rect 21082 27860 21088 27872
rect 20947 27832 21088 27860
rect 20947 27829 20959 27832
rect 20901 27823 20959 27829
rect 21082 27820 21088 27832
rect 21140 27820 21146 27872
rect 22005 27863 22063 27869
rect 22005 27829 22017 27863
rect 22051 27860 22063 27863
rect 22649 27863 22707 27869
rect 22649 27860 22661 27863
rect 22051 27832 22661 27860
rect 22051 27829 22063 27832
rect 22005 27823 22063 27829
rect 22649 27829 22661 27832
rect 22695 27829 22707 27863
rect 23014 27860 23020 27872
rect 22975 27832 23020 27860
rect 22649 27823 22707 27829
rect 23014 27820 23020 27832
rect 23072 27820 23078 27872
rect 23934 27860 23940 27872
rect 23895 27832 23940 27860
rect 23934 27820 23940 27832
rect 23992 27820 23998 27872
rect 24780 27869 24808 27900
rect 24946 27888 24952 27900
rect 25004 27928 25010 27940
rect 25130 27928 25136 27940
rect 25004 27900 25136 27928
rect 25004 27888 25010 27900
rect 25130 27888 25136 27900
rect 25188 27888 25194 27940
rect 24765 27863 24823 27869
rect 24765 27829 24777 27863
rect 24811 27829 24823 27863
rect 24765 27823 24823 27829
rect 24854 27820 24860 27872
rect 24912 27860 24918 27872
rect 25041 27863 25099 27869
rect 25041 27860 25053 27863
rect 24912 27832 25053 27860
rect 24912 27820 24918 27832
rect 25041 27829 25053 27832
rect 25087 27829 25099 27863
rect 30006 27860 30012 27872
rect 29967 27832 30012 27860
rect 25041 27823 25099 27829
rect 30006 27820 30012 27832
rect 30064 27820 30070 27872
rect 38746 27820 38752 27872
rect 38804 27860 38810 27872
rect 41386 27860 41414 28036
rect 46290 28024 46296 28036
rect 46348 28064 46354 28076
rect 46845 28067 46903 28073
rect 46845 28064 46857 28067
rect 46348 28036 46857 28064
rect 46348 28024 46354 28036
rect 46845 28033 46857 28036
rect 46891 28033 46903 28067
rect 46845 28027 46903 28033
rect 46934 27860 46940 27872
rect 38804 27832 41414 27860
rect 46895 27832 46940 27860
rect 38804 27820 38810 27832
rect 46934 27820 46940 27832
rect 46992 27820 46998 27872
rect 47762 27860 47768 27872
rect 47723 27832 47768 27860
rect 47762 27820 47768 27832
rect 47820 27820 47826 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 3326 27616 3332 27668
rect 3384 27656 3390 27668
rect 15102 27656 15108 27668
rect 3384 27628 15108 27656
rect 3384 27616 3390 27628
rect 15102 27616 15108 27628
rect 15160 27616 15166 27668
rect 19518 27616 19524 27668
rect 19576 27656 19582 27668
rect 20346 27656 20352 27668
rect 19576 27628 20352 27656
rect 19576 27616 19582 27628
rect 20346 27616 20352 27628
rect 20404 27616 20410 27668
rect 20714 27616 20720 27668
rect 20772 27656 20778 27668
rect 20993 27659 21051 27665
rect 20993 27656 21005 27659
rect 20772 27628 21005 27656
rect 20772 27616 20778 27628
rect 20993 27625 21005 27628
rect 21039 27625 21051 27659
rect 21450 27656 21456 27668
rect 21411 27628 21456 27656
rect 20993 27619 21051 27625
rect 21450 27616 21456 27628
rect 21508 27616 21514 27668
rect 23753 27659 23811 27665
rect 23753 27625 23765 27659
rect 23799 27656 23811 27659
rect 24670 27656 24676 27668
rect 23799 27628 24676 27656
rect 23799 27625 23811 27628
rect 23753 27619 23811 27625
rect 24670 27616 24676 27628
rect 24728 27616 24734 27668
rect 24765 27659 24823 27665
rect 24765 27625 24777 27659
rect 24811 27656 24823 27659
rect 26510 27656 26516 27668
rect 24811 27628 26516 27656
rect 24811 27625 24823 27628
rect 24765 27619 24823 27625
rect 26510 27616 26516 27628
rect 26568 27616 26574 27668
rect 30374 27616 30380 27668
rect 30432 27656 30438 27668
rect 30929 27659 30987 27665
rect 30929 27656 30941 27659
rect 30432 27628 30941 27656
rect 30432 27616 30438 27628
rect 30929 27625 30941 27628
rect 30975 27656 30987 27659
rect 30975 27628 31754 27656
rect 30975 27625 30987 27628
rect 30929 27619 30987 27625
rect 2222 27548 2228 27600
rect 2280 27588 2286 27600
rect 2280 27560 24624 27588
rect 2280 27548 2286 27560
rect 15010 27480 15016 27532
rect 15068 27520 15074 27532
rect 16114 27520 16120 27532
rect 15068 27492 15700 27520
rect 16075 27492 16120 27520
rect 15068 27480 15074 27492
rect 12986 27412 12992 27464
rect 13044 27452 13050 27464
rect 14277 27455 14335 27461
rect 14277 27452 14289 27455
rect 13044 27424 14289 27452
rect 13044 27412 13050 27424
rect 14277 27421 14289 27424
rect 14323 27421 14335 27455
rect 15672 27452 15700 27492
rect 16114 27480 16120 27492
rect 16172 27480 16178 27532
rect 16850 27520 16856 27532
rect 16224 27492 16856 27520
rect 16224 27452 16252 27492
rect 16850 27480 16856 27492
rect 16908 27480 16914 27532
rect 17034 27520 17040 27532
rect 16995 27492 17040 27520
rect 17034 27480 17040 27492
rect 17092 27480 17098 27532
rect 20714 27480 20720 27532
rect 20772 27520 20778 27532
rect 21177 27523 21235 27529
rect 21177 27520 21189 27523
rect 20772 27492 21189 27520
rect 20772 27480 20778 27492
rect 21177 27489 21189 27492
rect 21223 27520 21235 27523
rect 21223 27492 23704 27520
rect 21223 27489 21235 27492
rect 21177 27483 21235 27489
rect 15672 27424 16252 27452
rect 16577 27455 16635 27461
rect 14277 27415 14335 27421
rect 16577 27421 16589 27455
rect 16623 27421 16635 27455
rect 19242 27452 19248 27464
rect 19203 27424 19248 27452
rect 16577 27415 16635 27421
rect 14458 27384 14464 27396
rect 14419 27356 14464 27384
rect 14458 27344 14464 27356
rect 14516 27344 14522 27396
rect 13262 27276 13268 27328
rect 13320 27316 13326 27328
rect 16592 27316 16620 27415
rect 19242 27412 19248 27424
rect 19300 27412 19306 27464
rect 19334 27412 19340 27464
rect 19392 27452 19398 27464
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 19392 27424 19441 27452
rect 19392 27412 19398 27424
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 20254 27452 20260 27464
rect 20215 27424 20260 27452
rect 19429 27415 19487 27421
rect 20254 27412 20260 27424
rect 20312 27412 20318 27464
rect 20349 27455 20407 27461
rect 20349 27421 20361 27455
rect 20395 27421 20407 27455
rect 20349 27415 20407 27421
rect 21269 27455 21327 27461
rect 21269 27421 21281 27455
rect 21315 27452 21327 27455
rect 22278 27452 22284 27464
rect 21315 27424 22284 27452
rect 21315 27421 21327 27424
rect 21269 27415 21327 27421
rect 16758 27384 16764 27396
rect 16719 27356 16764 27384
rect 16758 27344 16764 27356
rect 16816 27344 16822 27396
rect 16850 27344 16856 27396
rect 16908 27384 16914 27396
rect 20364 27384 20392 27415
rect 22278 27412 22284 27424
rect 22336 27412 22342 27464
rect 22756 27461 22784 27492
rect 22741 27455 22799 27461
rect 22741 27421 22753 27455
rect 22787 27421 22799 27455
rect 22741 27415 22799 27421
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27452 22983 27455
rect 23014 27452 23020 27464
rect 22971 27424 23020 27452
rect 22971 27421 22983 27424
rect 22925 27415 22983 27421
rect 20990 27384 20996 27396
rect 16908 27356 20392 27384
rect 20951 27356 20996 27384
rect 16908 27344 16914 27356
rect 20990 27344 20996 27356
rect 21048 27344 21054 27396
rect 21082 27344 21088 27396
rect 21140 27384 21146 27396
rect 22940 27384 22968 27415
rect 23014 27412 23020 27424
rect 23072 27452 23078 27464
rect 23569 27455 23627 27461
rect 23569 27452 23581 27455
rect 23072 27424 23581 27452
rect 23072 27412 23078 27424
rect 23569 27421 23581 27424
rect 23615 27421 23627 27455
rect 23569 27415 23627 27421
rect 21140 27356 22968 27384
rect 23385 27387 23443 27393
rect 21140 27344 21146 27356
rect 23385 27353 23397 27387
rect 23431 27384 23443 27387
rect 23676 27384 23704 27492
rect 23934 27384 23940 27396
rect 23431 27356 23940 27384
rect 23431 27353 23443 27356
rect 23385 27347 23443 27353
rect 23934 27344 23940 27356
rect 23992 27344 23998 27396
rect 24596 27384 24624 27560
rect 24688 27520 24716 27616
rect 25590 27588 25596 27600
rect 25240 27560 25596 27588
rect 24688 27492 25176 27520
rect 24946 27412 24952 27464
rect 25004 27452 25010 27464
rect 25148 27461 25176 27492
rect 25240 27461 25268 27560
rect 25590 27548 25596 27560
rect 25648 27548 25654 27600
rect 25774 27548 25780 27600
rect 25832 27588 25838 27600
rect 26237 27591 26295 27597
rect 26237 27588 26249 27591
rect 25832 27560 26249 27588
rect 25832 27548 25838 27560
rect 26237 27557 26249 27560
rect 26283 27557 26295 27591
rect 31110 27588 31116 27600
rect 31071 27560 31116 27588
rect 26237 27551 26295 27557
rect 31110 27548 31116 27560
rect 31168 27548 31174 27600
rect 31386 27548 31392 27600
rect 31444 27588 31450 27600
rect 31573 27591 31631 27597
rect 31573 27588 31585 27591
rect 31444 27560 31585 27588
rect 31444 27548 31450 27560
rect 31573 27557 31585 27560
rect 31619 27557 31631 27591
rect 31573 27551 31631 27557
rect 28445 27523 28503 27529
rect 25332 27492 27384 27520
rect 25041 27455 25099 27461
rect 25041 27452 25053 27455
rect 25004 27424 25053 27452
rect 25004 27412 25010 27424
rect 25041 27421 25053 27424
rect 25087 27421 25099 27455
rect 25041 27415 25099 27421
rect 25133 27455 25191 27461
rect 25133 27421 25145 27455
rect 25179 27421 25191 27455
rect 25133 27415 25191 27421
rect 25225 27455 25283 27461
rect 25225 27421 25237 27455
rect 25271 27421 25283 27455
rect 25225 27415 25283 27421
rect 25332 27384 25360 27492
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27452 25467 27455
rect 25590 27452 25596 27464
rect 25455 27424 25596 27452
rect 25455 27421 25467 27424
rect 25409 27415 25467 27421
rect 25590 27412 25596 27424
rect 25648 27412 25654 27464
rect 25961 27455 26019 27461
rect 25961 27421 25973 27455
rect 26007 27421 26019 27455
rect 25961 27415 26019 27421
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27452 26111 27455
rect 26326 27452 26332 27464
rect 26099 27424 26332 27452
rect 26099 27421 26111 27424
rect 26053 27415 26111 27421
rect 24596 27356 25360 27384
rect 25976 27384 26004 27415
rect 26326 27412 26332 27424
rect 26384 27412 26390 27464
rect 27356 27461 27384 27492
rect 28445 27489 28457 27523
rect 28491 27520 28503 27523
rect 28902 27520 28908 27532
rect 28491 27492 28908 27520
rect 28491 27489 28503 27492
rect 28445 27483 28503 27489
rect 28902 27480 28908 27492
rect 28960 27520 28966 27532
rect 30837 27523 30895 27529
rect 30837 27520 30849 27523
rect 28960 27492 29868 27520
rect 28960 27480 28966 27492
rect 27065 27455 27123 27461
rect 27065 27421 27077 27455
rect 27111 27421 27123 27455
rect 27065 27415 27123 27421
rect 27341 27455 27399 27461
rect 27341 27421 27353 27455
rect 27387 27421 27399 27455
rect 27341 27415 27399 27421
rect 26142 27384 26148 27396
rect 25976 27356 26148 27384
rect 26142 27344 26148 27356
rect 26200 27344 26206 27396
rect 27080 27384 27108 27415
rect 27890 27412 27896 27464
rect 27948 27452 27954 27464
rect 29840 27461 29868 27492
rect 30024 27492 30849 27520
rect 30024 27461 30052 27492
rect 30837 27489 30849 27492
rect 30883 27520 30895 27523
rect 31202 27520 31208 27532
rect 30883 27492 31208 27520
rect 30883 27489 30895 27492
rect 30837 27483 30895 27489
rect 31202 27480 31208 27492
rect 31260 27480 31266 27532
rect 31726 27520 31754 27628
rect 42426 27616 42432 27668
rect 42484 27656 42490 27668
rect 45554 27656 45560 27668
rect 42484 27628 45560 27656
rect 42484 27616 42490 27628
rect 45554 27616 45560 27628
rect 45612 27616 45618 27668
rect 47762 27588 47768 27600
rect 46308 27560 47768 27588
rect 46308 27529 46336 27560
rect 47762 27548 47768 27560
rect 47820 27548 47826 27600
rect 46293 27523 46351 27529
rect 31726 27492 32076 27520
rect 28169 27455 28227 27461
rect 28169 27452 28181 27455
rect 27948 27424 28181 27452
rect 27948 27412 27954 27424
rect 28169 27421 28181 27424
rect 28215 27421 28227 27455
rect 28169 27415 28227 27421
rect 29825 27455 29883 27461
rect 29825 27421 29837 27455
rect 29871 27421 29883 27455
rect 29825 27415 29883 27421
rect 30009 27455 30067 27461
rect 30009 27421 30021 27455
rect 30055 27421 30067 27455
rect 30190 27452 30196 27464
rect 30103 27424 30196 27452
rect 30009 27415 30067 27421
rect 27080 27356 27844 27384
rect 19334 27316 19340 27328
rect 13320 27288 16620 27316
rect 19295 27288 19340 27316
rect 13320 27276 13326 27288
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 20533 27319 20591 27325
rect 20533 27285 20545 27319
rect 20579 27316 20591 27319
rect 21358 27316 21364 27328
rect 20579 27288 21364 27316
rect 20579 27285 20591 27288
rect 20533 27279 20591 27285
rect 21358 27276 21364 27288
rect 21416 27276 21422 27328
rect 22833 27319 22891 27325
rect 22833 27285 22845 27319
rect 22879 27316 22891 27319
rect 22922 27316 22928 27328
rect 22879 27288 22928 27316
rect 22879 27285 22891 27288
rect 22833 27279 22891 27285
rect 22922 27276 22928 27288
rect 22980 27276 22986 27328
rect 24946 27276 24952 27328
rect 25004 27316 25010 27328
rect 25498 27316 25504 27328
rect 25004 27288 25504 27316
rect 25004 27276 25010 27288
rect 25498 27276 25504 27288
rect 25556 27316 25562 27328
rect 25958 27316 25964 27328
rect 25556 27288 25964 27316
rect 25556 27276 25562 27288
rect 25958 27276 25964 27288
rect 26016 27276 26022 27328
rect 26878 27316 26884 27328
rect 26839 27288 26884 27316
rect 26878 27276 26884 27288
rect 26936 27276 26942 27328
rect 26970 27276 26976 27328
rect 27028 27316 27034 27328
rect 27816 27325 27844 27356
rect 27249 27319 27307 27325
rect 27249 27316 27261 27319
rect 27028 27288 27261 27316
rect 27028 27276 27034 27288
rect 27249 27285 27261 27288
rect 27295 27285 27307 27319
rect 27249 27279 27307 27285
rect 27801 27319 27859 27325
rect 27801 27285 27813 27319
rect 27847 27285 27859 27319
rect 28258 27316 28264 27328
rect 28219 27288 28264 27316
rect 27801 27279 27859 27285
rect 28258 27276 28264 27288
rect 28316 27276 28322 27328
rect 29840 27316 29868 27415
rect 30190 27412 30196 27424
rect 30248 27452 30254 27464
rect 30929 27455 30987 27461
rect 30248 27424 30788 27452
rect 30248 27412 30254 27424
rect 30653 27387 30711 27393
rect 30653 27353 30665 27387
rect 30699 27353 30711 27387
rect 30760 27384 30788 27424
rect 30929 27421 30941 27455
rect 30975 27452 30987 27455
rect 31754 27452 31760 27464
rect 30975 27424 31760 27452
rect 30975 27421 30987 27424
rect 30929 27415 30987 27421
rect 31754 27412 31760 27424
rect 31812 27452 31818 27464
rect 31938 27452 31944 27464
rect 31812 27424 31857 27452
rect 31899 27424 31944 27452
rect 31812 27412 31818 27424
rect 31938 27412 31944 27424
rect 31996 27412 32002 27464
rect 32048 27461 32076 27492
rect 46293 27489 46305 27523
rect 46339 27489 46351 27523
rect 46293 27483 46351 27489
rect 46477 27523 46535 27529
rect 46477 27489 46489 27523
rect 46523 27520 46535 27523
rect 46934 27520 46940 27532
rect 46523 27492 46940 27520
rect 46523 27489 46535 27492
rect 46477 27483 46535 27489
rect 46934 27480 46940 27492
rect 46992 27480 46998 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 32033 27455 32091 27461
rect 32033 27421 32045 27455
rect 32079 27452 32091 27455
rect 32306 27452 32312 27464
rect 32079 27424 32312 27452
rect 32079 27421 32091 27424
rect 32033 27415 32091 27421
rect 32306 27412 32312 27424
rect 32364 27412 32370 27464
rect 31956 27384 31984 27412
rect 30760 27356 31984 27384
rect 30653 27347 30711 27353
rect 30668 27316 30696 27347
rect 31386 27316 31392 27328
rect 29840 27288 31392 27316
rect 31386 27276 31392 27288
rect 31444 27276 31450 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 10965 27115 11023 27121
rect 10965 27081 10977 27115
rect 11011 27081 11023 27115
rect 13262 27112 13268 27124
rect 13223 27084 13268 27112
rect 10965 27075 11023 27081
rect 10980 27044 11008 27075
rect 13262 27072 13268 27084
rect 13320 27072 13326 27124
rect 14369 27115 14427 27121
rect 14369 27081 14381 27115
rect 14415 27112 14427 27115
rect 14458 27112 14464 27124
rect 14415 27084 14464 27112
rect 14415 27081 14427 27084
rect 14369 27075 14427 27081
rect 14458 27072 14464 27084
rect 14516 27072 14522 27124
rect 15657 27115 15715 27121
rect 15657 27081 15669 27115
rect 15703 27112 15715 27115
rect 16758 27112 16764 27124
rect 15703 27084 16764 27112
rect 15703 27081 15715 27084
rect 15657 27075 15715 27081
rect 16758 27072 16764 27084
rect 16816 27072 16822 27124
rect 19426 27112 19432 27124
rect 19387 27084 19432 27112
rect 19426 27072 19432 27084
rect 19484 27072 19490 27124
rect 20254 27072 20260 27124
rect 20312 27112 20318 27124
rect 20312 27084 22876 27112
rect 20312 27072 20318 27084
rect 11793 27047 11851 27053
rect 11793 27044 11805 27047
rect 10980 27016 11805 27044
rect 11793 27013 11805 27016
rect 11839 27013 11851 27047
rect 11793 27007 11851 27013
rect 12434 27004 12440 27056
rect 12492 27004 12498 27056
rect 10597 26979 10655 26985
rect 10597 26945 10609 26979
rect 10643 26945 10655 26979
rect 10597 26939 10655 26945
rect 10612 26840 10640 26939
rect 10689 26911 10747 26917
rect 10689 26877 10701 26911
rect 10735 26908 10747 26911
rect 11238 26908 11244 26920
rect 10735 26880 11244 26908
rect 10735 26877 10747 26880
rect 10689 26871 10747 26877
rect 11238 26868 11244 26880
rect 11296 26868 11302 26920
rect 11514 26908 11520 26920
rect 11475 26880 11520 26908
rect 11514 26868 11520 26880
rect 11572 26868 11578 26920
rect 12342 26908 12348 26920
rect 11624 26880 12348 26908
rect 11624 26840 11652 26880
rect 12342 26868 12348 26880
rect 12400 26908 12406 26920
rect 13280 26908 13308 27072
rect 17402 27004 17408 27056
rect 17460 27044 17466 27056
rect 21450 27044 21456 27056
rect 17460 27016 21456 27044
rect 17460 27004 17466 27016
rect 21450 27004 21456 27016
rect 21508 27004 21514 27056
rect 22186 27004 22192 27056
rect 22244 27044 22250 27056
rect 22848 27044 22876 27084
rect 22922 27072 22928 27124
rect 22980 27112 22986 27124
rect 26970 27112 26976 27124
rect 22980 27084 24900 27112
rect 22980 27072 22986 27084
rect 24486 27044 24492 27056
rect 22244 27016 22289 27044
rect 22848 27016 24492 27044
rect 22244 27004 22250 27016
rect 24486 27004 24492 27016
rect 24544 27004 24550 27056
rect 14274 26976 14280 26988
rect 14235 26948 14280 26976
rect 14274 26936 14280 26948
rect 14332 26976 14338 26988
rect 14921 26979 14979 26985
rect 14921 26976 14933 26979
rect 14332 26948 14933 26976
rect 14332 26936 14338 26948
rect 14921 26945 14933 26948
rect 14967 26945 14979 26979
rect 14921 26939 14979 26945
rect 15565 26979 15623 26985
rect 15565 26945 15577 26979
rect 15611 26976 15623 26979
rect 17218 26976 17224 26988
rect 15611 26948 17224 26976
rect 15611 26945 15623 26948
rect 15565 26939 15623 26945
rect 17218 26936 17224 26948
rect 17276 26936 17282 26988
rect 19334 26976 19340 26988
rect 19295 26948 19340 26976
rect 19334 26936 19340 26948
rect 19392 26936 19398 26988
rect 19521 26979 19579 26985
rect 19521 26945 19533 26979
rect 19567 26976 19579 26979
rect 19978 26976 19984 26988
rect 19567 26948 19984 26976
rect 19567 26945 19579 26948
rect 19521 26939 19579 26945
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 20441 26979 20499 26985
rect 20441 26945 20453 26979
rect 20487 26945 20499 26979
rect 20441 26939 20499 26945
rect 20625 26979 20683 26985
rect 20625 26945 20637 26979
rect 20671 26976 20683 26979
rect 20714 26976 20720 26988
rect 20671 26948 20720 26976
rect 20671 26945 20683 26948
rect 20625 26939 20683 26945
rect 12400 26880 13308 26908
rect 12400 26868 12406 26880
rect 17954 26868 17960 26920
rect 18012 26908 18018 26920
rect 20456 26908 20484 26939
rect 20714 26936 20720 26948
rect 20772 26936 20778 26988
rect 20809 26979 20867 26985
rect 20809 26945 20821 26979
rect 20855 26976 20867 26979
rect 21266 26976 21272 26988
rect 20855 26948 21272 26976
rect 20855 26945 20867 26948
rect 20809 26939 20867 26945
rect 21266 26936 21272 26948
rect 21324 26936 21330 26988
rect 21358 26936 21364 26988
rect 21416 26976 21422 26988
rect 21821 26979 21879 26985
rect 21821 26976 21833 26979
rect 21416 26948 21833 26976
rect 21416 26936 21422 26948
rect 21821 26945 21833 26948
rect 21867 26945 21879 26979
rect 21821 26939 21879 26945
rect 21910 26936 21916 26988
rect 21968 26976 21974 26988
rect 22094 26976 22100 26988
rect 21968 26948 22013 26976
rect 22055 26948 22100 26976
rect 21968 26936 21974 26948
rect 22094 26936 22100 26948
rect 22152 26936 22158 26988
rect 22327 26979 22385 26985
rect 22327 26945 22339 26979
rect 22373 26976 22385 26979
rect 22554 26976 22560 26988
rect 22373 26948 22560 26976
rect 22373 26945 22385 26948
rect 22327 26939 22385 26945
rect 22554 26936 22560 26948
rect 22612 26936 22618 26988
rect 24673 26979 24731 26985
rect 24673 26945 24685 26979
rect 24719 26976 24731 26979
rect 24762 26976 24768 26988
rect 24719 26948 24768 26976
rect 24719 26945 24731 26948
rect 24673 26939 24731 26945
rect 24762 26936 24768 26948
rect 24820 26936 24826 26988
rect 24872 26976 24900 27084
rect 26252 27084 26976 27112
rect 25130 27044 25136 27056
rect 25188 27053 25194 27056
rect 25188 27047 25216 27053
rect 25068 27016 25136 27044
rect 25130 27004 25136 27016
rect 25204 27044 25216 27047
rect 25774 27044 25780 27056
rect 25204 27016 25780 27044
rect 25204 27013 25216 27016
rect 25188 27007 25216 27013
rect 25188 27004 25194 27007
rect 25774 27004 25780 27016
rect 25832 27004 25838 27056
rect 26252 27044 26280 27084
rect 26970 27072 26976 27084
rect 27028 27072 27034 27124
rect 27614 27072 27620 27124
rect 27672 27112 27678 27124
rect 27709 27115 27767 27121
rect 27709 27112 27721 27115
rect 27672 27084 27721 27112
rect 27672 27072 27678 27084
rect 27709 27081 27721 27084
rect 27755 27081 27767 27115
rect 27709 27075 27767 27081
rect 28629 27115 28687 27121
rect 28629 27081 28641 27115
rect 28675 27112 28687 27115
rect 30466 27112 30472 27124
rect 28675 27084 30472 27112
rect 28675 27081 28687 27084
rect 28629 27075 28687 27081
rect 30466 27072 30472 27084
rect 30524 27072 30530 27124
rect 30929 27115 30987 27121
rect 30929 27112 30941 27115
rect 30576 27084 30941 27112
rect 30576 27044 30604 27084
rect 30929 27081 30941 27084
rect 30975 27081 30987 27115
rect 31478 27112 31484 27124
rect 31439 27084 31484 27112
rect 30929 27075 30987 27081
rect 31478 27072 31484 27084
rect 31536 27072 31542 27124
rect 26160 27016 26280 27044
rect 29656 27016 30604 27044
rect 26160 26985 26188 27016
rect 25041 26979 25099 26985
rect 25041 26976 25053 26979
rect 24872 26948 25053 26976
rect 25041 26945 25053 26948
rect 25087 26945 25099 26979
rect 26126 26979 26188 26985
rect 25041 26939 25099 26945
rect 25975 26969 26033 26975
rect 25975 26935 25987 26969
rect 26021 26966 26033 26969
rect 26021 26938 26096 26966
rect 26126 26945 26138 26979
rect 26172 26948 26188 26979
rect 26222 26979 26280 26985
rect 26172 26945 26184 26948
rect 26126 26939 26184 26945
rect 26222 26945 26234 26979
rect 26268 26945 26280 26979
rect 26222 26939 26280 26945
rect 26329 26979 26387 26985
rect 26329 26945 26341 26979
rect 26375 26976 26387 26979
rect 26510 26976 26516 26988
rect 26375 26948 26516 26976
rect 26375 26945 26387 26948
rect 26329 26939 26387 26945
rect 26021 26935 26033 26938
rect 25975 26929 26033 26935
rect 24946 26908 24952 26920
rect 18012 26880 20484 26908
rect 24907 26880 24952 26908
rect 18012 26868 18018 26880
rect 24946 26868 24952 26880
rect 25004 26868 25010 26920
rect 25682 26908 25688 26920
rect 25332 26880 25688 26908
rect 10612 26812 11652 26840
rect 20533 26843 20591 26849
rect 20533 26809 20545 26843
rect 20579 26840 20591 26843
rect 20990 26840 20996 26852
rect 20579 26812 20996 26840
rect 20579 26809 20591 26812
rect 20533 26803 20591 26809
rect 20990 26800 20996 26812
rect 21048 26840 21054 26852
rect 25332 26849 25360 26880
rect 25682 26868 25688 26880
rect 25740 26868 25746 26920
rect 25317 26843 25375 26849
rect 21048 26812 25268 26840
rect 21048 26800 21054 26812
rect 15013 26775 15071 26781
rect 15013 26741 15025 26775
rect 15059 26772 15071 26775
rect 15194 26772 15200 26784
rect 15059 26744 15200 26772
rect 15059 26741 15071 26744
rect 15013 26735 15071 26741
rect 15194 26732 15200 26744
rect 15252 26732 15258 26784
rect 19978 26732 19984 26784
rect 20036 26772 20042 26784
rect 20165 26775 20223 26781
rect 20165 26772 20177 26775
rect 20036 26744 20177 26772
rect 20036 26732 20042 26744
rect 20165 26741 20177 26744
rect 20211 26741 20223 26775
rect 20165 26735 20223 26741
rect 20717 26775 20775 26781
rect 20717 26741 20729 26775
rect 20763 26772 20775 26775
rect 20806 26772 20812 26784
rect 20763 26744 20812 26772
rect 20763 26741 20775 26744
rect 20717 26735 20775 26741
rect 20806 26732 20812 26744
rect 20864 26732 20870 26784
rect 22094 26732 22100 26784
rect 22152 26772 22158 26784
rect 22465 26775 22523 26781
rect 22465 26772 22477 26775
rect 22152 26744 22477 26772
rect 22152 26732 22158 26744
rect 22465 26741 22477 26744
rect 22511 26741 22523 26775
rect 25240 26772 25268 26812
rect 25317 26809 25329 26843
rect 25363 26809 25375 26843
rect 26068 26840 26096 26938
rect 26252 26908 26280 26939
rect 26510 26936 26516 26948
rect 26568 26936 26574 26988
rect 27522 26976 27528 26988
rect 27435 26948 27528 26976
rect 27522 26936 27528 26948
rect 27580 26976 27586 26988
rect 28258 26976 28264 26988
rect 27580 26948 28264 26976
rect 27580 26936 27586 26948
rect 28258 26936 28264 26948
rect 28316 26976 28322 26988
rect 29656 26985 29684 27016
rect 30650 27004 30656 27056
rect 30708 27044 30714 27056
rect 30708 27016 30753 27044
rect 30708 27004 30714 27016
rect 31202 27004 31208 27056
rect 31260 27044 31266 27056
rect 31260 27016 31616 27044
rect 31260 27004 31266 27016
rect 31588 26988 31616 27016
rect 28445 26979 28503 26985
rect 28445 26976 28457 26979
rect 28316 26948 28457 26976
rect 28316 26936 28322 26948
rect 28445 26945 28457 26948
rect 28491 26945 28503 26979
rect 28445 26939 28503 26945
rect 29641 26979 29699 26985
rect 29641 26945 29653 26979
rect 29687 26945 29699 26979
rect 29641 26939 29699 26945
rect 29825 26979 29883 26985
rect 29825 26945 29837 26979
rect 29871 26945 29883 26979
rect 29825 26939 29883 26945
rect 29917 26979 29975 26985
rect 29917 26945 29929 26979
rect 29963 26945 29975 26979
rect 30374 26976 30380 26988
rect 30335 26948 30380 26976
rect 29917 26939 29975 26945
rect 28460 26908 28488 26939
rect 29730 26908 29736 26920
rect 26252 26880 26372 26908
rect 28460 26880 29736 26908
rect 26344 26852 26372 26880
rect 29730 26868 29736 26880
rect 29788 26868 29794 26920
rect 26234 26840 26240 26852
rect 26068 26812 26240 26840
rect 25317 26803 25375 26809
rect 26234 26800 26240 26812
rect 26292 26800 26298 26852
rect 26326 26800 26332 26852
rect 26384 26800 26390 26852
rect 29840 26840 29868 26939
rect 28966 26812 29868 26840
rect 29932 26840 29960 26939
rect 30374 26936 30380 26948
rect 30432 26936 30438 26988
rect 30558 26976 30564 26988
rect 30519 26948 30564 26976
rect 30558 26936 30564 26948
rect 30616 26936 30622 26988
rect 30745 26979 30803 26985
rect 30745 26945 30757 26979
rect 30791 26945 30803 26979
rect 31386 26976 31392 26988
rect 31347 26948 31392 26976
rect 30745 26939 30803 26945
rect 30466 26868 30472 26920
rect 30524 26908 30530 26920
rect 30760 26908 30788 26939
rect 31386 26936 31392 26948
rect 31444 26936 31450 26988
rect 31570 26976 31576 26988
rect 31531 26948 31576 26976
rect 31570 26936 31576 26948
rect 31628 26936 31634 26988
rect 32306 26976 32312 26988
rect 32267 26948 32312 26976
rect 32306 26936 32312 26948
rect 32364 26936 32370 26988
rect 30524 26880 30788 26908
rect 30524 26868 30530 26880
rect 31938 26868 31944 26920
rect 31996 26908 32002 26920
rect 32217 26911 32275 26917
rect 32217 26908 32229 26911
rect 31996 26880 32229 26908
rect 31996 26868 32002 26880
rect 32217 26877 32229 26880
rect 32263 26877 32275 26911
rect 32217 26871 32275 26877
rect 46566 26868 46572 26920
rect 46624 26908 46630 26920
rect 46750 26908 46756 26920
rect 46624 26880 46756 26908
rect 46624 26868 46630 26880
rect 46750 26868 46756 26880
rect 46808 26868 46814 26920
rect 32677 26843 32735 26849
rect 32677 26840 32689 26843
rect 29932 26812 32689 26840
rect 25682 26772 25688 26784
rect 25240 26744 25688 26772
rect 22465 26735 22523 26741
rect 25682 26732 25688 26744
rect 25740 26732 25746 26784
rect 25774 26732 25780 26784
rect 25832 26772 25838 26784
rect 25832 26744 25877 26772
rect 25832 26732 25838 26744
rect 25958 26732 25964 26784
rect 26016 26772 26022 26784
rect 28966 26772 28994 26812
rect 32677 26809 32689 26812
rect 32723 26809 32735 26843
rect 32677 26803 32735 26809
rect 26016 26744 28994 26772
rect 29457 26775 29515 26781
rect 26016 26732 26022 26744
rect 29457 26741 29469 26775
rect 29503 26772 29515 26775
rect 31294 26772 31300 26784
rect 29503 26744 31300 26772
rect 29503 26741 29515 26744
rect 29457 26735 29515 26741
rect 31294 26732 31300 26744
rect 31352 26732 31358 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 11238 26568 11244 26580
rect 11199 26540 11244 26568
rect 11238 26528 11244 26540
rect 11296 26528 11302 26580
rect 20346 26568 20352 26580
rect 20307 26540 20352 26568
rect 20346 26528 20352 26540
rect 20404 26528 20410 26580
rect 21361 26571 21419 26577
rect 21361 26537 21373 26571
rect 21407 26568 21419 26571
rect 21910 26568 21916 26580
rect 21407 26540 21916 26568
rect 21407 26537 21419 26540
rect 21361 26531 21419 26537
rect 21910 26528 21916 26540
rect 21968 26528 21974 26580
rect 25130 26568 25136 26580
rect 24596 26540 25136 26568
rect 15102 26460 15108 26512
rect 15160 26500 15166 26512
rect 15160 26472 15516 26500
rect 15160 26460 15166 26472
rect 12618 26432 12624 26444
rect 11164 26404 12624 26432
rect 11164 26373 11192 26404
rect 12618 26392 12624 26404
rect 12676 26392 12682 26444
rect 15194 26432 15200 26444
rect 15155 26404 15200 26432
rect 15194 26392 15200 26404
rect 15252 26392 15258 26444
rect 15488 26441 15516 26472
rect 21082 26460 21088 26512
rect 21140 26460 21146 26512
rect 15473 26435 15531 26441
rect 15473 26401 15485 26435
rect 15519 26401 15531 26435
rect 15473 26395 15531 26401
rect 19981 26435 20039 26441
rect 19981 26401 19993 26435
rect 20027 26432 20039 26435
rect 20254 26432 20260 26444
rect 20027 26404 20260 26432
rect 20027 26401 20039 26404
rect 19981 26395 20039 26401
rect 20254 26392 20260 26404
rect 20312 26392 20318 26444
rect 21100 26432 21128 26460
rect 21177 26435 21235 26441
rect 21177 26432 21189 26435
rect 21100 26404 21189 26432
rect 21177 26401 21189 26404
rect 21223 26401 21235 26435
rect 21177 26395 21235 26401
rect 11149 26367 11207 26373
rect 11149 26333 11161 26367
rect 11195 26333 11207 26367
rect 11149 26327 11207 26333
rect 11333 26367 11391 26373
rect 11333 26333 11345 26367
rect 11379 26364 11391 26367
rect 12710 26364 12716 26376
rect 11379 26336 12716 26364
rect 11379 26333 11391 26336
rect 11333 26327 11391 26333
rect 12710 26324 12716 26336
rect 12768 26364 12774 26376
rect 12986 26364 12992 26376
rect 12768 26336 12992 26364
rect 12768 26324 12774 26336
rect 12986 26324 12992 26336
rect 13044 26324 13050 26376
rect 13265 26367 13323 26373
rect 13265 26333 13277 26367
rect 13311 26364 13323 26367
rect 14734 26364 14740 26376
rect 13311 26336 14740 26364
rect 13311 26333 13323 26336
rect 13265 26327 13323 26333
rect 14734 26324 14740 26336
rect 14792 26324 14798 26376
rect 15013 26367 15071 26373
rect 15013 26333 15025 26367
rect 15059 26333 15071 26367
rect 15013 26327 15071 26333
rect 20165 26367 20223 26373
rect 20165 26333 20177 26367
rect 20211 26364 20223 26367
rect 20346 26364 20352 26376
rect 20211 26336 20352 26364
rect 20211 26333 20223 26336
rect 20165 26327 20223 26333
rect 12526 26256 12532 26308
rect 12584 26296 12590 26308
rect 13357 26299 13415 26305
rect 13357 26296 13369 26299
rect 12584 26268 13369 26296
rect 12584 26256 12590 26268
rect 13357 26265 13369 26268
rect 13403 26265 13415 26299
rect 15028 26296 15056 26327
rect 20346 26324 20352 26336
rect 20404 26324 20410 26376
rect 21085 26367 21143 26373
rect 21085 26333 21097 26367
rect 21131 26364 21143 26367
rect 22186 26364 22192 26376
rect 21131 26336 22192 26364
rect 21131 26333 21143 26336
rect 21085 26327 21143 26333
rect 22186 26324 22192 26336
rect 22244 26324 22250 26376
rect 24596 26364 24624 26540
rect 25130 26528 25136 26540
rect 25188 26528 25194 26580
rect 26878 26528 26884 26580
rect 26936 26568 26942 26580
rect 27414 26571 27472 26577
rect 27414 26568 27426 26571
rect 26936 26540 27426 26568
rect 26936 26528 26942 26540
rect 27414 26537 27426 26540
rect 27460 26537 27472 26571
rect 28902 26568 28908 26580
rect 28863 26540 28908 26568
rect 27414 26531 27472 26537
rect 28902 26528 28908 26540
rect 28960 26528 28966 26580
rect 32306 26528 32312 26580
rect 32364 26568 32370 26580
rect 32769 26571 32827 26577
rect 32769 26568 32781 26571
rect 32364 26540 32781 26568
rect 32364 26528 32370 26540
rect 32769 26537 32781 26540
rect 32815 26537 32827 26571
rect 32769 26531 32827 26537
rect 24670 26460 24676 26512
rect 24728 26500 24734 26512
rect 25225 26503 25283 26509
rect 25225 26500 25237 26503
rect 24728 26472 25237 26500
rect 24728 26460 24734 26472
rect 25225 26469 25237 26472
rect 25271 26469 25283 26503
rect 25225 26463 25283 26469
rect 25682 26460 25688 26512
rect 25740 26500 25746 26512
rect 26053 26503 26111 26509
rect 26053 26500 26065 26503
rect 25740 26472 26065 26500
rect 25740 26460 25746 26472
rect 26053 26469 26065 26472
rect 26099 26469 26111 26503
rect 26053 26463 26111 26469
rect 29454 26460 29460 26512
rect 29512 26500 29518 26512
rect 29512 26472 29868 26500
rect 29512 26460 29518 26472
rect 24946 26392 24952 26444
rect 25004 26432 25010 26444
rect 25004 26404 25084 26432
rect 25004 26392 25010 26404
rect 24673 26367 24731 26373
rect 24673 26364 24685 26367
rect 24596 26336 24685 26364
rect 24673 26333 24685 26336
rect 24719 26333 24731 26367
rect 24854 26364 24860 26376
rect 24815 26336 24860 26364
rect 24673 26327 24731 26333
rect 24854 26324 24860 26336
rect 24912 26324 24918 26376
rect 25056 26373 25084 26404
rect 25041 26367 25099 26373
rect 25041 26333 25053 26367
rect 25087 26333 25099 26367
rect 26970 26364 26976 26376
rect 25041 26327 25099 26333
rect 25516 26336 26976 26364
rect 16482 26296 16488 26308
rect 15028 26268 16488 26296
rect 13357 26259 13415 26265
rect 16482 26256 16488 26268
rect 16540 26256 16546 26308
rect 24762 26256 24768 26308
rect 24820 26296 24826 26308
rect 24949 26299 25007 26305
rect 24820 26268 24900 26296
rect 24820 26256 24826 26268
rect 24872 26228 24900 26268
rect 24949 26265 24961 26299
rect 24995 26296 25007 26299
rect 25516 26296 25544 26336
rect 26970 26324 26976 26336
rect 27028 26324 27034 26376
rect 27154 26364 27160 26376
rect 27115 26336 27160 26364
rect 27154 26324 27160 26336
rect 27212 26324 27218 26376
rect 29549 26367 29607 26373
rect 29549 26333 29561 26367
rect 29595 26333 29607 26367
rect 29730 26364 29736 26376
rect 29691 26336 29736 26364
rect 29549 26327 29607 26333
rect 25682 26296 25688 26308
rect 24995 26268 25544 26296
rect 25643 26268 25688 26296
rect 24995 26265 25007 26268
rect 24949 26259 25007 26265
rect 25682 26256 25688 26268
rect 25740 26256 25746 26308
rect 25869 26299 25927 26305
rect 25869 26265 25881 26299
rect 25915 26296 25927 26299
rect 26142 26296 26148 26308
rect 25915 26268 26148 26296
rect 25915 26265 25927 26268
rect 25869 26259 25927 26265
rect 26142 26256 26148 26268
rect 26200 26256 26206 26308
rect 29086 26296 29092 26308
rect 28658 26268 29092 26296
rect 29086 26256 29092 26268
rect 29144 26256 29150 26308
rect 29564 26296 29592 26327
rect 29730 26324 29736 26336
rect 29788 26324 29794 26376
rect 29840 26373 29868 26472
rect 29914 26460 29920 26512
rect 29972 26460 29978 26512
rect 29932 26373 29960 26460
rect 30374 26392 30380 26444
rect 30432 26432 30438 26444
rect 31021 26435 31079 26441
rect 31021 26432 31033 26435
rect 30432 26404 31033 26432
rect 30432 26392 30438 26404
rect 31021 26401 31033 26404
rect 31067 26401 31079 26435
rect 31294 26432 31300 26444
rect 31255 26404 31300 26432
rect 31021 26395 31079 26401
rect 31294 26392 31300 26404
rect 31352 26392 31358 26444
rect 29825 26367 29883 26373
rect 29825 26333 29837 26367
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 29917 26367 29975 26373
rect 29917 26333 29929 26367
rect 29963 26333 29975 26367
rect 29917 26327 29975 26333
rect 45186 26324 45192 26376
rect 45244 26364 45250 26376
rect 47673 26367 47731 26373
rect 47673 26364 47685 26367
rect 45244 26336 47685 26364
rect 45244 26324 45250 26336
rect 47673 26333 47685 26336
rect 47719 26333 47731 26367
rect 47673 26327 47731 26333
rect 31570 26296 31576 26308
rect 29564 26268 31576 26296
rect 31570 26256 31576 26268
rect 31628 26256 31634 26308
rect 31754 26256 31760 26308
rect 31812 26256 31818 26308
rect 25700 26228 25728 26256
rect 30098 26228 30104 26240
rect 24872 26200 25728 26228
rect 30059 26200 30104 26228
rect 30098 26188 30104 26200
rect 30156 26188 30162 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 10781 26027 10839 26033
rect 10781 25993 10793 26027
rect 10827 26024 10839 26027
rect 11514 26024 11520 26036
rect 10827 25996 11520 26024
rect 10827 25993 10839 25996
rect 10781 25987 10839 25993
rect 11514 25984 11520 25996
rect 11572 25984 11578 26036
rect 12069 26027 12127 26033
rect 12069 25993 12081 26027
rect 12115 26024 12127 26027
rect 12434 26024 12440 26036
rect 12115 25996 12440 26024
rect 12115 25993 12127 25996
rect 12069 25987 12127 25993
rect 12434 25984 12440 25996
rect 12492 25984 12498 26036
rect 16850 25984 16856 26036
rect 16908 25984 16914 26036
rect 22186 25984 22192 26036
rect 22244 26024 22250 26036
rect 23569 26027 23627 26033
rect 23569 26024 23581 26027
rect 22244 25996 23581 26024
rect 22244 25984 22250 25996
rect 23569 25993 23581 25996
rect 23615 25993 23627 26027
rect 23569 25987 23627 25993
rect 24026 25984 24032 26036
rect 24084 26024 24090 26036
rect 24121 26027 24179 26033
rect 24121 26024 24133 26027
rect 24084 25996 24133 26024
rect 24084 25984 24090 25996
rect 24121 25993 24133 25996
rect 24167 25993 24179 26027
rect 27522 26024 27528 26036
rect 27483 25996 27528 26024
rect 24121 25987 24179 25993
rect 27522 25984 27528 25996
rect 27580 25984 27586 26036
rect 29086 26024 29092 26036
rect 29047 25996 29092 26024
rect 29086 25984 29092 25996
rect 29144 25984 29150 26036
rect 31481 26027 31539 26033
rect 31481 25993 31493 26027
rect 31527 26024 31539 26027
rect 31754 26024 31760 26036
rect 31527 25996 31760 26024
rect 31527 25993 31539 25996
rect 31481 25987 31539 25993
rect 31754 25984 31760 25996
rect 31812 25984 31818 26036
rect 16868 25956 16896 25984
rect 12452 25928 15056 25956
rect 12452 25900 12480 25928
rect 10686 25888 10692 25900
rect 10647 25860 10692 25888
rect 10686 25848 10692 25860
rect 10744 25848 10750 25900
rect 11977 25891 12035 25897
rect 11977 25857 11989 25891
rect 12023 25888 12035 25891
rect 12434 25888 12440 25900
rect 12023 25860 12440 25888
rect 12023 25857 12035 25860
rect 11977 25851 12035 25857
rect 12434 25848 12440 25860
rect 12492 25848 12498 25900
rect 12805 25891 12863 25897
rect 12805 25857 12817 25891
rect 12851 25888 12863 25891
rect 13817 25891 13875 25897
rect 12851 25860 13492 25888
rect 12851 25857 12863 25860
rect 12805 25851 12863 25857
rect 13464 25832 13492 25860
rect 13817 25857 13829 25891
rect 13863 25888 13875 25891
rect 13998 25888 14004 25900
rect 13863 25860 14004 25888
rect 13863 25857 13875 25860
rect 13817 25851 13875 25857
rect 13998 25848 14004 25860
rect 14056 25848 14062 25900
rect 15028 25897 15056 25928
rect 16684 25928 18184 25956
rect 16684 25897 16712 25928
rect 15013 25891 15071 25897
rect 15013 25857 15025 25891
rect 15059 25857 15071 25891
rect 15013 25851 15071 25857
rect 16669 25891 16727 25897
rect 16669 25857 16681 25891
rect 16715 25857 16727 25891
rect 16669 25851 16727 25857
rect 16758 25848 16764 25900
rect 16816 25888 16822 25900
rect 16853 25891 16911 25897
rect 16853 25888 16865 25891
rect 16816 25860 16865 25888
rect 16816 25848 16822 25860
rect 16853 25857 16865 25860
rect 16899 25857 16911 25891
rect 17681 25891 17739 25897
rect 17681 25888 17693 25891
rect 16853 25851 16911 25857
rect 16960 25860 17693 25888
rect 13081 25823 13139 25829
rect 13081 25789 13093 25823
rect 13127 25820 13139 25823
rect 13170 25820 13176 25832
rect 13127 25792 13176 25820
rect 13127 25789 13139 25792
rect 13081 25783 13139 25789
rect 13170 25780 13176 25792
rect 13228 25780 13234 25832
rect 13446 25780 13452 25832
rect 13504 25820 13510 25832
rect 13725 25823 13783 25829
rect 13725 25820 13737 25823
rect 13504 25792 13737 25820
rect 13504 25780 13510 25792
rect 13725 25789 13737 25792
rect 13771 25789 13783 25823
rect 13725 25783 13783 25789
rect 11790 25712 11796 25764
rect 11848 25752 11854 25764
rect 12989 25755 13047 25761
rect 12989 25752 13001 25755
rect 11848 25724 13001 25752
rect 11848 25712 11854 25724
rect 12989 25721 13001 25724
rect 13035 25721 13047 25755
rect 12989 25715 13047 25721
rect 14734 25712 14740 25764
rect 14792 25752 14798 25764
rect 16960 25752 16988 25860
rect 17681 25857 17693 25860
rect 17727 25857 17739 25891
rect 17681 25851 17739 25857
rect 18156 25832 18184 25928
rect 22094 25916 22100 25968
rect 22152 25956 22158 25968
rect 22152 25928 22197 25956
rect 22152 25916 22158 25928
rect 22830 25916 22836 25968
rect 22888 25916 22894 25968
rect 28537 25959 28595 25965
rect 28537 25956 28549 25959
rect 27632 25928 28549 25956
rect 18230 25848 18236 25900
rect 18288 25888 18294 25900
rect 18417 25891 18475 25897
rect 18417 25888 18429 25891
rect 18288 25860 18429 25888
rect 18288 25848 18294 25860
rect 18417 25857 18429 25860
rect 18463 25857 18475 25891
rect 18417 25851 18475 25857
rect 18601 25891 18659 25897
rect 18601 25857 18613 25891
rect 18647 25888 18659 25891
rect 19978 25888 19984 25900
rect 18647 25860 19984 25888
rect 18647 25857 18659 25860
rect 18601 25851 18659 25857
rect 19978 25848 19984 25860
rect 20036 25848 20042 25900
rect 21818 25888 21824 25900
rect 21779 25860 21824 25888
rect 21818 25848 21824 25860
rect 21876 25848 21882 25900
rect 23382 25848 23388 25900
rect 23440 25888 23446 25900
rect 24029 25891 24087 25897
rect 24029 25888 24041 25891
rect 23440 25860 24041 25888
rect 23440 25848 23446 25860
rect 24029 25857 24041 25860
rect 24075 25888 24087 25891
rect 24765 25891 24823 25897
rect 24765 25888 24777 25891
rect 24075 25860 24777 25888
rect 24075 25857 24087 25860
rect 24029 25851 24087 25857
rect 24765 25857 24777 25860
rect 24811 25888 24823 25891
rect 25409 25891 25467 25897
rect 25409 25888 25421 25891
rect 24811 25860 25421 25888
rect 24811 25857 24823 25860
rect 24765 25851 24823 25857
rect 25409 25857 25421 25860
rect 25455 25857 25467 25891
rect 25409 25851 25467 25857
rect 25498 25848 25504 25900
rect 25556 25888 25562 25900
rect 27632 25897 27660 25928
rect 28537 25925 28549 25928
rect 28583 25956 28595 25959
rect 29454 25956 29460 25968
rect 28583 25928 29460 25956
rect 28583 25925 28595 25928
rect 28537 25919 28595 25925
rect 29454 25916 29460 25928
rect 29512 25916 29518 25968
rect 30006 25956 30012 25968
rect 29967 25928 30012 25956
rect 30006 25916 30012 25928
rect 30064 25916 30070 25968
rect 27249 25891 27307 25897
rect 27249 25888 27261 25891
rect 25556 25860 27261 25888
rect 25556 25848 25562 25860
rect 27249 25857 27261 25860
rect 27295 25857 27307 25891
rect 27249 25851 27307 25857
rect 27617 25891 27675 25897
rect 27617 25857 27629 25891
rect 27663 25857 27675 25891
rect 27617 25851 27675 25857
rect 28353 25891 28411 25897
rect 28353 25857 28365 25891
rect 28399 25857 28411 25891
rect 28353 25851 28411 25857
rect 28997 25891 29055 25897
rect 28997 25857 29009 25891
rect 29043 25857 29055 25891
rect 28997 25851 29055 25857
rect 29825 25891 29883 25897
rect 29825 25857 29837 25891
rect 29871 25888 29883 25891
rect 30098 25888 30104 25900
rect 29871 25860 30104 25888
rect 29871 25857 29883 25860
rect 29825 25851 29883 25857
rect 18138 25820 18144 25832
rect 18051 25792 18144 25820
rect 18138 25780 18144 25792
rect 18196 25820 18202 25832
rect 27065 25823 27123 25829
rect 27065 25820 27077 25823
rect 18196 25792 27077 25820
rect 18196 25780 18202 25792
rect 27065 25789 27077 25792
rect 27111 25789 27123 25823
rect 28368 25820 28396 25851
rect 28534 25820 28540 25832
rect 28368 25792 28540 25820
rect 27065 25783 27123 25789
rect 28534 25780 28540 25792
rect 28592 25780 28598 25832
rect 29012 25820 29040 25851
rect 30098 25848 30104 25860
rect 30156 25848 30162 25900
rect 30193 25891 30251 25897
rect 30193 25857 30205 25891
rect 30239 25888 30251 25891
rect 30837 25891 30895 25897
rect 30837 25888 30849 25891
rect 30239 25860 30849 25888
rect 30239 25857 30251 25860
rect 30193 25851 30251 25857
rect 30837 25857 30849 25860
rect 30883 25857 30895 25891
rect 30837 25851 30895 25857
rect 31389 25891 31447 25897
rect 31389 25857 31401 25891
rect 31435 25857 31447 25891
rect 46290 25888 46296 25900
rect 46251 25860 46296 25888
rect 31389 25851 31447 25857
rect 30282 25820 30288 25832
rect 29012 25792 30288 25820
rect 30282 25780 30288 25792
rect 30340 25820 30346 25832
rect 31404 25820 31432 25851
rect 46290 25848 46296 25860
rect 46348 25848 46354 25900
rect 30340 25792 31432 25820
rect 30340 25780 30346 25792
rect 14792 25724 16988 25752
rect 14792 25712 14798 25724
rect 12621 25687 12679 25693
rect 12621 25653 12633 25687
rect 12667 25684 12679 25687
rect 12802 25684 12808 25696
rect 12667 25656 12808 25684
rect 12667 25653 12679 25656
rect 12621 25647 12679 25653
rect 12802 25644 12808 25656
rect 12860 25644 12866 25696
rect 14093 25687 14151 25693
rect 14093 25653 14105 25687
rect 14139 25684 14151 25687
rect 14458 25684 14464 25696
rect 14139 25656 14464 25684
rect 14139 25653 14151 25656
rect 14093 25647 14151 25653
rect 14458 25644 14464 25656
rect 14516 25644 14522 25696
rect 15102 25684 15108 25696
rect 15063 25656 15108 25684
rect 15102 25644 15108 25656
rect 15160 25644 15166 25696
rect 15930 25644 15936 25696
rect 15988 25684 15994 25696
rect 17037 25687 17095 25693
rect 17037 25684 17049 25687
rect 15988 25656 17049 25684
rect 15988 25644 15994 25656
rect 17037 25653 17049 25656
rect 17083 25653 17095 25687
rect 17037 25647 17095 25653
rect 17865 25687 17923 25693
rect 17865 25653 17877 25687
rect 17911 25684 17923 25687
rect 18046 25684 18052 25696
rect 17911 25656 18052 25684
rect 17911 25653 17923 25656
rect 17865 25647 17923 25653
rect 18046 25644 18052 25656
rect 18104 25644 18110 25696
rect 18414 25684 18420 25696
rect 18375 25656 18420 25684
rect 18414 25644 18420 25656
rect 18472 25644 18478 25696
rect 24857 25687 24915 25693
rect 24857 25653 24869 25687
rect 24903 25684 24915 25687
rect 25130 25684 25136 25696
rect 24903 25656 25136 25684
rect 24903 25653 24915 25656
rect 24857 25647 24915 25653
rect 25130 25644 25136 25656
rect 25188 25644 25194 25696
rect 25406 25644 25412 25696
rect 25464 25684 25470 25696
rect 25501 25687 25559 25693
rect 25501 25684 25513 25687
rect 25464 25656 25513 25684
rect 25464 25644 25470 25656
rect 25501 25653 25513 25656
rect 25547 25653 25559 25687
rect 25501 25647 25559 25653
rect 29914 25644 29920 25696
rect 29972 25684 29978 25696
rect 30653 25687 30711 25693
rect 30653 25684 30665 25687
rect 29972 25656 30665 25684
rect 29972 25644 29978 25656
rect 30653 25653 30665 25656
rect 30699 25653 30711 25687
rect 30653 25647 30711 25653
rect 46385 25687 46443 25693
rect 46385 25653 46397 25687
rect 46431 25684 46443 25687
rect 46474 25684 46480 25696
rect 46431 25656 46480 25684
rect 46431 25653 46443 25656
rect 46385 25647 46443 25653
rect 46474 25644 46480 25656
rect 46532 25644 46538 25696
rect 47762 25684 47768 25696
rect 47723 25656 47768 25684
rect 47762 25644 47768 25656
rect 47820 25644 47826 25696
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 11790 25480 11796 25492
rect 11751 25452 11796 25480
rect 11790 25440 11796 25452
rect 11848 25440 11854 25492
rect 16758 25480 16764 25492
rect 16719 25452 16764 25480
rect 16758 25440 16764 25452
rect 16816 25440 16822 25492
rect 17773 25483 17831 25489
rect 17773 25449 17785 25483
rect 17819 25480 17831 25483
rect 17954 25480 17960 25492
rect 17819 25452 17960 25480
rect 17819 25449 17831 25452
rect 17773 25443 17831 25449
rect 17954 25440 17960 25452
rect 18012 25440 18018 25492
rect 18230 25480 18236 25492
rect 18191 25452 18236 25480
rect 18230 25440 18236 25452
rect 18288 25440 18294 25492
rect 22830 25440 22836 25492
rect 22888 25480 22894 25492
rect 22925 25483 22983 25489
rect 22925 25480 22937 25483
rect 22888 25452 22937 25480
rect 22888 25440 22894 25452
rect 22925 25449 22937 25452
rect 22971 25449 22983 25483
rect 22925 25443 22983 25449
rect 24660 25483 24718 25489
rect 24660 25449 24672 25483
rect 24706 25480 24718 25483
rect 25774 25480 25780 25492
rect 24706 25452 25780 25480
rect 24706 25449 24718 25452
rect 24660 25443 24718 25449
rect 25774 25440 25780 25452
rect 25832 25440 25838 25492
rect 30374 25480 30380 25492
rect 29656 25452 30380 25480
rect 11606 25372 11612 25424
rect 11664 25412 11670 25424
rect 12618 25412 12624 25424
rect 11664 25384 12624 25412
rect 11664 25372 11670 25384
rect 12618 25372 12624 25384
rect 12676 25412 12682 25424
rect 13354 25412 13360 25424
rect 12676 25384 13360 25412
rect 12676 25372 12682 25384
rect 13354 25372 13360 25384
rect 13412 25372 13418 25424
rect 16482 25372 16488 25424
rect 16540 25412 16546 25424
rect 17221 25415 17279 25421
rect 17221 25412 17233 25415
rect 16540 25384 17233 25412
rect 16540 25372 16546 25384
rect 17221 25381 17233 25384
rect 17267 25381 17279 25415
rect 17221 25375 17279 25381
rect 8294 25304 8300 25356
rect 8352 25344 8358 25356
rect 9401 25347 9459 25353
rect 9401 25344 9413 25347
rect 8352 25316 9413 25344
rect 8352 25304 8358 25316
rect 9401 25313 9413 25316
rect 9447 25313 9459 25347
rect 14458 25344 14464 25356
rect 9401 25307 9459 25313
rect 11164 25316 12848 25344
rect 14419 25316 14464 25344
rect 8941 25279 8999 25285
rect 8941 25245 8953 25279
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 1949 25143 2007 25149
rect 1949 25109 1961 25143
rect 1995 25140 2007 25143
rect 2038 25140 2044 25152
rect 1995 25112 2044 25140
rect 1995 25109 2007 25112
rect 1949 25103 2007 25109
rect 2038 25100 2044 25112
rect 2096 25100 2102 25152
rect 8956 25140 8984 25239
rect 9122 25208 9128 25220
rect 9083 25180 9128 25208
rect 9122 25168 9128 25180
rect 9180 25168 9186 25220
rect 11164 25140 11192 25316
rect 11425 25279 11483 25285
rect 11425 25245 11437 25279
rect 11471 25276 11483 25279
rect 11698 25276 11704 25288
rect 11471 25248 11704 25276
rect 11471 25245 11483 25248
rect 11425 25239 11483 25245
rect 11698 25236 11704 25248
rect 11756 25276 11762 25288
rect 12342 25276 12348 25288
rect 11756 25248 12348 25276
rect 11756 25236 11762 25248
rect 12342 25236 12348 25248
rect 12400 25276 12406 25288
rect 12713 25279 12771 25285
rect 12713 25276 12725 25279
rect 12400 25248 12725 25276
rect 12400 25236 12406 25248
rect 12713 25245 12725 25248
rect 12759 25245 12771 25279
rect 12713 25239 12771 25245
rect 11241 25211 11299 25217
rect 11241 25177 11253 25211
rect 11287 25208 11299 25211
rect 12066 25208 12072 25220
rect 11287 25180 12072 25208
rect 11287 25177 11299 25180
rect 11241 25171 11299 25177
rect 12066 25168 12072 25180
rect 12124 25168 12130 25220
rect 12437 25211 12495 25217
rect 12437 25177 12449 25211
rect 12483 25208 12495 25211
rect 12820 25208 12848 25316
rect 14458 25304 14464 25316
rect 14516 25304 14522 25356
rect 17236 25344 17264 25375
rect 25682 25372 25688 25424
rect 25740 25412 25746 25424
rect 26145 25415 26203 25421
rect 26145 25412 26157 25415
rect 25740 25384 26157 25412
rect 25740 25372 25746 25384
rect 26145 25381 26157 25384
rect 26191 25381 26203 25415
rect 26145 25375 26203 25381
rect 24397 25347 24455 25353
rect 17236 25316 18644 25344
rect 14182 25276 14188 25288
rect 14143 25248 14188 25276
rect 14182 25236 14188 25248
rect 14240 25236 14246 25288
rect 16482 25276 16488 25288
rect 16443 25248 16488 25276
rect 16482 25236 16488 25248
rect 16540 25236 16546 25288
rect 16577 25279 16635 25285
rect 16577 25245 16589 25279
rect 16623 25276 16635 25279
rect 17589 25279 17647 25285
rect 16623 25248 17540 25276
rect 16623 25245 16635 25248
rect 16577 25239 16635 25245
rect 13170 25208 13176 25220
rect 12483 25180 13176 25208
rect 12483 25177 12495 25180
rect 12437 25171 12495 25177
rect 13170 25168 13176 25180
rect 13228 25168 13234 25220
rect 15102 25168 15108 25220
rect 15160 25168 15166 25220
rect 11514 25140 11520 25152
rect 8956 25112 11192 25140
rect 11475 25112 11520 25140
rect 11514 25100 11520 25112
rect 11572 25100 11578 25152
rect 11606 25100 11612 25152
rect 11664 25140 11670 25152
rect 12084 25140 12112 25168
rect 17512 25152 17540 25248
rect 17589 25245 17601 25279
rect 17635 25276 17647 25279
rect 18506 25276 18512 25288
rect 17635 25248 17816 25276
rect 18467 25248 18512 25276
rect 17635 25245 17647 25248
rect 17589 25239 17647 25245
rect 12621 25143 12679 25149
rect 12621 25140 12633 25143
rect 11664 25112 11709 25140
rect 12084 25112 12633 25140
rect 11664 25100 11670 25112
rect 12621 25109 12633 25112
rect 12667 25109 12679 25143
rect 12621 25103 12679 25109
rect 12710 25100 12716 25152
rect 12768 25140 12774 25152
rect 12805 25143 12863 25149
rect 12805 25140 12817 25143
rect 12768 25112 12817 25140
rect 12768 25100 12774 25112
rect 12805 25109 12817 25112
rect 12851 25109 12863 25143
rect 12805 25103 12863 25109
rect 12989 25143 13047 25149
rect 12989 25109 13001 25143
rect 13035 25140 13047 25143
rect 13538 25140 13544 25152
rect 13035 25112 13544 25140
rect 13035 25109 13047 25112
rect 12989 25103 13047 25109
rect 13538 25100 13544 25112
rect 13596 25100 13602 25152
rect 13998 25100 14004 25152
rect 14056 25140 14062 25152
rect 15933 25143 15991 25149
rect 15933 25140 15945 25143
rect 14056 25112 15945 25140
rect 14056 25100 14062 25112
rect 15933 25109 15945 25112
rect 15979 25140 15991 25143
rect 16390 25140 16396 25152
rect 15979 25112 16396 25140
rect 15979 25109 15991 25112
rect 15933 25103 15991 25109
rect 16390 25100 16396 25112
rect 16448 25100 16454 25152
rect 16482 25100 16488 25152
rect 16540 25140 16546 25152
rect 17405 25143 17463 25149
rect 17405 25140 17417 25143
rect 16540 25112 17417 25140
rect 16540 25100 16546 25112
rect 17405 25109 17417 25112
rect 17451 25109 17463 25143
rect 17405 25103 17463 25109
rect 17494 25100 17500 25152
rect 17552 25140 17558 25152
rect 17788 25140 17816 25248
rect 18506 25236 18512 25248
rect 18564 25236 18570 25288
rect 18233 25211 18291 25217
rect 18233 25177 18245 25211
rect 18279 25208 18291 25211
rect 18616 25208 18644 25316
rect 24397 25313 24409 25347
rect 24443 25344 24455 25347
rect 27154 25344 27160 25356
rect 24443 25316 27160 25344
rect 24443 25313 24455 25316
rect 24397 25307 24455 25313
rect 27154 25304 27160 25316
rect 27212 25344 27218 25356
rect 29656 25353 29684 25452
rect 30374 25440 30380 25452
rect 30432 25440 30438 25492
rect 31389 25483 31447 25489
rect 31389 25449 31401 25483
rect 31435 25480 31447 25483
rect 31570 25480 31576 25492
rect 31435 25452 31576 25480
rect 31435 25449 31447 25452
rect 31389 25443 31447 25449
rect 31570 25440 31576 25452
rect 31628 25440 31634 25492
rect 29641 25347 29699 25353
rect 29641 25344 29653 25347
rect 27212 25316 29653 25344
rect 27212 25304 27218 25316
rect 29641 25313 29653 25316
rect 29687 25313 29699 25347
rect 29914 25344 29920 25356
rect 29875 25316 29920 25344
rect 29641 25307 29699 25313
rect 29914 25304 29920 25316
rect 29972 25304 29978 25356
rect 46474 25344 46480 25356
rect 46435 25316 46480 25344
rect 46474 25304 46480 25316
rect 46532 25304 46538 25356
rect 48130 25344 48136 25356
rect 48091 25316 48136 25344
rect 48130 25304 48136 25316
rect 48188 25304 48194 25356
rect 22833 25279 22891 25285
rect 22833 25245 22845 25279
rect 22879 25276 22891 25279
rect 23382 25276 23388 25288
rect 22879 25248 23388 25276
rect 22879 25245 22891 25248
rect 22833 25239 22891 25245
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 45830 25236 45836 25288
rect 45888 25276 45894 25288
rect 46293 25279 46351 25285
rect 46293 25276 46305 25279
rect 45888 25248 46305 25276
rect 45888 25236 45894 25248
rect 46293 25245 46305 25248
rect 46339 25245 46351 25279
rect 46293 25239 46351 25245
rect 19334 25208 19340 25220
rect 18279 25180 19340 25208
rect 18279 25177 18291 25180
rect 18233 25171 18291 25177
rect 19334 25168 19340 25180
rect 19392 25168 19398 25220
rect 25130 25168 25136 25220
rect 25188 25168 25194 25220
rect 30926 25168 30932 25220
rect 30984 25168 30990 25220
rect 17862 25140 17868 25152
rect 17552 25112 17597 25140
rect 17775 25112 17868 25140
rect 17552 25100 17558 25112
rect 17862 25100 17868 25112
rect 17920 25140 17926 25152
rect 18417 25143 18475 25149
rect 18417 25140 18429 25143
rect 17920 25112 18429 25140
rect 17920 25100 17926 25112
rect 18417 25109 18429 25112
rect 18463 25109 18475 25143
rect 18417 25103 18475 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 8849 24939 8907 24945
rect 8849 24905 8861 24939
rect 8895 24936 8907 24939
rect 9122 24936 9128 24948
rect 8895 24908 9128 24936
rect 8895 24905 8907 24908
rect 8849 24899 8907 24905
rect 9122 24896 9128 24908
rect 9180 24896 9186 24948
rect 11514 24896 11520 24948
rect 11572 24936 11578 24948
rect 11609 24939 11667 24945
rect 11609 24936 11621 24939
rect 11572 24908 11621 24936
rect 11572 24896 11578 24908
rect 11609 24905 11621 24908
rect 11655 24936 11667 24939
rect 12710 24936 12716 24948
rect 11655 24908 12716 24936
rect 11655 24905 11667 24908
rect 11609 24899 11667 24905
rect 12710 24896 12716 24908
rect 12768 24896 12774 24948
rect 13538 24896 13544 24948
rect 13596 24936 13602 24948
rect 13596 24908 14141 24936
rect 13596 24896 13602 24908
rect 11790 24868 11796 24880
rect 11440 24840 11796 24868
rect 8757 24803 8815 24809
rect 8757 24769 8769 24803
rect 8803 24800 8815 24803
rect 8938 24800 8944 24812
rect 8803 24772 8944 24800
rect 8803 24769 8815 24772
rect 8757 24763 8815 24769
rect 8938 24760 8944 24772
rect 8996 24760 9002 24812
rect 9677 24803 9735 24809
rect 9677 24769 9689 24803
rect 9723 24769 9735 24803
rect 9677 24763 9735 24769
rect 9861 24803 9919 24809
rect 9861 24769 9873 24803
rect 9907 24769 9919 24803
rect 9861 24763 9919 24769
rect 10505 24803 10563 24809
rect 10505 24769 10517 24803
rect 10551 24800 10563 24803
rect 10686 24800 10692 24812
rect 10551 24772 10692 24800
rect 10551 24769 10563 24772
rect 10505 24763 10563 24769
rect 9692 24664 9720 24763
rect 9876 24732 9904 24763
rect 10686 24760 10692 24772
rect 10744 24760 10750 24812
rect 11440 24732 11468 24840
rect 11790 24828 11796 24840
rect 11848 24828 11854 24880
rect 12802 24868 12808 24880
rect 12763 24840 12808 24868
rect 12802 24828 12808 24840
rect 12860 24828 12866 24880
rect 14113 24868 14141 24908
rect 14182 24896 14188 24948
rect 14240 24936 14246 24948
rect 14921 24939 14979 24945
rect 14921 24936 14933 24939
rect 14240 24908 14933 24936
rect 14240 24896 14246 24908
rect 14921 24905 14933 24908
rect 14967 24905 14979 24939
rect 14921 24899 14979 24905
rect 16758 24896 16764 24948
rect 16816 24936 16822 24948
rect 17037 24939 17095 24945
rect 17037 24936 17049 24939
rect 16816 24908 17049 24936
rect 16816 24896 16822 24908
rect 17037 24905 17049 24908
rect 17083 24905 17095 24939
rect 17037 24899 17095 24905
rect 19334 24896 19340 24948
rect 19392 24936 19398 24948
rect 19797 24939 19855 24945
rect 19797 24936 19809 24939
rect 19392 24908 19809 24936
rect 19392 24896 19398 24908
rect 19797 24905 19809 24908
rect 19843 24905 19855 24939
rect 19797 24899 19855 24905
rect 23109 24939 23167 24945
rect 23109 24905 23121 24939
rect 23155 24936 23167 24939
rect 23382 24936 23388 24948
rect 23155 24908 23388 24936
rect 23155 24905 23167 24908
rect 23109 24899 23167 24905
rect 23382 24896 23388 24908
rect 23440 24896 23446 24948
rect 26142 24936 26148 24948
rect 26103 24908 26148 24936
rect 26142 24896 26148 24908
rect 26200 24896 26206 24948
rect 16945 24871 17003 24877
rect 16945 24868 16957 24871
rect 14113 24840 16957 24868
rect 16945 24837 16957 24840
rect 16991 24868 17003 24871
rect 18325 24871 18383 24877
rect 16991 24840 17080 24868
rect 16991 24837 17003 24840
rect 16945 24831 17003 24837
rect 17052 24812 17080 24840
rect 18325 24837 18337 24871
rect 18371 24868 18383 24871
rect 18414 24868 18420 24880
rect 18371 24840 18420 24868
rect 18371 24837 18383 24840
rect 18325 24831 18383 24837
rect 18414 24828 18420 24840
rect 18472 24828 18478 24880
rect 25406 24828 25412 24880
rect 25464 24828 25470 24880
rect 39577 24871 39635 24877
rect 39577 24868 39589 24871
rect 39408 24840 39589 24868
rect 11517 24803 11575 24809
rect 11517 24769 11529 24803
rect 11563 24800 11575 24803
rect 11606 24800 11612 24812
rect 11563 24772 11612 24800
rect 11563 24769 11575 24772
rect 11517 24763 11575 24769
rect 11606 24760 11612 24772
rect 11664 24760 11670 24812
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24800 11943 24803
rect 12066 24800 12072 24812
rect 11931 24772 12072 24800
rect 11931 24769 11943 24772
rect 11885 24763 11943 24769
rect 12066 24760 12072 24772
rect 12124 24760 12130 24812
rect 12526 24800 12532 24812
rect 12487 24772 12532 24800
rect 12526 24760 12532 24772
rect 12584 24760 12590 24812
rect 14182 24800 14188 24812
rect 13938 24772 14188 24800
rect 14182 24760 14188 24772
rect 14240 24760 14246 24812
rect 14734 24800 14740 24812
rect 14695 24772 14740 24800
rect 14734 24760 14740 24772
rect 14792 24760 14798 24812
rect 15930 24800 15936 24812
rect 15891 24772 15936 24800
rect 15930 24760 15936 24772
rect 15988 24760 15994 24812
rect 16390 24760 16396 24812
rect 16448 24800 16454 24812
rect 16669 24803 16727 24809
rect 16669 24800 16681 24803
rect 16448 24772 16681 24800
rect 16448 24760 16454 24772
rect 16669 24769 16681 24772
rect 16715 24769 16727 24803
rect 16850 24800 16856 24812
rect 16811 24772 16856 24800
rect 16669 24763 16727 24769
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 17034 24760 17040 24812
rect 17092 24760 17098 24812
rect 18046 24800 18052 24812
rect 18007 24772 18052 24800
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 20257 24803 20315 24809
rect 11698 24732 11704 24744
rect 9876 24704 11468 24732
rect 11659 24704 11704 24732
rect 11698 24692 11704 24704
rect 11756 24692 11762 24744
rect 13170 24692 13176 24744
rect 13228 24732 13234 24744
rect 14277 24735 14335 24741
rect 14277 24732 14289 24735
rect 13228 24704 14289 24732
rect 13228 24692 13234 24704
rect 14277 24701 14289 24704
rect 14323 24701 14335 24735
rect 14277 24695 14335 24701
rect 11885 24667 11943 24673
rect 11885 24664 11897 24667
rect 9692 24636 11897 24664
rect 11885 24633 11897 24636
rect 11931 24633 11943 24667
rect 15948 24664 15976 24760
rect 19444 24732 19472 24786
rect 20257 24769 20269 24803
rect 20303 24800 20315 24803
rect 20901 24803 20959 24809
rect 20303 24772 20484 24800
rect 20303 24769 20315 24772
rect 20257 24763 20315 24769
rect 20349 24735 20407 24741
rect 20349 24732 20361 24735
rect 19444 24704 20361 24732
rect 20349 24701 20361 24704
rect 20395 24701 20407 24735
rect 20349 24695 20407 24701
rect 11885 24627 11943 24633
rect 14113 24636 15976 24664
rect 9674 24596 9680 24608
rect 9635 24568 9680 24596
rect 9674 24556 9680 24568
rect 9732 24556 9738 24608
rect 10318 24596 10324 24608
rect 10279 24568 10324 24596
rect 10318 24556 10324 24568
rect 10376 24556 10382 24608
rect 13354 24556 13360 24608
rect 13412 24596 13418 24608
rect 14113 24596 14141 24636
rect 19518 24624 19524 24676
rect 19576 24664 19582 24676
rect 20456 24664 20484 24772
rect 20901 24769 20913 24803
rect 20947 24769 20959 24803
rect 20901 24763 20959 24769
rect 22189 24803 22247 24809
rect 22189 24769 22201 24803
rect 22235 24800 22247 24803
rect 22922 24800 22928 24812
rect 22235 24772 22928 24800
rect 22235 24769 22247 24772
rect 22189 24763 22247 24769
rect 20530 24692 20536 24744
rect 20588 24732 20594 24744
rect 20916 24732 20944 24763
rect 22922 24760 22928 24772
rect 22980 24760 22986 24812
rect 27617 24803 27675 24809
rect 27617 24769 27629 24803
rect 27663 24800 27675 24803
rect 28258 24800 28264 24812
rect 27663 24772 28264 24800
rect 27663 24769 27675 24772
rect 27617 24763 27675 24769
rect 28258 24760 28264 24772
rect 28316 24760 28322 24812
rect 30282 24760 30288 24812
rect 30340 24800 30346 24812
rect 30653 24803 30711 24809
rect 30653 24800 30665 24803
rect 30340 24772 30665 24800
rect 30340 24760 30346 24772
rect 30653 24769 30665 24772
rect 30699 24769 30711 24803
rect 30653 24763 30711 24769
rect 30745 24803 30803 24809
rect 30745 24769 30757 24803
rect 30791 24800 30803 24803
rect 30926 24800 30932 24812
rect 30791 24772 30932 24800
rect 30791 24769 30803 24772
rect 30745 24763 30803 24769
rect 30926 24760 30932 24772
rect 30984 24760 30990 24812
rect 38746 24800 38752 24812
rect 38707 24772 38752 24800
rect 38746 24760 38752 24772
rect 38804 24760 38810 24812
rect 38841 24803 38899 24809
rect 38841 24769 38853 24803
rect 38887 24800 38899 24803
rect 39408 24800 39436 24840
rect 39577 24837 39589 24840
rect 39623 24837 39635 24871
rect 39577 24831 39635 24837
rect 45186 24800 45192 24812
rect 38887 24772 39436 24800
rect 45147 24772 45192 24800
rect 38887 24769 38899 24772
rect 38841 24763 38899 24769
rect 45186 24760 45192 24772
rect 45244 24760 45250 24812
rect 46750 24760 46756 24812
rect 46808 24800 46814 24812
rect 47578 24800 47584 24812
rect 46808 24772 47584 24800
rect 46808 24760 46814 24772
rect 47578 24760 47584 24772
rect 47636 24760 47642 24812
rect 20588 24704 20944 24732
rect 20588 24692 20594 24704
rect 21818 24692 21824 24744
rect 21876 24732 21882 24744
rect 24397 24735 24455 24741
rect 24397 24732 24409 24735
rect 21876 24704 24409 24732
rect 21876 24692 21882 24704
rect 24397 24701 24409 24704
rect 24443 24701 24455 24735
rect 24670 24732 24676 24744
rect 24631 24704 24676 24732
rect 24397 24695 24455 24701
rect 24670 24692 24676 24704
rect 24728 24692 24734 24744
rect 25038 24692 25044 24744
rect 25096 24732 25102 24744
rect 39393 24735 39451 24741
rect 25096 24704 36584 24732
rect 25096 24692 25102 24704
rect 22094 24664 22100 24676
rect 19576 24636 22100 24664
rect 19576 24624 19582 24636
rect 22094 24624 22100 24636
rect 22152 24624 22158 24676
rect 26418 24624 26424 24676
rect 26476 24664 26482 24676
rect 36556 24664 36584 24704
rect 39393 24701 39405 24735
rect 39439 24732 39451 24735
rect 40586 24732 40592 24744
rect 39439 24704 40592 24732
rect 39439 24701 39451 24704
rect 39393 24695 39451 24701
rect 40586 24692 40592 24704
rect 40644 24692 40650 24744
rect 40696 24704 40908 24732
rect 40696 24664 40724 24704
rect 26476 24636 31754 24664
rect 36556 24636 40724 24664
rect 40880 24664 40908 24704
rect 40954 24692 40960 24744
rect 41012 24732 41018 24744
rect 45370 24732 45376 24744
rect 41012 24704 41057 24732
rect 45331 24704 45376 24732
rect 41012 24692 41018 24704
rect 45370 24692 45376 24704
rect 45428 24692 45434 24744
rect 46842 24732 46848 24744
rect 46803 24704 46848 24732
rect 46842 24692 46848 24704
rect 46900 24692 46906 24744
rect 45554 24664 45560 24676
rect 40880 24636 45560 24664
rect 26476 24624 26482 24636
rect 16022 24596 16028 24608
rect 13412 24568 14141 24596
rect 15983 24568 16028 24596
rect 13412 24556 13418 24568
rect 16022 24556 16028 24568
rect 16080 24556 16086 24608
rect 17126 24556 17132 24608
rect 17184 24596 17190 24608
rect 17221 24599 17279 24605
rect 17221 24596 17233 24599
rect 17184 24568 17233 24596
rect 17184 24556 17190 24568
rect 17221 24565 17233 24568
rect 17267 24565 17279 24599
rect 17221 24559 17279 24565
rect 20438 24556 20444 24608
rect 20496 24596 20502 24608
rect 20993 24599 21051 24605
rect 20993 24596 21005 24599
rect 20496 24568 21005 24596
rect 20496 24556 20502 24568
rect 20993 24565 21005 24568
rect 21039 24565 21051 24599
rect 22370 24596 22376 24608
rect 22283 24568 22376 24596
rect 20993 24559 21051 24565
rect 22370 24556 22376 24568
rect 22428 24596 22434 24608
rect 23014 24596 23020 24608
rect 22428 24568 23020 24596
rect 22428 24556 22434 24568
rect 23014 24556 23020 24568
rect 23072 24556 23078 24608
rect 27338 24556 27344 24608
rect 27396 24596 27402 24608
rect 27709 24599 27767 24605
rect 27709 24596 27721 24599
rect 27396 24568 27721 24596
rect 27396 24556 27402 24568
rect 27709 24565 27721 24568
rect 27755 24565 27767 24599
rect 28350 24596 28356 24608
rect 28311 24568 28356 24596
rect 27709 24559 27767 24565
rect 28350 24556 28356 24568
rect 28408 24556 28414 24608
rect 31726 24596 31754 24636
rect 45554 24624 45560 24636
rect 45612 24624 45618 24676
rect 40954 24596 40960 24608
rect 31726 24568 40960 24596
rect 40954 24556 40960 24568
rect 41012 24556 41018 24608
rect 46474 24556 46480 24608
rect 46532 24596 46538 24608
rect 47673 24599 47731 24605
rect 47673 24596 47685 24599
rect 46532 24568 47685 24596
rect 46532 24556 46538 24568
rect 47673 24565 47685 24568
rect 47719 24565 47731 24599
rect 47673 24559 47731 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 10778 24352 10784 24404
rect 10836 24392 10842 24404
rect 13446 24392 13452 24404
rect 10836 24364 11652 24392
rect 13407 24364 13452 24392
rect 10836 24352 10842 24364
rect 11624 24336 11652 24364
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 14182 24392 14188 24404
rect 14143 24364 14188 24392
rect 14182 24352 14188 24364
rect 14240 24352 14246 24404
rect 47486 24392 47492 24404
rect 45756 24364 47492 24392
rect 9674 24284 9680 24336
rect 9732 24324 9738 24336
rect 9732 24296 10456 24324
rect 9732 24284 9738 24296
rect 10318 24256 10324 24268
rect 10279 24228 10324 24256
rect 10318 24216 10324 24228
rect 10376 24216 10382 24268
rect 10428 24256 10456 24296
rect 11606 24284 11612 24336
rect 11664 24324 11670 24336
rect 16022 24324 16028 24336
rect 11664 24296 16028 24324
rect 11664 24284 11670 24296
rect 16022 24284 16028 24296
rect 16080 24324 16086 24336
rect 18506 24324 18512 24336
rect 16080 24296 18512 24324
rect 16080 24284 16086 24296
rect 10597 24259 10655 24265
rect 10597 24256 10609 24259
rect 10428 24228 10609 24256
rect 10597 24225 10609 24228
rect 10643 24225 10655 24259
rect 13722 24256 13728 24268
rect 10597 24219 10655 24225
rect 12544 24228 13728 24256
rect 12434 24148 12440 24200
rect 12492 24188 12498 24200
rect 12544 24197 12572 24228
rect 13722 24216 13728 24228
rect 13780 24256 13786 24268
rect 16577 24259 16635 24265
rect 13780 24228 14136 24256
rect 13780 24216 13786 24228
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 12492 24160 12541 24188
rect 12492 24148 12498 24160
rect 12529 24157 12541 24160
rect 12575 24157 12587 24191
rect 13354 24188 13360 24200
rect 13315 24160 13360 24188
rect 12529 24151 12587 24157
rect 13354 24148 13360 24160
rect 13412 24148 13418 24200
rect 13538 24188 13544 24200
rect 13499 24160 13544 24188
rect 13538 24148 13544 24160
rect 13596 24148 13602 24200
rect 14108 24197 14136 24228
rect 16577 24225 16589 24259
rect 16623 24256 16635 24259
rect 16850 24256 16856 24268
rect 16623 24228 16856 24256
rect 16623 24225 16635 24228
rect 16577 24219 16635 24225
rect 16850 24216 16856 24228
rect 16908 24216 16914 24268
rect 17129 24259 17187 24265
rect 17129 24225 17141 24259
rect 17175 24256 17187 24259
rect 17175 24228 17908 24256
rect 17175 24225 17187 24228
rect 17129 24219 17187 24225
rect 17880 24200 17908 24228
rect 14093 24191 14151 24197
rect 14093 24157 14105 24191
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 16666 24148 16672 24200
rect 16724 24188 16730 24200
rect 17589 24191 17647 24197
rect 17589 24188 17601 24191
rect 16724 24160 17601 24188
rect 16724 24148 16730 24160
rect 17589 24157 17601 24160
rect 17635 24157 17647 24191
rect 17589 24151 17647 24157
rect 17862 24148 17868 24200
rect 17920 24188 17926 24200
rect 18064 24197 18092 24296
rect 18506 24284 18512 24296
rect 18564 24284 18570 24336
rect 45646 24324 45652 24336
rect 22112 24296 45652 24324
rect 20438 24256 20444 24268
rect 20399 24228 20444 24256
rect 20438 24216 20444 24228
rect 20496 24216 20502 24268
rect 22112 24265 22140 24296
rect 45646 24284 45652 24296
rect 45704 24284 45710 24336
rect 22097 24259 22155 24265
rect 22097 24225 22109 24259
rect 22143 24225 22155 24259
rect 27338 24256 27344 24268
rect 27299 24228 27344 24256
rect 22097 24219 22155 24225
rect 27338 24216 27344 24228
rect 27396 24216 27402 24268
rect 28997 24259 29055 24265
rect 28997 24225 29009 24259
rect 29043 24256 29055 24259
rect 37274 24256 37280 24268
rect 29043 24228 37280 24256
rect 29043 24225 29055 24228
rect 28997 24219 29055 24225
rect 37274 24216 37280 24228
rect 37332 24216 37338 24268
rect 45756 24256 45784 24364
rect 47486 24352 47492 24364
rect 47544 24352 47550 24404
rect 47762 24324 47768 24336
rect 46308 24296 47768 24324
rect 46308 24265 46336 24296
rect 47762 24284 47768 24296
rect 47820 24284 47826 24336
rect 41386 24228 45784 24256
rect 46293 24259 46351 24265
rect 17957 24191 18015 24197
rect 17957 24188 17969 24191
rect 17920 24160 17969 24188
rect 17920 24148 17926 24160
rect 17957 24157 17969 24160
rect 18003 24157 18015 24191
rect 17957 24151 18015 24157
rect 18049 24191 18107 24197
rect 18049 24157 18061 24191
rect 18095 24157 18107 24191
rect 19518 24188 19524 24200
rect 19479 24160 19524 24188
rect 18049 24151 18107 24157
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 20254 24188 20260 24200
rect 20215 24160 20260 24188
rect 20254 24148 20260 24160
rect 20312 24148 20318 24200
rect 22649 24191 22707 24197
rect 22649 24157 22661 24191
rect 22695 24188 22707 24191
rect 22922 24188 22928 24200
rect 22695 24160 22928 24188
rect 22695 24157 22707 24160
rect 22649 24151 22707 24157
rect 22922 24148 22928 24160
rect 22980 24148 22986 24200
rect 23382 24148 23388 24200
rect 23440 24188 23446 24200
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 23440 24160 24409 24188
rect 23440 24148 23446 24160
rect 24397 24157 24409 24160
rect 24443 24157 24455 24191
rect 27154 24188 27160 24200
rect 27115 24160 27160 24188
rect 24397 24151 24455 24157
rect 27154 24148 27160 24160
rect 27212 24148 27218 24200
rect 12621 24123 12679 24129
rect 12621 24120 12633 24123
rect 11822 24092 12633 24120
rect 12621 24089 12633 24092
rect 12667 24089 12679 24123
rect 12621 24083 12679 24089
rect 16390 24080 16396 24132
rect 16448 24120 16454 24132
rect 16853 24123 16911 24129
rect 16853 24120 16865 24123
rect 16448 24092 16865 24120
rect 16448 24080 16454 24092
rect 16853 24089 16865 24092
rect 16899 24089 16911 24123
rect 16853 24083 16911 24089
rect 16945 24123 17003 24129
rect 16945 24089 16957 24123
rect 16991 24120 17003 24123
rect 17034 24120 17040 24132
rect 16991 24092 17040 24120
rect 16991 24089 17003 24092
rect 16945 24083 17003 24089
rect 17034 24080 17040 24092
rect 17092 24080 17098 24132
rect 39206 24080 39212 24132
rect 39264 24120 39270 24132
rect 41386 24120 41414 24228
rect 46293 24225 46305 24259
rect 46339 24225 46351 24259
rect 46474 24256 46480 24268
rect 46435 24228 46480 24256
rect 46293 24219 46351 24225
rect 46474 24216 46480 24228
rect 46532 24216 46538 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 42978 24148 42984 24200
rect 43036 24188 43042 24200
rect 43073 24191 43131 24197
rect 43073 24188 43085 24191
rect 43036 24160 43085 24188
rect 43036 24148 43042 24160
rect 43073 24157 43085 24160
rect 43119 24157 43131 24191
rect 43073 24151 43131 24157
rect 43257 24191 43315 24197
rect 43257 24157 43269 24191
rect 43303 24157 43315 24191
rect 43257 24151 43315 24157
rect 45833 24191 45891 24197
rect 45833 24157 45845 24191
rect 45879 24188 45891 24191
rect 45922 24188 45928 24200
rect 45879 24160 45928 24188
rect 45879 24157 45891 24160
rect 45833 24151 45891 24157
rect 39264 24092 41414 24120
rect 39264 24080 39270 24092
rect 42794 24080 42800 24132
rect 42852 24120 42858 24132
rect 43272 24120 43300 24151
rect 45922 24148 45928 24160
rect 45980 24148 45986 24200
rect 42852 24092 43300 24120
rect 42852 24080 42858 24092
rect 12066 24052 12072 24064
rect 12027 24024 12072 24052
rect 12066 24012 12072 24024
rect 12124 24012 12130 24064
rect 16758 24052 16764 24064
rect 16719 24024 16764 24052
rect 16758 24012 16764 24024
rect 16816 24012 16822 24064
rect 17862 24052 17868 24064
rect 17823 24024 17868 24052
rect 17862 24012 17868 24024
rect 17920 24012 17926 24064
rect 19426 24012 19432 24064
rect 19484 24052 19490 24064
rect 19613 24055 19671 24061
rect 19613 24052 19625 24055
rect 19484 24024 19625 24052
rect 19484 24012 19490 24024
rect 19613 24021 19625 24024
rect 19659 24021 19671 24055
rect 22738 24052 22744 24064
rect 22699 24024 22744 24052
rect 19613 24015 19671 24021
rect 22738 24012 22744 24024
rect 22796 24012 22802 24064
rect 24118 24012 24124 24064
rect 24176 24052 24182 24064
rect 24489 24055 24547 24061
rect 24489 24052 24501 24055
rect 24176 24024 24501 24052
rect 24176 24012 24182 24024
rect 24489 24021 24501 24024
rect 24535 24021 24547 24055
rect 24489 24015 24547 24021
rect 26050 24012 26056 24064
rect 26108 24052 26114 24064
rect 41230 24052 41236 24064
rect 26108 24024 41236 24052
rect 26108 24012 26114 24024
rect 41230 24012 41236 24024
rect 41288 24012 41294 24064
rect 43162 24052 43168 24064
rect 43123 24024 43168 24052
rect 43162 24012 43168 24024
rect 43220 24012 43226 24064
rect 45649 24055 45707 24061
rect 45649 24021 45661 24055
rect 45695 24052 45707 24055
rect 47578 24052 47584 24064
rect 45695 24024 47584 24052
rect 45695 24021 45707 24024
rect 45649 24015 45707 24021
rect 47578 24012 47584 24024
rect 47636 24012 47642 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 3602 23808 3608 23860
rect 3660 23848 3666 23860
rect 25590 23848 25596 23860
rect 3660 23820 25596 23848
rect 3660 23808 3666 23820
rect 25590 23808 25596 23820
rect 25648 23808 25654 23860
rect 26329 23851 26387 23857
rect 26329 23848 26341 23851
rect 26160 23820 26341 23848
rect 12066 23780 12072 23792
rect 8404 23752 12072 23780
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 8404 23721 8432 23752
rect 12066 23740 12072 23752
rect 12124 23740 12130 23792
rect 16666 23780 16672 23792
rect 16627 23752 16672 23780
rect 16666 23740 16672 23752
rect 16724 23740 16730 23792
rect 16868 23752 17632 23780
rect 16868 23724 16896 23752
rect 8389 23715 8447 23721
rect 8389 23681 8401 23715
rect 8435 23681 8447 23715
rect 8389 23675 8447 23681
rect 14182 23672 14188 23724
rect 14240 23712 14246 23724
rect 14553 23715 14611 23721
rect 14553 23712 14565 23715
rect 14240 23684 14565 23712
rect 14240 23672 14246 23684
rect 14553 23681 14565 23684
rect 14599 23681 14611 23715
rect 16850 23712 16856 23724
rect 16763 23684 16856 23712
rect 14553 23675 14611 23681
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23681 17095 23715
rect 17037 23675 17095 23681
rect 8570 23644 8576 23656
rect 8531 23616 8576 23644
rect 8570 23604 8576 23616
rect 8628 23604 8634 23656
rect 9766 23644 9772 23656
rect 9727 23616 9772 23644
rect 9766 23604 9772 23616
rect 9824 23604 9830 23656
rect 16574 23604 16580 23656
rect 16632 23644 16638 23656
rect 16758 23644 16764 23656
rect 16632 23616 16764 23644
rect 16632 23604 16638 23616
rect 16758 23604 16764 23616
rect 16816 23644 16822 23656
rect 17052 23644 17080 23675
rect 17126 23672 17132 23724
rect 17184 23712 17190 23724
rect 17184 23684 17229 23712
rect 17184 23672 17190 23684
rect 16816 23616 17080 23644
rect 16816 23604 16822 23616
rect 6886 23548 12434 23576
rect 1949 23511 2007 23517
rect 1949 23477 1961 23511
rect 1995 23508 2007 23511
rect 6886 23508 6914 23548
rect 1995 23480 6914 23508
rect 12406 23508 12434 23548
rect 13722 23536 13728 23588
rect 13780 23576 13786 23588
rect 14737 23579 14795 23585
rect 14737 23576 14749 23579
rect 13780 23548 14749 23576
rect 13780 23536 13786 23548
rect 14737 23545 14749 23548
rect 14783 23545 14795 23579
rect 17604 23576 17632 23752
rect 17862 23740 17868 23792
rect 17920 23780 17926 23792
rect 18325 23783 18383 23789
rect 18325 23780 18337 23783
rect 17920 23752 18337 23780
rect 17920 23740 17926 23752
rect 18325 23749 18337 23752
rect 18371 23749 18383 23783
rect 18325 23743 18383 23749
rect 20162 23740 20168 23792
rect 20220 23780 20226 23792
rect 20717 23783 20775 23789
rect 20717 23780 20729 23783
rect 20220 23752 20729 23780
rect 20220 23740 20226 23752
rect 20717 23749 20729 23752
rect 20763 23780 20775 23783
rect 20806 23780 20812 23792
rect 20763 23752 20812 23780
rect 20763 23749 20775 23752
rect 20717 23743 20775 23749
rect 20806 23740 20812 23752
rect 20864 23740 20870 23792
rect 26050 23780 26056 23792
rect 22066 23752 26056 23780
rect 19426 23672 19432 23724
rect 19484 23672 19490 23724
rect 19886 23672 19892 23724
rect 19944 23712 19950 23724
rect 20349 23715 20407 23721
rect 20349 23712 20361 23715
rect 19944 23684 20361 23712
rect 19944 23672 19950 23684
rect 20349 23681 20361 23684
rect 20395 23712 20407 23715
rect 21913 23715 21971 23721
rect 21913 23712 21925 23715
rect 20395 23684 21925 23712
rect 20395 23681 20407 23684
rect 20349 23675 20407 23681
rect 21913 23681 21925 23684
rect 21959 23712 21971 23715
rect 22066 23712 22094 23752
rect 26050 23740 26056 23752
rect 26108 23740 26114 23792
rect 23017 23715 23075 23721
rect 23017 23712 23029 23715
rect 21959 23684 22094 23712
rect 22296 23684 23029 23712
rect 21959 23681 21971 23684
rect 21913 23675 21971 23681
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 18046 23604 18052 23616
rect 18104 23604 18110 23656
rect 19797 23647 19855 23653
rect 19797 23644 19809 23647
rect 18156 23616 19809 23644
rect 18156 23576 18184 23616
rect 19797 23613 19809 23616
rect 19843 23644 19855 23647
rect 20254 23644 20260 23656
rect 19843 23616 20260 23644
rect 19843 23613 19855 23616
rect 19797 23607 19855 23613
rect 20254 23604 20260 23616
rect 20312 23604 20318 23656
rect 22094 23604 22100 23656
rect 22152 23644 22158 23656
rect 22296 23644 22324 23684
rect 23017 23681 23029 23684
rect 23063 23681 23075 23715
rect 23017 23675 23075 23681
rect 25317 23715 25375 23721
rect 25317 23681 25329 23715
rect 25363 23712 25375 23715
rect 26160 23712 26188 23820
rect 26329 23817 26341 23820
rect 26375 23848 26387 23851
rect 28258 23848 28264 23860
rect 26375 23820 28264 23848
rect 26375 23817 26387 23820
rect 26329 23811 26387 23817
rect 28258 23808 28264 23820
rect 28316 23808 28322 23860
rect 40586 23848 40592 23860
rect 40547 23820 40592 23848
rect 40586 23808 40592 23820
rect 40644 23808 40650 23860
rect 41325 23851 41383 23857
rect 41325 23817 41337 23851
rect 41371 23817 41383 23851
rect 41325 23811 41383 23817
rect 27709 23783 27767 23789
rect 27709 23749 27721 23783
rect 27755 23780 27767 23783
rect 28350 23780 28356 23792
rect 27755 23752 28356 23780
rect 27755 23749 27767 23752
rect 27709 23743 27767 23749
rect 28350 23740 28356 23752
rect 28408 23740 28414 23792
rect 37734 23712 37740 23724
rect 25363 23684 26188 23712
rect 37695 23684 37740 23712
rect 25363 23681 25375 23684
rect 25317 23675 25375 23681
rect 37734 23672 37740 23684
rect 37792 23672 37798 23724
rect 39206 23712 39212 23724
rect 39167 23684 39212 23712
rect 39206 23672 39212 23684
rect 39264 23672 39270 23724
rect 40221 23715 40279 23721
rect 40221 23681 40233 23715
rect 40267 23681 40279 23715
rect 41138 23712 41144 23724
rect 41099 23684 41144 23712
rect 40221 23675 40279 23681
rect 22152 23616 22324 23644
rect 22152 23604 22158 23616
rect 22370 23604 22376 23656
rect 22428 23644 22434 23656
rect 22465 23647 22523 23653
rect 22465 23644 22477 23647
rect 22428 23616 22477 23644
rect 22428 23604 22434 23616
rect 22465 23613 22477 23616
rect 22511 23644 22523 23647
rect 27525 23647 27583 23653
rect 22511 23616 25544 23644
rect 22511 23613 22523 23616
rect 22465 23607 22523 23613
rect 17604 23548 18184 23576
rect 14737 23539 14795 23545
rect 20070 23508 20076 23520
rect 12406 23480 20076 23508
rect 1995 23477 2007 23480
rect 1949 23471 2007 23477
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 23106 23508 23112 23520
rect 23067 23480 23112 23508
rect 23106 23468 23112 23480
rect 23164 23468 23170 23520
rect 25406 23508 25412 23520
rect 25367 23480 25412 23508
rect 25406 23468 25412 23480
rect 25464 23468 25470 23520
rect 25516 23508 25544 23616
rect 27525 23613 27537 23647
rect 27571 23644 27583 23647
rect 27798 23644 27804 23656
rect 27571 23616 27804 23644
rect 27571 23613 27583 23616
rect 27525 23607 27583 23613
rect 27798 23604 27804 23616
rect 27856 23604 27862 23656
rect 27985 23647 28043 23653
rect 27985 23613 27997 23647
rect 28031 23613 28043 23647
rect 27985 23607 28043 23613
rect 25590 23536 25596 23588
rect 25648 23576 25654 23588
rect 28000 23576 28028 23607
rect 38470 23604 38476 23656
rect 38528 23644 38534 23656
rect 39117 23647 39175 23653
rect 39117 23644 39129 23647
rect 38528 23616 39129 23644
rect 38528 23604 38534 23616
rect 39117 23613 39129 23616
rect 39163 23613 39175 23647
rect 39117 23607 39175 23613
rect 39577 23647 39635 23653
rect 39577 23613 39589 23647
rect 39623 23644 39635 23647
rect 40129 23647 40187 23653
rect 40129 23644 40141 23647
rect 39623 23616 40141 23644
rect 39623 23613 39635 23616
rect 39577 23607 39635 23613
rect 40129 23613 40141 23616
rect 40175 23613 40187 23647
rect 40236 23644 40264 23675
rect 41138 23672 41144 23684
rect 41196 23672 41202 23724
rect 41230 23672 41236 23724
rect 41288 23712 41294 23724
rect 41340 23712 41368 23811
rect 45370 23808 45376 23860
rect 45428 23848 45434 23860
rect 47673 23851 47731 23857
rect 47673 23848 47685 23851
rect 45428 23820 47685 23848
rect 45428 23808 45434 23820
rect 47673 23817 47685 23820
rect 47719 23817 47731 23851
rect 47673 23811 47731 23817
rect 42705 23783 42763 23789
rect 42705 23749 42717 23783
rect 42751 23780 42763 23783
rect 47486 23780 47492 23792
rect 42751 23752 47492 23780
rect 42751 23749 42763 23752
rect 42705 23743 42763 23749
rect 47486 23740 47492 23752
rect 47544 23740 47550 23792
rect 42429 23715 42487 23721
rect 42429 23712 42441 23715
rect 41288 23684 42441 23712
rect 41288 23672 41294 23684
rect 42429 23681 42441 23684
rect 42475 23681 42487 23715
rect 43346 23712 43352 23724
rect 43307 23684 43352 23712
rect 42429 23675 42487 23681
rect 43346 23672 43352 23684
rect 43404 23672 43410 23724
rect 43533 23715 43591 23721
rect 43533 23681 43545 23715
rect 43579 23712 43591 23715
rect 44818 23712 44824 23724
rect 43579 23684 44824 23712
rect 43579 23681 43591 23684
rect 43533 23675 43591 23681
rect 44818 23672 44824 23684
rect 44876 23672 44882 23724
rect 47581 23715 47639 23721
rect 47581 23681 47593 23715
rect 47627 23681 47639 23715
rect 47581 23675 47639 23681
rect 42518 23644 42524 23656
rect 40236 23616 42524 23644
rect 40129 23607 40187 23613
rect 42518 23604 42524 23616
rect 42576 23604 42582 23656
rect 45186 23644 45192 23656
rect 45147 23616 45192 23644
rect 45186 23604 45192 23616
rect 45244 23604 45250 23656
rect 45373 23647 45431 23653
rect 45373 23613 45385 23647
rect 45419 23644 45431 23647
rect 45646 23644 45652 23656
rect 45419 23616 45652 23644
rect 45419 23613 45431 23616
rect 45373 23607 45431 23613
rect 45646 23604 45652 23616
rect 45704 23604 45710 23656
rect 46658 23644 46664 23656
rect 46619 23616 46664 23644
rect 46658 23604 46664 23616
rect 46716 23604 46722 23656
rect 47394 23576 47400 23588
rect 25648 23548 28028 23576
rect 31726 23548 47400 23576
rect 25648 23536 25654 23548
rect 31726 23508 31754 23548
rect 47394 23536 47400 23548
rect 47452 23576 47458 23588
rect 47596 23576 47624 23675
rect 47452 23548 47624 23576
rect 47452 23536 47458 23548
rect 25516 23480 31754 23508
rect 38013 23511 38071 23517
rect 38013 23477 38025 23511
rect 38059 23508 38071 23511
rect 38562 23508 38568 23520
rect 38059 23480 38568 23508
rect 38059 23477 38071 23480
rect 38013 23471 38071 23477
rect 38562 23468 38568 23480
rect 38620 23468 38626 23520
rect 42978 23468 42984 23520
rect 43036 23508 43042 23520
rect 43441 23511 43499 23517
rect 43441 23508 43453 23511
rect 43036 23480 43453 23508
rect 43036 23468 43042 23480
rect 43441 23477 43453 23480
rect 43487 23477 43499 23511
rect 43441 23471 43499 23477
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 8570 23264 8576 23316
rect 8628 23304 8634 23316
rect 9033 23307 9091 23313
rect 9033 23304 9045 23307
rect 8628 23276 9045 23304
rect 8628 23264 8634 23276
rect 9033 23273 9045 23276
rect 9079 23273 9091 23307
rect 39482 23304 39488 23316
rect 9033 23267 9091 23273
rect 11716 23276 39488 23304
rect 2130 23196 2136 23248
rect 2188 23236 2194 23248
rect 11716 23236 11744 23276
rect 39482 23264 39488 23276
rect 39540 23264 39546 23316
rect 43162 23264 43168 23316
rect 43220 23304 43226 23316
rect 43441 23307 43499 23313
rect 43441 23304 43453 23307
rect 43220 23276 43453 23304
rect 43220 23264 43226 23276
rect 43441 23273 43453 23276
rect 43487 23273 43499 23307
rect 43441 23267 43499 23273
rect 43622 23264 43628 23316
rect 43680 23304 43686 23316
rect 47026 23304 47032 23316
rect 43680 23276 47032 23304
rect 43680 23264 43686 23276
rect 47026 23264 47032 23276
rect 47084 23264 47090 23316
rect 47762 23264 47768 23316
rect 47820 23304 47826 23316
rect 47946 23304 47952 23316
rect 47820 23276 47952 23304
rect 47820 23264 47826 23276
rect 47946 23264 47952 23276
rect 48004 23264 48010 23316
rect 17126 23236 17132 23248
rect 2188 23208 11744 23236
rect 16500 23208 17132 23236
rect 2188 23196 2194 23208
rect 13722 23128 13728 23180
rect 13780 23168 13786 23180
rect 16500 23177 16528 23208
rect 17126 23196 17132 23208
rect 17184 23196 17190 23248
rect 17865 23239 17923 23245
rect 17865 23205 17877 23239
rect 17911 23236 17923 23239
rect 18046 23236 18052 23248
rect 17911 23208 18052 23236
rect 17911 23205 17923 23208
rect 17865 23199 17923 23205
rect 18046 23196 18052 23208
rect 18104 23196 18110 23248
rect 20070 23236 20076 23248
rect 19983 23208 20076 23236
rect 20070 23196 20076 23208
rect 20128 23236 20134 23248
rect 20530 23236 20536 23248
rect 20128 23208 20536 23236
rect 20128 23196 20134 23208
rect 20530 23196 20536 23208
rect 20588 23196 20594 23248
rect 41138 23236 41144 23248
rect 37568 23208 41144 23236
rect 16485 23171 16543 23177
rect 13780 23140 15424 23168
rect 13780 23128 13786 23140
rect 8938 23100 8944 23112
rect 8899 23072 8944 23100
rect 8938 23060 8944 23072
rect 8996 23060 9002 23112
rect 10686 23100 10692 23112
rect 10647 23072 10692 23100
rect 10686 23060 10692 23072
rect 10744 23100 10750 23112
rect 11698 23100 11704 23112
rect 10744 23072 11704 23100
rect 10744 23060 10750 23072
rect 11698 23060 11704 23072
rect 11756 23060 11762 23112
rect 14734 23100 14740 23112
rect 14695 23072 14740 23100
rect 14734 23060 14740 23072
rect 14792 23060 14798 23112
rect 15396 23109 15424 23140
rect 16485 23137 16497 23171
rect 16531 23137 16543 23171
rect 16758 23168 16764 23180
rect 16719 23140 16764 23168
rect 16485 23131 16543 23137
rect 16758 23128 16764 23140
rect 16816 23128 16822 23180
rect 22738 23168 22744 23180
rect 20640 23140 22744 23168
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23069 15439 23103
rect 15381 23063 15439 23069
rect 16393 23103 16451 23109
rect 16393 23069 16405 23103
rect 16439 23100 16451 23103
rect 16574 23100 16580 23112
rect 16439 23072 16580 23100
rect 16439 23069 16451 23072
rect 16393 23063 16451 23069
rect 16574 23060 16580 23072
rect 16632 23060 16638 23112
rect 17681 23103 17739 23109
rect 17681 23069 17693 23103
rect 17727 23069 17739 23103
rect 19886 23100 19892 23112
rect 19847 23072 19892 23100
rect 17681 23063 17739 23069
rect 14752 23032 14780 23060
rect 17696 23032 17724 23063
rect 19886 23060 19892 23072
rect 19944 23060 19950 23112
rect 20640 23109 20668 23140
rect 22738 23128 22744 23140
rect 22796 23168 22802 23180
rect 23198 23168 23204 23180
rect 22796 23140 23204 23168
rect 22796 23128 22802 23140
rect 23198 23128 23204 23140
rect 23256 23128 23262 23180
rect 23477 23171 23535 23177
rect 23477 23137 23489 23171
rect 23523 23168 23535 23171
rect 25225 23171 25283 23177
rect 25225 23168 25237 23171
rect 23523 23140 25237 23168
rect 23523 23137 23535 23140
rect 23477 23131 23535 23137
rect 25225 23137 25237 23140
rect 25271 23137 25283 23171
rect 25406 23168 25412 23180
rect 25367 23140 25412 23168
rect 25225 23131 25283 23137
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23069 20683 23103
rect 21726 23100 21732 23112
rect 21687 23072 21732 23100
rect 20625 23063 20683 23069
rect 14752 23004 17724 23032
rect 17862 22992 17868 23044
rect 17920 23032 17926 23044
rect 20640 23032 20668 23063
rect 21726 23060 21732 23072
rect 21784 23060 21790 23112
rect 23106 23060 23112 23112
rect 23164 23060 23170 23112
rect 17920 23004 20668 23032
rect 22005 23035 22063 23041
rect 17920 22992 17926 23004
rect 22005 23001 22017 23035
rect 22051 23032 22063 23035
rect 22051 23004 22416 23032
rect 22051 23001 22063 23004
rect 22005 22995 22063 23001
rect 10873 22967 10931 22973
rect 10873 22933 10885 22967
rect 10919 22964 10931 22967
rect 11514 22964 11520 22976
rect 10919 22936 11520 22964
rect 10919 22933 10931 22936
rect 10873 22927 10931 22933
rect 11514 22924 11520 22936
rect 11572 22924 11578 22976
rect 14366 22924 14372 22976
rect 14424 22964 14430 22976
rect 14829 22967 14887 22973
rect 14829 22964 14841 22967
rect 14424 22936 14841 22964
rect 14424 22924 14430 22936
rect 14829 22933 14841 22936
rect 14875 22933 14887 22967
rect 14829 22927 14887 22933
rect 15378 22924 15384 22976
rect 15436 22964 15442 22976
rect 15473 22967 15531 22973
rect 15473 22964 15485 22967
rect 15436 22936 15485 22964
rect 15436 22924 15442 22936
rect 15473 22933 15485 22936
rect 15519 22933 15531 22967
rect 15473 22927 15531 22933
rect 20809 22967 20867 22973
rect 20809 22933 20821 22967
rect 20855 22964 20867 22967
rect 22094 22964 22100 22976
rect 20855 22936 22100 22964
rect 20855 22933 20867 22936
rect 20809 22927 20867 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 22388 22964 22416 23004
rect 22738 22964 22744 22976
rect 22388 22936 22744 22964
rect 22738 22924 22744 22936
rect 22796 22924 22802 22976
rect 22830 22924 22836 22976
rect 22888 22964 22894 22976
rect 23290 22964 23296 22976
rect 22888 22936 23296 22964
rect 22888 22924 22894 22936
rect 23290 22924 23296 22936
rect 23348 22964 23354 22976
rect 23492 22964 23520 23131
rect 25406 23128 25412 23140
rect 25464 23128 25470 23180
rect 25958 23128 25964 23180
rect 26016 23168 26022 23180
rect 26234 23168 26240 23180
rect 26016 23140 26240 23168
rect 26016 23128 26022 23140
rect 26234 23128 26240 23140
rect 26292 23128 26298 23180
rect 27890 23168 27896 23180
rect 27851 23140 27896 23168
rect 27890 23128 27896 23140
rect 27948 23128 27954 23180
rect 28074 23128 28080 23180
rect 28132 23168 28138 23180
rect 28169 23171 28227 23177
rect 28169 23168 28181 23171
rect 28132 23140 28181 23168
rect 28132 23128 28138 23140
rect 28169 23137 28181 23140
rect 28215 23137 28227 23171
rect 28169 23131 28227 23137
rect 27798 23100 27804 23112
rect 27711 23072 27804 23100
rect 27798 23060 27804 23072
rect 27856 23100 27862 23112
rect 28442 23100 28448 23112
rect 27856 23072 28448 23100
rect 27856 23060 27862 23072
rect 28442 23060 28448 23072
rect 28500 23060 28506 23112
rect 36446 23060 36452 23112
rect 36504 23100 36510 23112
rect 36817 23103 36875 23109
rect 36817 23100 36829 23103
rect 36504 23072 36829 23100
rect 36504 23060 36510 23072
rect 36817 23069 36829 23072
rect 36863 23100 36875 23103
rect 37568 23100 37596 23208
rect 41138 23196 41144 23208
rect 41196 23196 41202 23248
rect 42889 23239 42947 23245
rect 42889 23205 42901 23239
rect 42935 23236 42947 23239
rect 45186 23236 45192 23248
rect 42935 23208 45192 23236
rect 42935 23205 42947 23208
rect 42889 23199 42947 23205
rect 45186 23196 45192 23208
rect 45244 23236 45250 23248
rect 45244 23208 45416 23236
rect 45244 23196 45250 23208
rect 38378 23168 38384 23180
rect 38291 23140 38384 23168
rect 38378 23128 38384 23140
rect 38436 23168 38442 23180
rect 38930 23168 38936 23180
rect 38436 23140 38936 23168
rect 38436 23128 38442 23140
rect 38930 23128 38936 23140
rect 38988 23128 38994 23180
rect 40037 23171 40095 23177
rect 40037 23137 40049 23171
rect 40083 23168 40095 23171
rect 40586 23168 40592 23180
rect 40083 23140 40592 23168
rect 40083 23137 40095 23140
rect 40037 23131 40095 23137
rect 40586 23128 40592 23140
rect 40644 23128 40650 23180
rect 43346 23128 43352 23180
rect 43404 23168 43410 23180
rect 45388 23177 45416 23208
rect 45373 23171 45431 23177
rect 43404 23140 44036 23168
rect 43404 23128 43410 23140
rect 37734 23100 37740 23112
rect 36863 23072 37596 23100
rect 37695 23072 37740 23100
rect 36863 23069 36875 23072
rect 36817 23063 36875 23069
rect 37734 23060 37740 23072
rect 37792 23060 37798 23112
rect 42794 23060 42800 23112
rect 42852 23100 42858 23112
rect 44008 23109 44036 23140
rect 45373 23137 45385 23171
rect 45419 23137 45431 23171
rect 45373 23131 45431 23137
rect 43014 23103 43072 23109
rect 43014 23100 43026 23103
rect 42852 23072 43026 23100
rect 42852 23060 42858 23072
rect 43014 23069 43026 23072
rect 43060 23069 43072 23103
rect 43014 23063 43072 23069
rect 43533 23103 43591 23109
rect 43533 23069 43545 23103
rect 43579 23069 43591 23103
rect 43533 23063 43591 23069
rect 43993 23103 44051 23109
rect 43993 23069 44005 23103
rect 44039 23069 44051 23103
rect 43993 23063 44051 23069
rect 44177 23103 44235 23109
rect 44177 23069 44189 23103
rect 44223 23100 44235 23103
rect 44818 23100 44824 23112
rect 44223 23072 44824 23100
rect 44223 23069 44235 23072
rect 44177 23063 44235 23069
rect 27065 23035 27123 23041
rect 27065 23001 27077 23035
rect 27111 23032 27123 23035
rect 40034 23032 40040 23044
rect 27111 23004 40040 23032
rect 27111 23001 27123 23004
rect 27065 22995 27123 23001
rect 40034 22992 40040 23004
rect 40092 22992 40098 23044
rect 40221 23035 40279 23041
rect 40221 23001 40233 23035
rect 40267 23032 40279 23035
rect 40770 23032 40776 23044
rect 40267 23004 40776 23032
rect 40267 23001 40279 23004
rect 40221 22995 40279 23001
rect 40770 22992 40776 23004
rect 40828 22992 40834 23044
rect 41782 22992 41788 23044
rect 41840 23032 41846 23044
rect 41877 23035 41935 23041
rect 41877 23032 41889 23035
rect 41840 23004 41889 23032
rect 41840 22992 41846 23004
rect 41877 23001 41889 23004
rect 41923 23001 41935 23035
rect 41877 22995 41935 23001
rect 42518 22992 42524 23044
rect 42576 23032 42582 23044
rect 43548 23032 43576 23063
rect 44818 23060 44824 23072
rect 44876 23060 44882 23112
rect 47673 23103 47731 23109
rect 47673 23069 47685 23103
rect 47719 23100 47731 23103
rect 48130 23100 48136 23112
rect 47719 23072 48136 23100
rect 47719 23069 47731 23072
rect 47673 23063 47731 23069
rect 48130 23060 48136 23072
rect 48188 23060 48194 23112
rect 42576 23004 43576 23032
rect 42576 22992 42582 23004
rect 44266 22992 44272 23044
rect 44324 23032 44330 23044
rect 45557 23035 45615 23041
rect 45557 23032 45569 23035
rect 44324 23004 45569 23032
rect 44324 22992 44330 23004
rect 45557 23001 45569 23004
rect 45603 23001 45615 23035
rect 47210 23032 47216 23044
rect 47171 23004 47216 23032
rect 45557 22995 45615 23001
rect 47210 22992 47216 23004
rect 47268 22992 47274 23044
rect 23348 22936 23520 22964
rect 37001 22967 37059 22973
rect 23348 22924 23354 22936
rect 37001 22933 37013 22967
rect 37047 22964 37059 22967
rect 37734 22964 37740 22976
rect 37047 22936 37740 22964
rect 37047 22933 37059 22936
rect 37001 22927 37059 22933
rect 37734 22924 37740 22936
rect 37792 22924 37798 22976
rect 43073 22967 43131 22973
rect 43073 22933 43085 22967
rect 43119 22964 43131 22967
rect 43162 22964 43168 22976
rect 43119 22936 43168 22964
rect 43119 22933 43131 22936
rect 43073 22927 43131 22933
rect 43162 22924 43168 22936
rect 43220 22964 43226 22976
rect 44085 22967 44143 22973
rect 44085 22964 44097 22967
rect 43220 22936 44097 22964
rect 43220 22924 43226 22936
rect 44085 22933 44097 22936
rect 44131 22933 44143 22967
rect 44085 22927 44143 22933
rect 45094 22924 45100 22976
rect 45152 22964 45158 22976
rect 48133 22967 48191 22973
rect 48133 22964 48145 22967
rect 45152 22936 48145 22964
rect 45152 22924 45158 22936
rect 48133 22933 48145 22936
rect 48179 22933 48191 22967
rect 48133 22927 48191 22933
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 12710 22720 12716 22772
rect 12768 22760 12774 22772
rect 16758 22760 16764 22772
rect 12768 22732 13584 22760
rect 12768 22720 12774 22732
rect 3878 22652 3884 22704
rect 3936 22692 3942 22704
rect 12066 22692 12072 22704
rect 3936 22664 6914 22692
rect 3936 22652 3942 22664
rect 6886 22488 6914 22664
rect 8496 22664 12072 22692
rect 8496 22633 8524 22664
rect 12066 22652 12072 22664
rect 12124 22652 12130 22704
rect 12434 22652 12440 22704
rect 12492 22652 12498 22704
rect 13556 22701 13584 22732
rect 14660 22732 16764 22760
rect 14660 22701 14688 22732
rect 16758 22720 16764 22732
rect 16816 22720 16822 22772
rect 22112 22732 22600 22760
rect 13541 22695 13599 22701
rect 13541 22661 13553 22695
rect 13587 22661 13599 22695
rect 13541 22655 13599 22661
rect 14645 22695 14703 22701
rect 14645 22661 14657 22695
rect 14691 22661 14703 22695
rect 14645 22655 14703 22661
rect 15378 22652 15384 22704
rect 15436 22652 15442 22704
rect 22112 22701 22140 22732
rect 22087 22695 22145 22701
rect 22087 22661 22099 22695
rect 22133 22661 22145 22695
rect 22572 22692 22600 22732
rect 22738 22720 22744 22772
rect 22796 22760 22802 22772
rect 23753 22763 23811 22769
rect 23753 22760 23765 22763
rect 22796 22732 23765 22760
rect 22796 22720 22802 22732
rect 23753 22729 23765 22732
rect 23799 22729 23811 22763
rect 26234 22760 26240 22772
rect 26147 22732 26240 22760
rect 23753 22723 23811 22729
rect 26234 22720 26240 22732
rect 26292 22760 26298 22772
rect 27154 22760 27160 22772
rect 26292 22732 27160 22760
rect 26292 22720 26298 22732
rect 27154 22720 27160 22732
rect 27212 22720 27218 22772
rect 28442 22720 28448 22772
rect 28500 22760 28506 22772
rect 29273 22763 29331 22769
rect 29273 22760 29285 22763
rect 28500 22732 29285 22760
rect 28500 22720 28506 22732
rect 29273 22729 29285 22732
rect 29319 22729 29331 22763
rect 37734 22760 37740 22772
rect 29273 22723 29331 22729
rect 35820 22732 37740 22760
rect 22830 22692 22836 22704
rect 22572 22664 22836 22692
rect 22087 22655 22145 22661
rect 22830 22652 22836 22664
rect 22888 22652 22894 22704
rect 23063 22661 23121 22667
rect 23063 22658 23075 22661
rect 8481 22627 8539 22633
rect 8481 22593 8493 22627
rect 8527 22593 8539 22627
rect 11514 22624 11520 22636
rect 11475 22596 11520 22624
rect 8481 22587 8539 22593
rect 11514 22584 11520 22596
rect 11572 22584 11578 22636
rect 14366 22624 14372 22636
rect 14327 22596 14372 22624
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 21450 22584 21456 22636
rect 21508 22624 21514 22636
rect 22281 22630 22339 22633
rect 22204 22627 22339 22630
rect 22204 22624 22293 22627
rect 21508 22602 22293 22624
rect 21508 22596 22232 22602
rect 21508 22584 21514 22596
rect 8662 22556 8668 22568
rect 8623 22528 8668 22556
rect 8662 22516 8668 22528
rect 8720 22516 8726 22568
rect 8941 22559 8999 22565
rect 8941 22525 8953 22559
rect 8987 22525 8999 22559
rect 11790 22556 11796 22568
rect 11751 22528 11796 22556
rect 8941 22519 8999 22525
rect 8956 22488 8984 22519
rect 11790 22516 11796 22528
rect 11848 22516 11854 22568
rect 16117 22559 16175 22565
rect 16117 22525 16129 22559
rect 16163 22556 16175 22559
rect 16574 22556 16580 22568
rect 16163 22528 16580 22556
rect 16163 22525 16175 22528
rect 16117 22519 16175 22525
rect 16574 22516 16580 22528
rect 16632 22556 16638 22568
rect 17589 22559 17647 22565
rect 17589 22556 17601 22559
rect 16632 22528 17601 22556
rect 16632 22516 16638 22528
rect 17589 22525 17601 22528
rect 17635 22525 17647 22559
rect 17770 22556 17776 22568
rect 17731 22528 17776 22556
rect 17589 22519 17647 22525
rect 17770 22516 17776 22528
rect 17828 22516 17834 22568
rect 19058 22556 19064 22568
rect 19019 22528 19064 22556
rect 19058 22516 19064 22528
rect 19116 22516 19122 22568
rect 6886 22460 8984 22488
rect 22020 22420 22048 22596
rect 22281 22593 22293 22602
rect 22327 22593 22339 22627
rect 22281 22587 22339 22593
rect 22373 22627 22431 22633
rect 22373 22593 22385 22627
rect 22419 22624 22431 22627
rect 22462 22624 22468 22636
rect 22419 22596 22468 22624
rect 22419 22593 22431 22596
rect 22373 22587 22431 22593
rect 22462 22584 22468 22596
rect 22520 22624 22526 22636
rect 23048 22627 23075 22658
rect 23109 22627 23121 22661
rect 25774 22652 25780 22704
rect 25832 22652 25838 22704
rect 27801 22695 27859 22701
rect 27801 22661 27813 22695
rect 27847 22692 27859 22695
rect 28074 22692 28080 22704
rect 27847 22664 28080 22692
rect 27847 22661 27859 22664
rect 27801 22655 27859 22661
rect 28074 22652 28080 22664
rect 28132 22652 28138 22704
rect 28810 22652 28816 22704
rect 28868 22652 28874 22704
rect 23048 22624 23121 22627
rect 23566 22624 23572 22636
rect 22520 22596 23572 22624
rect 22520 22584 22526 22596
rect 23566 22584 23572 22596
rect 23624 22584 23630 22636
rect 23661 22627 23719 22633
rect 23661 22593 23673 22627
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 23845 22627 23903 22633
rect 23845 22593 23857 22627
rect 23891 22593 23903 22627
rect 34698 22624 34704 22636
rect 34659 22596 34704 22624
rect 23845 22587 23903 22593
rect 23676 22556 23704 22587
rect 22572 22528 23704 22556
rect 22097 22491 22155 22497
rect 22097 22457 22109 22491
rect 22143 22488 22155 22491
rect 22186 22488 22192 22500
rect 22143 22460 22192 22488
rect 22143 22457 22155 22460
rect 22097 22451 22155 22457
rect 22186 22448 22192 22460
rect 22244 22448 22250 22500
rect 22278 22448 22284 22500
rect 22336 22488 22342 22500
rect 22572 22488 22600 22528
rect 22336 22460 22600 22488
rect 22336 22448 22342 22460
rect 22646 22448 22652 22500
rect 22704 22488 22710 22500
rect 23201 22491 23259 22497
rect 23201 22488 23213 22491
rect 22704 22460 23213 22488
rect 22704 22448 22710 22460
rect 23201 22457 23213 22460
rect 23247 22488 23259 22491
rect 23860 22488 23888 22587
rect 34698 22584 34704 22596
rect 34756 22584 34762 22636
rect 35820 22633 35848 22732
rect 37734 22720 37740 22732
rect 37792 22720 37798 22772
rect 39482 22760 39488 22772
rect 39443 22732 39488 22760
rect 39482 22720 39488 22732
rect 39540 22720 39546 22772
rect 40770 22760 40776 22772
rect 40731 22732 40776 22760
rect 40770 22720 40776 22732
rect 40828 22720 40834 22772
rect 42518 22720 42524 22772
rect 42576 22760 42582 22772
rect 42797 22763 42855 22769
rect 42797 22760 42809 22763
rect 42576 22732 42809 22760
rect 42576 22720 42582 22732
rect 42797 22729 42809 22732
rect 42843 22729 42855 22763
rect 44266 22760 44272 22772
rect 44227 22732 44272 22760
rect 42797 22723 42855 22729
rect 44266 22720 44272 22732
rect 44324 22720 44330 22772
rect 45646 22760 45652 22772
rect 45607 22732 45652 22760
rect 45646 22720 45652 22732
rect 45704 22720 45710 22772
rect 35897 22695 35955 22701
rect 35897 22661 35909 22695
rect 35943 22692 35955 22695
rect 37553 22695 37611 22701
rect 37553 22692 37565 22695
rect 35943 22664 37565 22692
rect 35943 22661 35955 22664
rect 35897 22655 35955 22661
rect 37553 22661 37565 22664
rect 37599 22661 37611 22695
rect 37553 22655 37611 22661
rect 39209 22695 39267 22701
rect 39209 22661 39221 22695
rect 39255 22692 39267 22695
rect 45738 22692 45744 22704
rect 39255 22664 45744 22692
rect 39255 22661 39267 22664
rect 39209 22655 39267 22661
rect 45738 22652 45744 22664
rect 45796 22652 45802 22704
rect 35805 22627 35863 22633
rect 35805 22593 35817 22627
rect 35851 22593 35863 22627
rect 36446 22624 36452 22636
rect 36407 22596 36452 22624
rect 35805 22587 35863 22593
rect 36446 22584 36452 22596
rect 36504 22584 36510 22636
rect 39758 22584 39764 22636
rect 39816 22624 39822 22636
rect 39853 22627 39911 22633
rect 39853 22624 39865 22627
rect 39816 22596 39865 22624
rect 39816 22584 39822 22596
rect 39853 22593 39865 22596
rect 39899 22593 39911 22627
rect 40957 22627 41015 22633
rect 40957 22624 40969 22627
rect 39853 22587 39911 22593
rect 40328 22596 40969 22624
rect 24486 22556 24492 22568
rect 24447 22528 24492 22556
rect 24486 22516 24492 22528
rect 24544 22516 24550 22568
rect 24762 22556 24768 22568
rect 24723 22528 24768 22556
rect 24762 22516 24768 22528
rect 24820 22516 24826 22568
rect 27522 22556 27528 22568
rect 27483 22528 27528 22556
rect 27522 22516 27528 22528
rect 27580 22516 27586 22568
rect 40328 22565 40356 22596
rect 40957 22593 40969 22596
rect 41003 22593 41015 22627
rect 42978 22624 42984 22636
rect 42939 22596 42984 22624
rect 40957 22587 41015 22593
rect 42978 22584 42984 22596
rect 43036 22584 43042 22636
rect 43162 22624 43168 22636
rect 43123 22596 43168 22624
rect 43162 22584 43168 22596
rect 43220 22584 43226 22636
rect 44453 22627 44511 22633
rect 44453 22593 44465 22627
rect 44499 22593 44511 22627
rect 45094 22624 45100 22636
rect 45055 22596 45100 22624
rect 44453 22587 44511 22593
rect 37369 22559 37427 22565
rect 37369 22556 37381 22559
rect 28920 22528 37381 22556
rect 28920 22500 28948 22528
rect 37369 22525 37381 22528
rect 37415 22525 37427 22559
rect 37369 22519 37427 22525
rect 40313 22559 40371 22565
rect 40313 22525 40325 22559
rect 40359 22525 40371 22559
rect 40313 22519 40371 22525
rect 42794 22516 42800 22568
rect 42852 22556 42858 22568
rect 43257 22559 43315 22565
rect 43257 22556 43269 22559
rect 42852 22528 43269 22556
rect 42852 22516 42858 22528
rect 43257 22525 43269 22528
rect 43303 22525 43315 22559
rect 43257 22519 43315 22525
rect 23247 22460 23888 22488
rect 23247 22457 23259 22460
rect 23201 22451 23259 22457
rect 28902 22448 28908 22500
rect 28960 22448 28966 22500
rect 44468 22488 44496 22587
rect 45094 22584 45100 22596
rect 45152 22584 45158 22636
rect 45554 22624 45560 22636
rect 45515 22596 45560 22624
rect 45554 22584 45560 22596
rect 45612 22584 45618 22636
rect 47578 22624 47584 22636
rect 47539 22596 47584 22624
rect 47578 22584 47584 22596
rect 47636 22584 47642 22636
rect 46198 22556 46204 22568
rect 46159 22528 46204 22556
rect 46198 22516 46204 22528
rect 46256 22516 46262 22568
rect 46474 22556 46480 22568
rect 46435 22528 46480 22556
rect 46474 22516 46480 22528
rect 46532 22516 46538 22568
rect 47854 22556 47860 22568
rect 47815 22528 47860 22556
rect 47854 22516 47860 22528
rect 47912 22516 47918 22568
rect 48133 22491 48191 22497
rect 48133 22488 48145 22491
rect 44468 22460 48145 22488
rect 48133 22457 48145 22460
rect 48179 22457 48191 22491
rect 48133 22451 48191 22457
rect 23017 22423 23075 22429
rect 23017 22420 23029 22423
rect 22020 22392 23029 22420
rect 23017 22389 23029 22392
rect 23063 22420 23075 22423
rect 23474 22420 23480 22432
rect 23063 22392 23480 22420
rect 23063 22389 23075 22392
rect 23017 22383 23075 22389
rect 23474 22380 23480 22392
rect 23532 22380 23538 22432
rect 34514 22420 34520 22432
rect 34475 22392 34520 22420
rect 34514 22380 34520 22392
rect 34572 22380 34578 22432
rect 36630 22420 36636 22432
rect 36591 22392 36636 22420
rect 36630 22380 36636 22392
rect 36688 22380 36694 22432
rect 39482 22380 39488 22432
rect 39540 22420 39546 22432
rect 39945 22423 40003 22429
rect 39945 22420 39957 22423
rect 39540 22392 39957 22420
rect 39540 22380 39546 22392
rect 39945 22389 39957 22392
rect 39991 22420 40003 22423
rect 40034 22420 40040 22432
rect 39991 22392 40040 22420
rect 39991 22389 40003 22392
rect 39945 22383 40003 22389
rect 40034 22380 40040 22392
rect 40092 22380 40098 22432
rect 44913 22423 44971 22429
rect 44913 22389 44925 22423
rect 44959 22420 44971 22423
rect 45922 22420 45928 22432
rect 44959 22392 45928 22420
rect 44959 22389 44971 22392
rect 44913 22383 44971 22389
rect 45922 22380 45928 22392
rect 45980 22380 45986 22432
rect 46658 22380 46664 22432
rect 46716 22420 46722 22432
rect 47673 22423 47731 22429
rect 47673 22420 47685 22423
rect 46716 22392 47685 22420
rect 46716 22380 46722 22392
rect 47673 22389 47685 22392
rect 47719 22389 47731 22423
rect 47673 22383 47731 22389
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 8662 22176 8668 22228
rect 8720 22216 8726 22228
rect 9033 22219 9091 22225
rect 9033 22216 9045 22219
rect 8720 22188 9045 22216
rect 8720 22176 8726 22188
rect 9033 22185 9045 22188
rect 9079 22185 9091 22219
rect 9033 22179 9091 22185
rect 13170 22176 13176 22228
rect 13228 22216 13234 22228
rect 14274 22216 14280 22228
rect 13228 22188 14280 22216
rect 13228 22176 13234 22188
rect 14274 22176 14280 22188
rect 14332 22216 14338 22228
rect 14458 22216 14464 22228
rect 14332 22188 14464 22216
rect 14332 22176 14338 22188
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 17770 22216 17776 22228
rect 17731 22188 17776 22216
rect 17770 22176 17776 22188
rect 17828 22176 17834 22228
rect 19978 22176 19984 22228
rect 20036 22176 20042 22228
rect 21726 22176 21732 22228
rect 21784 22216 21790 22228
rect 21821 22219 21879 22225
rect 21821 22216 21833 22219
rect 21784 22188 21833 22216
rect 21784 22176 21790 22188
rect 21821 22185 21833 22188
rect 21867 22185 21879 22219
rect 21821 22179 21879 22185
rect 22373 22219 22431 22225
rect 22373 22185 22385 22219
rect 22419 22216 22431 22219
rect 23934 22216 23940 22228
rect 22419 22188 23940 22216
rect 22419 22185 22431 22188
rect 22373 22179 22431 22185
rect 23934 22176 23940 22188
rect 23992 22176 23998 22228
rect 24486 22216 24492 22228
rect 24447 22188 24492 22216
rect 24486 22176 24492 22188
rect 24544 22176 24550 22228
rect 27249 22219 27307 22225
rect 27249 22185 27261 22219
rect 27295 22216 27307 22219
rect 27522 22216 27528 22228
rect 27295 22188 27528 22216
rect 27295 22185 27307 22188
rect 27249 22179 27307 22185
rect 27522 22176 27528 22188
rect 27580 22176 27586 22228
rect 34698 22216 34704 22228
rect 34659 22188 34704 22216
rect 34698 22176 34704 22188
rect 34756 22176 34762 22228
rect 34790 22176 34796 22228
rect 34848 22216 34854 22228
rect 34885 22219 34943 22225
rect 34885 22216 34897 22219
rect 34848 22188 34897 22216
rect 34848 22176 34854 22188
rect 34885 22185 34897 22188
rect 34931 22216 34943 22219
rect 35437 22219 35495 22225
rect 35437 22216 35449 22219
rect 34931 22188 35449 22216
rect 34931 22185 34943 22188
rect 34885 22179 34943 22185
rect 35437 22185 35449 22188
rect 35483 22185 35495 22219
rect 35437 22179 35495 22185
rect 45186 22176 45192 22228
rect 45244 22216 45250 22228
rect 48130 22216 48136 22228
rect 45244 22188 48136 22216
rect 45244 22176 45250 22188
rect 48130 22176 48136 22188
rect 48188 22176 48194 22228
rect 10612 22120 10916 22148
rect 10612 22080 10640 22120
rect 10520 22052 10640 22080
rect 10689 22083 10747 22089
rect 8938 22012 8944 22024
rect 8851 21984 8944 22012
rect 8938 21972 8944 21984
rect 8996 22012 9002 22024
rect 10520 22012 10548 22052
rect 10689 22049 10701 22083
rect 10735 22080 10747 22083
rect 10778 22080 10784 22092
rect 10735 22052 10784 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 10778 22040 10784 22052
rect 10836 22040 10842 22092
rect 8996 21984 10548 22012
rect 10597 22015 10655 22021
rect 8996 21972 9002 21984
rect 10597 21981 10609 22015
rect 10643 22014 10655 22015
rect 10643 21986 10732 22014
rect 10643 21981 10655 21986
rect 10597 21975 10655 21981
rect 10704 21944 10732 21986
rect 10888 22012 10916 22120
rect 11992 22120 12572 22148
rect 10965 22083 11023 22089
rect 10965 22049 10977 22083
rect 11011 22080 11023 22083
rect 11790 22080 11796 22092
rect 11011 22052 11796 22080
rect 11011 22049 11023 22052
rect 10965 22043 11023 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 11992 22080 12020 22120
rect 11900 22052 12020 22080
rect 12069 22083 12127 22089
rect 11900 22012 11928 22052
rect 12069 22049 12081 22083
rect 12115 22080 12127 22083
rect 12434 22080 12440 22092
rect 12115 22052 12440 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 12434 22040 12440 22052
rect 12492 22040 12498 22092
rect 12544 22080 12572 22120
rect 13924 22120 14320 22148
rect 13722 22080 13728 22092
rect 12544 22052 13728 22080
rect 13722 22040 13728 22052
rect 13780 22040 13786 22092
rect 10888 21984 11928 22012
rect 11977 22015 12035 22021
rect 11977 21981 11989 22015
rect 12023 22012 12035 22015
rect 12250 22012 12256 22024
rect 12023 21984 12256 22012
rect 12023 21981 12035 21984
rect 11977 21975 12035 21981
rect 12250 21972 12256 21984
rect 12308 21972 12314 22024
rect 12621 22015 12679 22021
rect 12621 21981 12633 22015
rect 12667 22012 12679 22015
rect 13170 22012 13176 22024
rect 12667 21984 13176 22012
rect 12667 21981 12679 21984
rect 12621 21975 12679 21981
rect 13170 21972 13176 21984
rect 13228 21972 13234 22024
rect 13262 21972 13268 22024
rect 13320 22012 13326 22024
rect 13924 22012 13952 22120
rect 13998 22040 14004 22092
rect 14056 22080 14062 22092
rect 14098 22083 14156 22089
rect 14098 22080 14110 22083
rect 14056 22052 14110 22080
rect 14056 22040 14062 22052
rect 14098 22049 14110 22052
rect 14144 22049 14156 22083
rect 14292 22080 14320 22120
rect 14366 22108 14372 22160
rect 14424 22148 14430 22160
rect 17862 22148 17868 22160
rect 14424 22120 17868 22148
rect 14424 22108 14430 22120
rect 17862 22108 17868 22120
rect 17920 22108 17926 22160
rect 19996 22148 20024 22176
rect 43070 22148 43076 22160
rect 19536 22120 20024 22148
rect 22480 22120 23428 22148
rect 19242 22080 19248 22092
rect 14292 22052 19248 22080
rect 14098 22043 14156 22049
rect 19242 22040 19248 22052
rect 19300 22040 19306 22092
rect 19536 22089 19564 22120
rect 19521 22083 19579 22089
rect 19521 22049 19533 22083
rect 19567 22049 19579 22083
rect 19521 22043 19579 22049
rect 19797 22083 19855 22089
rect 19797 22049 19809 22083
rect 19843 22080 19855 22083
rect 19978 22080 19984 22092
rect 19843 22052 19984 22080
rect 19843 22049 19855 22052
rect 19797 22043 19855 22049
rect 19978 22040 19984 22052
rect 20036 22040 20042 22092
rect 22480 22080 22508 22120
rect 20456 22052 22508 22080
rect 23400 22080 23428 22120
rect 25516 22120 25912 22148
rect 43031 22120 43076 22148
rect 25516 22080 25544 22120
rect 25884 22092 25912 22120
rect 43070 22108 43076 22120
rect 43128 22108 43134 22160
rect 45922 22108 45928 22160
rect 45980 22148 45986 22160
rect 45980 22120 46060 22148
rect 45980 22108 45986 22120
rect 23400 22052 25544 22080
rect 25593 22083 25651 22089
rect 20456 22024 20484 22052
rect 16390 22012 16396 22024
rect 13320 21984 13952 22012
rect 16351 21984 16396 22012
rect 13320 21972 13326 21984
rect 16390 21972 16396 21984
rect 16448 21972 16454 22024
rect 17678 22012 17684 22024
rect 17639 21984 17684 22012
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 19334 21972 19340 22024
rect 19392 22012 19398 22024
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 19392 21984 19441 22012
rect 19392 21972 19398 21984
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 20438 22012 20444 22024
rect 20399 21984 20444 22012
rect 19429 21975 19487 21981
rect 20438 21972 20444 21984
rect 20496 21972 20502 22024
rect 21652 22021 21680 22052
rect 20993 22015 21051 22021
rect 20993 21981 21005 22015
rect 21039 21981 21051 22015
rect 20993 21975 21051 21981
rect 21637 22015 21695 22021
rect 21637 21981 21649 22015
rect 21683 21981 21695 22015
rect 21637 21975 21695 21981
rect 12526 21944 12532 21956
rect 10704 21916 12532 21944
rect 12526 21904 12532 21916
rect 12584 21904 12590 21956
rect 12713 21947 12771 21953
rect 12713 21913 12725 21947
rect 12759 21944 12771 21947
rect 14277 21947 14335 21953
rect 14277 21944 14289 21947
rect 12759 21916 14289 21944
rect 12759 21913 12771 21916
rect 12713 21907 12771 21913
rect 14277 21913 14289 21916
rect 14323 21913 14335 21947
rect 15930 21944 15936 21956
rect 15891 21916 15936 21944
rect 14277 21907 14335 21913
rect 15930 21904 15936 21916
rect 15988 21904 15994 21956
rect 17696 21944 17724 21972
rect 20070 21944 20076 21956
rect 17696 21916 20076 21944
rect 20070 21904 20076 21916
rect 20128 21904 20134 21956
rect 21008 21944 21036 21975
rect 22002 21972 22008 22024
rect 22060 22012 22066 22024
rect 22646 22012 22652 22024
rect 22060 21984 22508 22012
rect 22607 21984 22652 22012
rect 22060 21972 22066 21984
rect 22094 21944 22100 21956
rect 21008 21916 22100 21944
rect 22094 21904 22100 21916
rect 22152 21944 22158 21956
rect 22278 21944 22284 21956
rect 22152 21916 22284 21944
rect 22152 21904 22158 21916
rect 22278 21904 22284 21916
rect 22336 21904 22342 21956
rect 22373 21947 22431 21953
rect 22373 21913 22385 21947
rect 22419 21913 22431 21947
rect 22480 21944 22508 21984
rect 22646 21972 22652 21984
rect 22704 21972 22710 22024
rect 23106 22012 23112 22024
rect 23067 21984 23112 22012
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 23474 22012 23480 22024
rect 23435 21984 23480 22012
rect 23474 21972 23480 21984
rect 23532 21972 23538 22024
rect 24504 22021 24532 22052
rect 25593 22049 25605 22083
rect 25639 22080 25651 22083
rect 25774 22080 25780 22092
rect 25639 22052 25780 22080
rect 25639 22049 25651 22052
rect 25593 22043 25651 22049
rect 25774 22040 25780 22052
rect 25832 22040 25838 22092
rect 25866 22040 25872 22092
rect 25924 22040 25930 22092
rect 28828 22080 28948 22094
rect 46032 22089 46060 22120
rect 34057 22083 34115 22089
rect 25976 22066 34008 22080
rect 25976 22052 28856 22066
rect 28920 22052 34008 22066
rect 24489 22015 24547 22021
rect 24489 21981 24501 22015
rect 24535 21981 24547 22015
rect 24489 21975 24547 21981
rect 24670 21972 24676 22024
rect 24728 22012 24734 22024
rect 25498 22012 25504 22024
rect 24728 21984 25504 22012
rect 24728 21972 24734 21984
rect 25498 21972 25504 21984
rect 25556 21972 25562 22024
rect 25976 22012 26004 22052
rect 25608 21984 26004 22012
rect 22480 21916 22600 21944
rect 22373 21907 22431 21913
rect 11514 21836 11520 21888
rect 11572 21876 11578 21888
rect 13262 21876 13268 21888
rect 11572 21848 13268 21876
rect 11572 21836 11578 21848
rect 13262 21836 13268 21848
rect 13320 21836 13326 21888
rect 13449 21879 13507 21885
rect 13449 21845 13461 21879
rect 13495 21876 13507 21879
rect 14642 21876 14648 21888
rect 13495 21848 14648 21876
rect 13495 21845 13507 21848
rect 13449 21839 13507 21845
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 16574 21876 16580 21888
rect 16535 21848 16580 21876
rect 16574 21836 16580 21848
rect 16632 21876 16638 21888
rect 17034 21876 17040 21888
rect 16632 21848 17040 21876
rect 16632 21836 16638 21848
rect 17034 21836 17040 21848
rect 17092 21836 17098 21888
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 20441 21879 20499 21885
rect 20441 21876 20453 21879
rect 19484 21848 20453 21876
rect 19484 21836 19490 21848
rect 20441 21845 20453 21848
rect 20487 21845 20499 21879
rect 21082 21876 21088 21888
rect 21043 21848 21088 21876
rect 20441 21839 20499 21845
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 22388 21876 22416 21907
rect 22462 21876 22468 21888
rect 22388 21848 22468 21876
rect 22462 21836 22468 21848
rect 22520 21836 22526 21888
rect 22572 21885 22600 21916
rect 24302 21904 24308 21956
rect 24360 21944 24366 21956
rect 25608 21944 25636 21984
rect 26970 21972 26976 22024
rect 27028 22012 27034 22024
rect 27157 22015 27215 22021
rect 27157 22012 27169 22015
rect 27028 21984 27169 22012
rect 27028 21972 27034 21984
rect 27157 21981 27169 21984
rect 27203 21981 27215 22015
rect 27157 21975 27215 21981
rect 27798 21972 27804 22024
rect 27856 22012 27862 22024
rect 28721 22015 28779 22021
rect 28721 22012 28733 22015
rect 27856 21984 28733 22012
rect 27856 21972 27862 21984
rect 28721 21981 28733 21984
rect 28767 22012 28779 22015
rect 29362 22012 29368 22024
rect 28767 22006 28856 22012
rect 28920 22006 29368 22012
rect 28767 21984 29368 22006
rect 28767 21981 28779 21984
rect 28721 21975 28779 21981
rect 28828 21978 28948 21984
rect 29362 21972 29368 21984
rect 29420 21972 29426 22024
rect 29549 22015 29607 22021
rect 29549 22012 29561 22015
rect 29472 21984 29561 22012
rect 24360 21916 25636 21944
rect 24360 21904 24366 21916
rect 25866 21904 25872 21956
rect 25924 21944 25930 21956
rect 29472 21944 29500 21984
rect 29549 21981 29561 21984
rect 29595 21981 29607 22015
rect 29549 21975 29607 21981
rect 29730 21972 29736 22024
rect 29788 22012 29794 22024
rect 30285 22015 30343 22021
rect 30285 22012 30297 22015
rect 29788 21984 30297 22012
rect 29788 21972 29794 21984
rect 30285 21981 30297 21984
rect 30331 21981 30343 22015
rect 30285 21975 30343 21981
rect 31202 21972 31208 22024
rect 31260 22012 31266 22024
rect 32217 22015 32275 22021
rect 32217 22012 32229 22015
rect 31260 21984 32229 22012
rect 31260 21972 31266 21984
rect 32217 21981 32229 21984
rect 32263 21981 32275 22015
rect 32217 21975 32275 21981
rect 32398 21944 32404 21956
rect 25924 21916 29500 21944
rect 32359 21916 32404 21944
rect 25924 21904 25930 21916
rect 32398 21904 32404 21916
rect 32456 21904 32462 21956
rect 22557 21879 22615 21885
rect 22557 21845 22569 21879
rect 22603 21876 22615 21879
rect 23106 21876 23112 21888
rect 22603 21848 23112 21876
rect 22603 21845 22615 21848
rect 22557 21839 22615 21845
rect 23106 21836 23112 21848
rect 23164 21876 23170 21888
rect 23293 21879 23351 21885
rect 23293 21876 23305 21879
rect 23164 21848 23305 21876
rect 23164 21836 23170 21848
rect 23293 21845 23305 21848
rect 23339 21845 23351 21879
rect 23293 21839 23351 21845
rect 23382 21836 23388 21888
rect 23440 21876 23446 21888
rect 23440 21848 23485 21876
rect 23440 21836 23446 21848
rect 23566 21836 23572 21888
rect 23624 21876 23630 21888
rect 23661 21879 23719 21885
rect 23661 21876 23673 21879
rect 23624 21848 23673 21876
rect 23624 21836 23630 21848
rect 23661 21845 23673 21848
rect 23707 21845 23719 21879
rect 23661 21839 23719 21845
rect 28810 21836 28816 21888
rect 28868 21876 28874 21888
rect 28868 21848 28913 21876
rect 28868 21836 28874 21848
rect 29454 21836 29460 21888
rect 29512 21876 29518 21888
rect 29733 21879 29791 21885
rect 29733 21876 29745 21879
rect 29512 21848 29745 21876
rect 29512 21836 29518 21848
rect 29733 21845 29745 21848
rect 29779 21845 29791 21879
rect 30374 21876 30380 21888
rect 30335 21848 30380 21876
rect 29733 21839 29791 21845
rect 30374 21836 30380 21848
rect 30432 21836 30438 21888
rect 33980 21876 34008 22052
rect 34057 22049 34069 22083
rect 34103 22080 34115 22083
rect 46017 22083 46075 22089
rect 34103 22052 37872 22080
rect 34103 22049 34115 22052
rect 34057 22043 34115 22049
rect 35161 22015 35219 22021
rect 35161 21981 35173 22015
rect 35207 22012 35219 22015
rect 35342 22012 35348 22024
rect 35207 21984 35348 22012
rect 35207 21981 35219 21984
rect 35161 21975 35219 21981
rect 35342 21972 35348 21984
rect 35400 21972 35406 22024
rect 36265 22015 36323 22021
rect 36265 21981 36277 22015
rect 36311 22012 36323 22015
rect 36354 22012 36360 22024
rect 36311 21984 36360 22012
rect 36311 21981 36323 21984
rect 36265 21975 36323 21981
rect 36354 21972 36360 21984
rect 36412 22012 36418 22024
rect 36630 22012 36636 22024
rect 36412 21984 36636 22012
rect 36412 21972 36418 21984
rect 36630 21972 36636 21984
rect 36688 21972 36694 22024
rect 37553 22015 37611 22021
rect 37553 21981 37565 22015
rect 37599 22012 37611 22015
rect 37734 22012 37740 22024
rect 37599 21984 37740 22012
rect 37599 21981 37611 21984
rect 37553 21975 37611 21981
rect 37734 21972 37740 21984
rect 37792 21972 37798 22024
rect 36909 21947 36967 21953
rect 36909 21913 36921 21947
rect 36955 21944 36967 21947
rect 36998 21944 37004 21956
rect 36955 21916 37004 21944
rect 36955 21913 36967 21916
rect 36909 21907 36967 21913
rect 36998 21904 37004 21916
rect 37056 21904 37062 21956
rect 37844 21944 37872 22052
rect 46017 22049 46029 22083
rect 46063 22049 46075 22083
rect 46017 22043 46075 22049
rect 38838 21972 38844 22024
rect 38896 22012 38902 22024
rect 39117 22015 39175 22021
rect 39117 22012 39129 22015
rect 38896 21984 39129 22012
rect 38896 21972 38902 21984
rect 39117 21981 39129 21984
rect 39163 21981 39175 22015
rect 39117 21975 39175 21981
rect 39758 21972 39764 22024
rect 39816 22012 39822 22024
rect 39853 22015 39911 22021
rect 39853 22012 39865 22015
rect 39816 21984 39865 22012
rect 39816 21972 39822 21984
rect 39853 21981 39865 21984
rect 39899 21981 39911 22015
rect 40034 22012 40040 22024
rect 39995 21984 40040 22012
rect 39853 21975 39911 21981
rect 40034 21972 40040 21984
rect 40092 21972 40098 22024
rect 42426 22012 42432 22024
rect 40144 21984 42432 22012
rect 40144 21944 40172 21984
rect 42426 21972 42432 21984
rect 42484 21972 42490 22024
rect 45186 22012 45192 22024
rect 45147 21984 45192 22012
rect 45186 21972 45192 21984
rect 45244 21972 45250 22024
rect 45370 22012 45376 22024
rect 45331 21984 45376 22012
rect 45370 21972 45376 21984
rect 45428 21972 45434 22024
rect 45830 22012 45836 22024
rect 45791 21984 45836 22012
rect 45830 21972 45836 21984
rect 45888 21972 45894 22024
rect 37844 21916 40172 21944
rect 40221 21947 40279 21953
rect 40221 21913 40233 21947
rect 40267 21944 40279 21947
rect 40310 21944 40316 21956
rect 40267 21916 40316 21944
rect 40267 21913 40279 21916
rect 40221 21907 40279 21913
rect 40310 21904 40316 21916
rect 40368 21904 40374 21956
rect 42702 21944 42708 21956
rect 42663 21916 42708 21944
rect 42702 21904 42708 21916
rect 42760 21904 42766 21956
rect 45554 21944 45560 21956
rect 43029 21916 45560 21944
rect 38286 21876 38292 21888
rect 33980 21848 38292 21876
rect 38286 21836 38292 21848
rect 38344 21836 38350 21888
rect 38562 21836 38568 21888
rect 38620 21876 38626 21888
rect 43029 21876 43057 21916
rect 45554 21904 45560 21916
rect 45612 21904 45618 21956
rect 45738 21904 45744 21956
rect 45796 21944 45802 21956
rect 46566 21944 46572 21956
rect 45796 21916 46572 21944
rect 45796 21904 45802 21916
rect 46566 21904 46572 21916
rect 46624 21904 46630 21956
rect 47210 21904 47216 21956
rect 47268 21944 47274 21956
rect 47673 21947 47731 21953
rect 47673 21944 47685 21947
rect 47268 21916 47685 21944
rect 47268 21904 47274 21916
rect 47673 21913 47685 21916
rect 47719 21913 47731 21947
rect 47673 21907 47731 21913
rect 43162 21876 43168 21888
rect 38620 21848 43057 21876
rect 43123 21848 43168 21876
rect 38620 21836 38626 21848
rect 43162 21836 43168 21848
rect 43220 21836 43226 21888
rect 45373 21879 45431 21885
rect 45373 21845 45385 21879
rect 45419 21876 45431 21879
rect 46658 21876 46664 21888
rect 45419 21848 46664 21876
rect 45419 21845 45431 21848
rect 45373 21839 45431 21845
rect 46658 21836 46664 21848
rect 46716 21836 46722 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 11698 21672 11704 21684
rect 11659 21644 11704 21672
rect 11698 21632 11704 21644
rect 11756 21632 11762 21684
rect 20438 21632 20444 21684
rect 20496 21672 20502 21684
rect 24302 21672 24308 21684
rect 20496 21644 21312 21672
rect 20496 21632 20502 21644
rect 6886 21576 12434 21604
rect 3786 21428 3792 21480
rect 3844 21468 3850 21480
rect 6886 21468 6914 21576
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21505 10839 21539
rect 10781 21499 10839 21505
rect 3844 21440 6914 21468
rect 10796 21468 10824 21499
rect 10870 21496 10876 21548
rect 10928 21536 10934 21548
rect 10965 21539 11023 21545
rect 10965 21536 10977 21539
rect 10928 21508 10977 21536
rect 10928 21496 10934 21508
rect 10965 21505 10977 21508
rect 11011 21505 11023 21539
rect 11514 21536 11520 21548
rect 11475 21508 11520 21536
rect 10965 21499 11023 21505
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 12250 21536 12256 21548
rect 12211 21508 12256 21536
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 12406 21536 12434 21576
rect 13722 21564 13728 21616
rect 13780 21604 13786 21616
rect 17678 21604 17684 21616
rect 13780 21576 17684 21604
rect 13780 21564 13786 21576
rect 17678 21564 17684 21576
rect 17736 21564 17742 21616
rect 19705 21607 19763 21613
rect 19705 21573 19717 21607
rect 19751 21604 19763 21607
rect 19978 21604 19984 21616
rect 19751 21576 19984 21604
rect 19751 21573 19763 21576
rect 19705 21567 19763 21573
rect 19978 21564 19984 21576
rect 20036 21564 20042 21616
rect 21082 21604 21088 21616
rect 20930 21576 21088 21604
rect 21082 21564 21088 21576
rect 21140 21564 21146 21616
rect 12406 21508 13492 21536
rect 12618 21468 12624 21480
rect 10796 21440 12624 21468
rect 3844 21428 3850 21440
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 10410 21360 10416 21412
rect 10468 21400 10474 21412
rect 13464 21400 13492 21508
rect 16390 21496 16396 21548
rect 16448 21536 16454 21548
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16448 21508 16865 21536
rect 16448 21496 16454 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 19426 21536 19432 21548
rect 19387 21508 19432 21536
rect 16853 21499 16911 21505
rect 13538 21428 13544 21480
rect 13596 21468 13602 21480
rect 13722 21468 13728 21480
rect 13596 21440 13641 21468
rect 13683 21440 13728 21468
rect 13596 21428 13602 21440
rect 13722 21428 13728 21440
rect 13780 21428 13786 21480
rect 14001 21471 14059 21477
rect 14001 21437 14013 21471
rect 14047 21437 14059 21471
rect 16868 21468 16896 21499
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 21284 21536 21312 21644
rect 22848 21644 24308 21672
rect 22848 21604 22876 21644
rect 24302 21632 24308 21644
rect 24360 21632 24366 21684
rect 24397 21675 24455 21681
rect 24397 21641 24409 21675
rect 24443 21672 24455 21675
rect 24762 21672 24768 21684
rect 24443 21644 24768 21672
rect 24443 21641 24455 21644
rect 24397 21635 24455 21641
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 27890 21632 27896 21684
rect 27948 21672 27954 21684
rect 28353 21675 28411 21681
rect 28353 21672 28365 21675
rect 27948 21644 28365 21672
rect 27948 21632 27954 21644
rect 28353 21641 28365 21644
rect 28399 21641 28411 21675
rect 28353 21635 28411 21641
rect 28442 21632 28448 21684
rect 28500 21672 28506 21684
rect 28500 21644 31754 21672
rect 28500 21632 28506 21644
rect 22020 21576 22876 21604
rect 23845 21607 23903 21613
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21284 21508 21833 21536
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 21910 21496 21916 21548
rect 21968 21536 21974 21548
rect 22020 21536 22048 21576
rect 23845 21573 23857 21607
rect 23891 21604 23903 21607
rect 28169 21607 28227 21613
rect 28169 21604 28181 21607
rect 23891 21576 28181 21604
rect 23891 21573 23903 21576
rect 23845 21567 23903 21573
rect 21968 21508 22048 21536
rect 21968 21496 21974 21508
rect 22278 21496 22284 21548
rect 22336 21536 22342 21548
rect 22557 21539 22615 21545
rect 22557 21536 22569 21539
rect 22336 21508 22569 21536
rect 22336 21496 22342 21508
rect 22557 21505 22569 21508
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 23106 21496 23112 21548
rect 23164 21536 23170 21548
rect 23290 21536 23296 21548
rect 23164 21508 23296 21536
rect 23164 21496 23170 21508
rect 23290 21496 23296 21508
rect 23348 21496 23354 21548
rect 23566 21536 23572 21548
rect 23527 21508 23572 21536
rect 23566 21496 23572 21508
rect 23624 21496 23630 21548
rect 23658 21496 23664 21548
rect 23716 21536 23722 21548
rect 23716 21508 23761 21536
rect 23716 21496 23722 21508
rect 23934 21496 23940 21548
rect 23992 21536 23998 21548
rect 24504 21545 24532 21576
rect 28169 21573 28181 21576
rect 28215 21604 28227 21607
rect 28215 21576 28396 21604
rect 28215 21573 28227 21576
rect 28169 21567 28227 21573
rect 28368 21548 28396 21576
rect 30374 21564 30380 21616
rect 30432 21564 30438 21616
rect 24305 21539 24363 21545
rect 24305 21536 24317 21539
rect 23992 21508 24317 21536
rect 23992 21496 23998 21508
rect 24305 21505 24317 21508
rect 24351 21505 24363 21539
rect 24305 21499 24363 21505
rect 24489 21539 24547 21545
rect 24489 21505 24501 21539
rect 24535 21505 24547 21539
rect 24489 21499 24547 21505
rect 25222 21496 25228 21548
rect 25280 21536 25286 21548
rect 25409 21539 25467 21545
rect 25409 21536 25421 21539
rect 25280 21508 25421 21536
rect 25280 21496 25286 21508
rect 25409 21505 25421 21508
rect 25455 21505 25467 21539
rect 25409 21499 25467 21505
rect 25498 21496 25504 21548
rect 25556 21536 25562 21548
rect 26973 21539 27031 21545
rect 26973 21536 26985 21539
rect 25556 21508 26985 21536
rect 25556 21496 25562 21508
rect 26973 21505 26985 21508
rect 27019 21536 27031 21539
rect 27798 21536 27804 21548
rect 27019 21508 27804 21536
rect 27019 21505 27031 21508
rect 26973 21499 27031 21505
rect 27798 21496 27804 21508
rect 27856 21496 27862 21548
rect 27890 21496 27896 21548
rect 27948 21536 27954 21548
rect 27985 21539 28043 21545
rect 27985 21536 27997 21539
rect 27948 21508 27997 21536
rect 27948 21496 27954 21508
rect 27985 21505 27997 21508
rect 28031 21505 28043 21539
rect 27985 21499 28043 21505
rect 28077 21539 28135 21545
rect 28077 21505 28089 21539
rect 28123 21505 28135 21539
rect 28077 21499 28135 21505
rect 21726 21468 21732 21480
rect 16868 21440 21732 21468
rect 14001 21431 14059 21437
rect 14016 21400 14044 21431
rect 21726 21428 21732 21440
rect 21784 21428 21790 21480
rect 28092 21468 28120 21499
rect 28350 21496 28356 21548
rect 28408 21496 28414 21548
rect 28810 21536 28816 21548
rect 28771 21508 28816 21536
rect 28810 21496 28816 21508
rect 28868 21496 28874 21548
rect 28994 21536 29000 21548
rect 28955 21508 29000 21536
rect 28994 21496 29000 21508
rect 29052 21496 29058 21548
rect 29454 21536 29460 21548
rect 29415 21508 29460 21536
rect 29454 21496 29460 21508
rect 29512 21496 29518 21548
rect 31726 21536 31754 21644
rect 34514 21632 34520 21684
rect 34572 21672 34578 21684
rect 42705 21675 42763 21681
rect 34572 21644 34744 21672
rect 34572 21632 34578 21644
rect 33410 21564 33416 21616
rect 33468 21604 33474 21616
rect 33505 21607 33563 21613
rect 33505 21604 33517 21607
rect 33468 21576 33517 21604
rect 33468 21564 33474 21576
rect 33505 21573 33517 21576
rect 33551 21573 33563 21607
rect 34606 21604 34612 21616
rect 34567 21576 34612 21604
rect 33505 21567 33563 21573
rect 34606 21564 34612 21576
rect 34664 21564 34670 21616
rect 34716 21613 34744 21644
rect 42705 21641 42717 21675
rect 42751 21672 42763 21675
rect 42794 21672 42800 21684
rect 42751 21644 42800 21672
rect 42751 21641 42763 21644
rect 42705 21635 42763 21641
rect 42794 21632 42800 21644
rect 42852 21632 42858 21684
rect 42886 21632 42892 21684
rect 42944 21672 42950 21684
rect 45557 21675 45615 21681
rect 42944 21644 44864 21672
rect 42944 21632 42950 21644
rect 34701 21607 34759 21613
rect 34701 21573 34713 21607
rect 34747 21573 34759 21607
rect 34701 21567 34759 21573
rect 34790 21564 34796 21616
rect 34848 21604 34854 21616
rect 38194 21604 38200 21616
rect 34848 21576 38200 21604
rect 34848 21564 34854 21576
rect 38194 21564 38200 21576
rect 38252 21564 38258 21616
rect 43717 21607 43775 21613
rect 43717 21604 43729 21607
rect 43180 21576 43729 21604
rect 32217 21539 32275 21545
rect 32217 21536 32229 21539
rect 31726 21508 32229 21536
rect 32217 21505 32229 21508
rect 32263 21505 32275 21539
rect 36354 21536 36360 21548
rect 36267 21508 36360 21536
rect 32217 21499 32275 21505
rect 28166 21468 28172 21480
rect 28092 21440 28172 21468
rect 28166 21428 28172 21440
rect 28224 21428 28230 21480
rect 29733 21471 29791 21477
rect 29733 21437 29745 21471
rect 29779 21468 29791 21471
rect 30098 21468 30104 21480
rect 29779 21440 30104 21468
rect 29779 21437 29791 21440
rect 29733 21431 29791 21437
rect 30098 21428 30104 21440
rect 30156 21428 30162 21480
rect 31202 21468 31208 21480
rect 31163 21440 31208 21468
rect 31202 21428 31208 21440
rect 31260 21428 31266 21480
rect 10468 21372 13400 21400
rect 13464 21372 14044 21400
rect 10468 21360 10474 21372
rect 10686 21292 10692 21344
rect 10744 21332 10750 21344
rect 10781 21335 10839 21341
rect 10781 21332 10793 21335
rect 10744 21304 10793 21332
rect 10744 21292 10750 21304
rect 10781 21301 10793 21304
rect 10827 21301 10839 21335
rect 12342 21332 12348 21344
rect 12303 21304 12348 21332
rect 10781 21295 10839 21301
rect 12342 21292 12348 21304
rect 12400 21292 12406 21344
rect 13372 21332 13400 21372
rect 14458 21360 14464 21412
rect 14516 21400 14522 21412
rect 17037 21403 17095 21409
rect 17037 21400 17049 21403
rect 14516 21372 17049 21400
rect 14516 21360 14522 21372
rect 17037 21369 17049 21372
rect 17083 21400 17095 21403
rect 18138 21400 18144 21412
rect 17083 21372 18144 21400
rect 17083 21369 17095 21372
rect 17037 21363 17095 21369
rect 18138 21360 18144 21372
rect 18196 21360 18202 21412
rect 27338 21360 27344 21412
rect 27396 21400 27402 21412
rect 27801 21403 27859 21409
rect 27801 21400 27813 21403
rect 27396 21372 27813 21400
rect 27396 21360 27402 21372
rect 27801 21369 27813 21372
rect 27847 21369 27859 21403
rect 27801 21363 27859 21369
rect 16850 21332 16856 21344
rect 13372 21304 16856 21332
rect 16850 21292 16856 21304
rect 16908 21292 16914 21344
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 21177 21335 21235 21341
rect 21177 21332 21189 21335
rect 19392 21304 21189 21332
rect 19392 21292 19398 21304
rect 21177 21301 21189 21304
rect 21223 21332 21235 21335
rect 21450 21332 21456 21344
rect 21223 21304 21456 21332
rect 21223 21301 21235 21304
rect 21177 21295 21235 21301
rect 21450 21292 21456 21304
rect 21508 21292 21514 21344
rect 21542 21292 21548 21344
rect 21600 21332 21606 21344
rect 21821 21335 21879 21341
rect 21821 21332 21833 21335
rect 21600 21304 21833 21332
rect 21600 21292 21606 21304
rect 21821 21301 21833 21304
rect 21867 21301 21879 21335
rect 21821 21295 21879 21301
rect 22554 21292 22560 21344
rect 22612 21332 22618 21344
rect 22649 21335 22707 21341
rect 22649 21332 22661 21335
rect 22612 21304 22661 21332
rect 22612 21292 22618 21304
rect 22649 21301 22661 21304
rect 22695 21301 22707 21335
rect 25498 21332 25504 21344
rect 25459 21304 25504 21332
rect 22649 21295 22707 21301
rect 25498 21292 25504 21304
rect 25556 21292 25562 21344
rect 26970 21292 26976 21344
rect 27028 21332 27034 21344
rect 27065 21335 27123 21341
rect 27065 21332 27077 21335
rect 27028 21304 27077 21332
rect 27028 21292 27034 21304
rect 27065 21301 27077 21304
rect 27111 21301 27123 21335
rect 27065 21295 27123 21301
rect 27982 21292 27988 21344
rect 28040 21332 28046 21344
rect 28813 21335 28871 21341
rect 28813 21332 28825 21335
rect 28040 21304 28825 21332
rect 28040 21292 28046 21304
rect 28813 21301 28825 21304
rect 28859 21301 28871 21335
rect 32232 21332 32260 21499
rect 36354 21496 36360 21508
rect 36412 21496 36418 21548
rect 37734 21536 37740 21548
rect 37695 21508 37740 21536
rect 37734 21496 37740 21508
rect 37792 21496 37798 21548
rect 41690 21536 41696 21548
rect 41651 21508 41696 21536
rect 41690 21496 41696 21508
rect 41748 21496 41754 21548
rect 41874 21536 41880 21548
rect 41835 21508 41880 21536
rect 41874 21496 41880 21508
rect 41932 21496 41938 21548
rect 42889 21539 42947 21545
rect 42889 21505 42901 21539
rect 42935 21536 42947 21539
rect 43070 21536 43076 21548
rect 42935 21508 43076 21536
rect 42935 21505 42947 21508
rect 42889 21499 42947 21505
rect 43070 21496 43076 21508
rect 43128 21536 43134 21548
rect 43180 21536 43208 21576
rect 43717 21573 43729 21576
rect 43763 21573 43775 21607
rect 43717 21567 43775 21573
rect 43622 21536 43628 21548
rect 43128 21508 43208 21536
rect 43583 21508 43628 21536
rect 43128 21496 43134 21508
rect 43622 21496 43628 21508
rect 43680 21496 43686 21548
rect 43806 21496 43812 21548
rect 43864 21536 43870 21548
rect 43864 21508 43909 21536
rect 43864 21496 43870 21508
rect 44266 21496 44272 21548
rect 44324 21536 44330 21548
rect 44729 21539 44787 21545
rect 44729 21536 44741 21539
rect 44324 21508 44741 21536
rect 44324 21496 44330 21508
rect 44729 21505 44741 21508
rect 44775 21505 44787 21539
rect 44836 21536 44864 21644
rect 45557 21641 45569 21675
rect 45603 21672 45615 21675
rect 45830 21672 45836 21684
rect 45603 21644 45836 21672
rect 45603 21641 45615 21644
rect 45557 21635 45615 21641
rect 45830 21632 45836 21644
rect 45888 21632 45894 21684
rect 47578 21632 47584 21684
rect 47636 21672 47642 21684
rect 47765 21675 47823 21681
rect 47765 21672 47777 21675
rect 47636 21644 47777 21672
rect 47636 21632 47642 21644
rect 47765 21641 47777 21644
rect 47811 21641 47823 21675
rect 47765 21635 47823 21641
rect 47949 21675 48007 21681
rect 47949 21641 47961 21675
rect 47995 21672 48007 21675
rect 48130 21672 48136 21684
rect 47995 21644 48136 21672
rect 47995 21641 48007 21644
rect 47949 21635 48007 21641
rect 45370 21564 45376 21616
rect 45428 21604 45434 21616
rect 46658 21604 46664 21616
rect 45428 21576 46520 21604
rect 46619 21576 46664 21604
rect 45428 21564 45434 21576
rect 45738 21536 45744 21548
rect 44836 21508 45744 21536
rect 44729 21499 44787 21505
rect 45738 21496 45744 21508
rect 45796 21496 45802 21548
rect 46201 21539 46259 21545
rect 46201 21505 46213 21539
rect 46247 21505 46259 21539
rect 46492 21536 46520 21576
rect 46658 21564 46664 21576
rect 46716 21564 46722 21616
rect 46845 21607 46903 21613
rect 46845 21573 46857 21607
rect 46891 21604 46903 21607
rect 47596 21604 47624 21632
rect 46891 21576 47624 21604
rect 46891 21573 46903 21576
rect 46845 21567 46903 21573
rect 47581 21539 47639 21545
rect 47581 21536 47593 21539
rect 46492 21508 47593 21536
rect 46201 21499 46259 21505
rect 47581 21505 47593 21508
rect 47627 21536 47639 21539
rect 47670 21536 47676 21548
rect 47627 21508 47676 21536
rect 47627 21505 47639 21508
rect 47581 21499 47639 21505
rect 32769 21471 32827 21477
rect 32769 21437 32781 21471
rect 32815 21468 32827 21471
rect 32858 21468 32864 21480
rect 32815 21440 32864 21468
rect 32815 21437 32827 21440
rect 32769 21431 32827 21437
rect 32858 21428 32864 21440
rect 32916 21428 32922 21480
rect 33413 21471 33471 21477
rect 33413 21437 33425 21471
rect 33459 21468 33471 21471
rect 35526 21468 35532 21480
rect 33459 21440 35532 21468
rect 33459 21437 33471 21440
rect 33413 21431 33471 21437
rect 35526 21428 35532 21440
rect 35584 21428 35590 21480
rect 35621 21471 35679 21477
rect 35621 21437 35633 21471
rect 35667 21468 35679 21471
rect 36262 21468 36268 21480
rect 35667 21440 36268 21468
rect 35667 21437 35679 21440
rect 35621 21431 35679 21437
rect 36262 21428 36268 21440
rect 36320 21428 36326 21480
rect 32306 21360 32312 21412
rect 32364 21400 32370 21412
rect 33965 21403 34023 21409
rect 33965 21400 33977 21403
rect 32364 21372 33977 21400
rect 32364 21360 32370 21372
rect 33965 21369 33977 21372
rect 34011 21369 34023 21403
rect 36372 21400 36400 21496
rect 38286 21468 38292 21480
rect 38247 21440 38292 21468
rect 38286 21428 38292 21440
rect 38344 21428 38350 21480
rect 41785 21471 41843 21477
rect 41785 21437 41797 21471
rect 41831 21468 41843 21471
rect 42702 21468 42708 21480
rect 41831 21440 42708 21468
rect 41831 21437 41843 21440
rect 41785 21431 41843 21437
rect 42702 21428 42708 21440
rect 42760 21468 42766 21480
rect 43165 21471 43223 21477
rect 43165 21468 43177 21471
rect 42760 21440 43177 21468
rect 42760 21428 42766 21440
rect 43165 21437 43177 21440
rect 43211 21437 43223 21471
rect 45002 21468 45008 21480
rect 44963 21440 45008 21468
rect 43165 21431 43223 21437
rect 45002 21428 45008 21440
rect 45060 21428 45066 21480
rect 46216 21468 46244 21499
rect 47670 21496 47676 21508
rect 47728 21496 47734 21548
rect 47854 21536 47860 21548
rect 47815 21508 47860 21536
rect 47854 21496 47860 21508
rect 47912 21496 47918 21548
rect 47029 21471 47087 21477
rect 47029 21468 47041 21471
rect 46216 21440 47041 21468
rect 47029 21437 47041 21440
rect 47075 21437 47087 21471
rect 47029 21431 47087 21437
rect 47762 21428 47768 21480
rect 47820 21468 47826 21480
rect 47964 21468 47992 21635
rect 48130 21632 48136 21644
rect 48188 21632 48194 21684
rect 47820 21440 47992 21468
rect 47820 21428 47826 21440
rect 33965 21363 34023 21369
rect 36280 21372 36400 21400
rect 36280 21332 36308 21372
rect 41874 21360 41880 21412
rect 41932 21400 41938 21412
rect 43806 21400 43812 21412
rect 41932 21372 43812 21400
rect 41932 21360 41938 21372
rect 43806 21360 43812 21372
rect 43864 21360 43870 21412
rect 48130 21400 48136 21412
rect 48091 21372 48136 21400
rect 48130 21360 48136 21372
rect 48188 21360 48194 21412
rect 36630 21332 36636 21344
rect 32232 21304 36308 21332
rect 36591 21304 36636 21332
rect 28813 21295 28871 21301
rect 36630 21292 36636 21304
rect 36688 21292 36694 21344
rect 36998 21292 37004 21344
rect 37056 21332 37062 21344
rect 42886 21332 42892 21344
rect 37056 21304 42892 21332
rect 37056 21292 37062 21304
rect 42886 21292 42892 21304
rect 42944 21292 42950 21344
rect 43070 21332 43076 21344
rect 43031 21304 43076 21332
rect 43070 21292 43076 21304
rect 43128 21292 43134 21344
rect 46014 21332 46020 21344
rect 45975 21304 46020 21332
rect 46014 21292 46020 21304
rect 46072 21292 46078 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 2590 21088 2596 21140
rect 2648 21128 2654 21140
rect 10410 21128 10416 21140
rect 2648 21100 10416 21128
rect 2648 21088 2654 21100
rect 10410 21088 10416 21100
rect 10468 21088 10474 21140
rect 12066 21088 12072 21140
rect 12124 21128 12130 21140
rect 12161 21131 12219 21137
rect 12161 21128 12173 21131
rect 12124 21100 12173 21128
rect 12124 21088 12130 21100
rect 12161 21097 12173 21100
rect 12207 21097 12219 21131
rect 12618 21128 12624 21140
rect 12579 21100 12624 21128
rect 12161 21091 12219 21097
rect 12618 21088 12624 21100
rect 12676 21088 12682 21140
rect 13722 21088 13728 21140
rect 13780 21128 13786 21140
rect 14921 21131 14979 21137
rect 14921 21128 14933 21131
rect 13780 21100 14933 21128
rect 13780 21088 13786 21100
rect 14921 21097 14933 21100
rect 14967 21097 14979 21131
rect 16206 21128 16212 21140
rect 16167 21100 16212 21128
rect 14921 21091 14979 21097
rect 16206 21088 16212 21100
rect 16264 21088 16270 21140
rect 16393 21131 16451 21137
rect 16393 21097 16405 21131
rect 16439 21128 16451 21131
rect 16482 21128 16488 21140
rect 16439 21100 16488 21128
rect 16439 21097 16451 21100
rect 16393 21091 16451 21097
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 16850 21088 16856 21140
rect 16908 21128 16914 21140
rect 23290 21128 23296 21140
rect 16908 21100 23152 21128
rect 23251 21100 23296 21128
rect 16908 21088 16914 21100
rect 3970 21020 3976 21072
rect 4028 21060 4034 21072
rect 10318 21060 10324 21072
rect 4028 21032 10324 21060
rect 4028 21020 4034 21032
rect 10318 21020 10324 21032
rect 10376 21020 10382 21072
rect 14366 21020 14372 21072
rect 14424 21060 14430 21072
rect 23124 21060 23152 21100
rect 23290 21088 23296 21100
rect 23348 21088 23354 21140
rect 24670 21128 24676 21140
rect 24631 21100 24676 21128
rect 24670 21088 24676 21100
rect 24728 21088 24734 21140
rect 27798 21128 27804 21140
rect 25240 21100 27804 21128
rect 25240 21060 25268 21100
rect 27798 21088 27804 21100
rect 27856 21088 27862 21140
rect 28166 21088 28172 21140
rect 28224 21128 28230 21140
rect 28261 21131 28319 21137
rect 28261 21128 28273 21131
rect 28224 21100 28273 21128
rect 28224 21088 28230 21100
rect 28261 21097 28273 21100
rect 28307 21128 28319 21131
rect 28442 21128 28448 21140
rect 28307 21100 28448 21128
rect 28307 21097 28319 21100
rect 28261 21091 28319 21097
rect 28442 21088 28448 21100
rect 28500 21088 28506 21140
rect 30098 21128 30104 21140
rect 28552 21100 29868 21128
rect 30059 21100 30104 21128
rect 28552 21060 28580 21100
rect 14424 21032 21680 21060
rect 23124 21032 25268 21060
rect 25332 21032 28580 21060
rect 29840 21060 29868 21100
rect 30098 21088 30104 21100
rect 30156 21088 30162 21140
rect 32674 21128 32680 21140
rect 32635 21100 32680 21128
rect 32674 21088 32680 21100
rect 32732 21088 32738 21140
rect 33410 21128 33416 21140
rect 33371 21100 33416 21128
rect 33410 21088 33416 21100
rect 33468 21088 33474 21140
rect 36262 21088 36268 21140
rect 36320 21128 36326 21140
rect 42702 21128 42708 21140
rect 36320 21100 42708 21128
rect 36320 21088 36326 21100
rect 42702 21088 42708 21100
rect 42760 21088 42766 21140
rect 42996 21100 43208 21128
rect 29840 21032 31892 21060
rect 14424 21020 14430 21032
rect 3418 20952 3424 21004
rect 3476 20992 3482 21004
rect 13998 20992 14004 21004
rect 3476 20964 14004 20992
rect 3476 20952 3482 20964
rect 13998 20952 14004 20964
rect 14056 20952 14062 21004
rect 20438 20952 20444 21004
rect 20496 20992 20502 21004
rect 20533 20995 20591 21001
rect 20533 20992 20545 20995
rect 20496 20964 20545 20992
rect 20496 20952 20502 20964
rect 20533 20961 20545 20964
rect 20579 20961 20591 20995
rect 21542 20992 21548 21004
rect 21503 20964 21548 20992
rect 20533 20955 20591 20961
rect 21542 20952 21548 20964
rect 21600 20952 21606 21004
rect 21652 20992 21680 21032
rect 25332 20992 25360 21032
rect 25498 20992 25504 21004
rect 21652 20964 25360 20992
rect 25459 20964 25504 20992
rect 25498 20952 25504 20964
rect 25556 20952 25562 21004
rect 26697 20995 26755 21001
rect 26697 20961 26709 20995
rect 26743 20961 26755 20995
rect 26697 20955 26755 20961
rect 10410 20924 10416 20936
rect 10371 20896 10416 20924
rect 10410 20884 10416 20896
rect 10468 20884 10474 20936
rect 12066 20884 12072 20936
rect 12124 20924 12130 20936
rect 12621 20927 12679 20933
rect 12621 20924 12633 20927
rect 12124 20896 12633 20924
rect 12124 20884 12130 20896
rect 12621 20893 12633 20896
rect 12667 20893 12679 20927
rect 12894 20924 12900 20936
rect 12855 20896 12900 20924
rect 12621 20887 12679 20893
rect 10686 20856 10692 20868
rect 10647 20828 10692 20856
rect 10686 20816 10692 20828
rect 10744 20816 10750 20868
rect 12342 20856 12348 20868
rect 11914 20828 12348 20856
rect 12342 20816 12348 20828
rect 12400 20816 12406 20868
rect 12636 20856 12664 20887
rect 12894 20884 12900 20896
rect 12952 20884 12958 20936
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20924 14151 20927
rect 14182 20924 14188 20936
rect 14139 20896 14188 20924
rect 14139 20893 14151 20896
rect 14093 20887 14151 20893
rect 14182 20884 14188 20896
rect 14240 20884 14246 20936
rect 14550 20924 14556 20936
rect 14292 20896 14556 20924
rect 12636 20828 14228 20856
rect 14200 20800 14228 20828
rect 12802 20788 12808 20800
rect 12763 20760 12808 20788
rect 12802 20748 12808 20760
rect 12860 20748 12866 20800
rect 14182 20748 14188 20800
rect 14240 20748 14246 20800
rect 14292 20797 14320 20896
rect 14550 20884 14556 20896
rect 14608 20884 14614 20936
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20924 14887 20927
rect 16574 20924 16580 20936
rect 14875 20896 16580 20924
rect 14875 20893 14887 20896
rect 14829 20887 14887 20893
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 17402 20924 17408 20936
rect 17363 20896 17408 20924
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 18138 20924 18144 20936
rect 18099 20896 18144 20924
rect 18138 20884 18144 20896
rect 18196 20884 18202 20936
rect 19242 20884 19248 20936
rect 19300 20924 19306 20936
rect 20257 20927 20315 20933
rect 20257 20924 20269 20927
rect 19300 20896 20269 20924
rect 19300 20884 19306 20896
rect 20257 20893 20269 20896
rect 20303 20924 20315 20927
rect 21450 20924 21456 20936
rect 20303 20896 21456 20924
rect 20303 20893 20315 20896
rect 20257 20887 20315 20893
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 23198 20884 23204 20936
rect 23256 20924 23262 20936
rect 24489 20927 24547 20933
rect 24489 20924 24501 20927
rect 23256 20896 24501 20924
rect 23256 20884 23262 20896
rect 24489 20893 24501 20896
rect 24535 20893 24547 20927
rect 25314 20924 25320 20936
rect 25275 20896 25320 20924
rect 24489 20887 24547 20893
rect 25314 20884 25320 20896
rect 25372 20884 25378 20936
rect 16025 20859 16083 20865
rect 16025 20825 16037 20859
rect 16071 20825 16083 20859
rect 16025 20819 16083 20825
rect 21821 20859 21879 20865
rect 21821 20825 21833 20859
rect 21867 20856 21879 20859
rect 22094 20856 22100 20868
rect 21867 20828 22100 20856
rect 21867 20825 21879 20828
rect 21821 20819 21879 20825
rect 14277 20791 14335 20797
rect 14277 20757 14289 20791
rect 14323 20757 14335 20791
rect 14277 20751 14335 20757
rect 14366 20748 14372 20800
rect 14424 20788 14430 20800
rect 16040 20788 16068 20819
rect 22094 20816 22100 20828
rect 22152 20816 22158 20868
rect 22554 20816 22560 20868
rect 22612 20816 22618 20868
rect 26712 20856 26740 20955
rect 28166 20952 28172 21004
rect 28224 20992 28230 21004
rect 28350 20992 28356 21004
rect 28224 20964 28356 20992
rect 28224 20952 28230 20964
rect 28350 20952 28356 20964
rect 28408 20992 28414 21004
rect 29641 20995 29699 21001
rect 29641 20992 29653 20995
rect 28408 20964 29653 20992
rect 28408 20952 28414 20964
rect 29641 20961 29653 20964
rect 29687 20961 29699 20995
rect 29641 20955 29699 20961
rect 31110 20952 31116 21004
rect 31168 20992 31174 21004
rect 31389 20995 31447 21001
rect 31389 20992 31401 20995
rect 31168 20964 31401 20992
rect 31168 20952 31174 20964
rect 31389 20961 31401 20964
rect 31435 20992 31447 20995
rect 31570 20992 31576 21004
rect 31435 20964 31576 20992
rect 31435 20961 31447 20964
rect 31389 20955 31447 20961
rect 31570 20952 31576 20964
rect 31628 20952 31634 21004
rect 31864 20992 31892 21032
rect 32214 21020 32220 21072
rect 32272 21060 32278 21072
rect 32272 21032 35296 21060
rect 32272 21020 32278 21032
rect 35268 21001 35296 21032
rect 35526 21020 35532 21072
rect 35584 21060 35590 21072
rect 42886 21060 42892 21072
rect 35584 21032 42892 21060
rect 35584 21020 35590 21032
rect 42886 21020 42892 21032
rect 42944 21020 42950 21072
rect 32953 20995 33011 21001
rect 31864 20964 32628 20992
rect 27798 20884 27804 20936
rect 27856 20924 27862 20936
rect 27856 20896 28396 20924
rect 27856 20884 27862 20896
rect 23216 20828 26740 20856
rect 14424 20760 16068 20788
rect 16235 20791 16293 20797
rect 14424 20748 14430 20760
rect 16235 20757 16247 20791
rect 16281 20788 16293 20791
rect 17034 20788 17040 20800
rect 16281 20760 17040 20788
rect 16281 20757 16293 20760
rect 16235 20751 16293 20757
rect 17034 20748 17040 20760
rect 17092 20748 17098 20800
rect 17589 20791 17647 20797
rect 17589 20757 17601 20791
rect 17635 20788 17647 20791
rect 17954 20788 17960 20800
rect 17635 20760 17960 20788
rect 17635 20757 17647 20760
rect 17589 20751 17647 20757
rect 17954 20748 17960 20760
rect 18012 20788 18018 20800
rect 18138 20788 18144 20800
rect 18012 20760 18144 20788
rect 18012 20748 18018 20760
rect 18138 20748 18144 20760
rect 18196 20748 18202 20800
rect 18233 20791 18291 20797
rect 18233 20757 18245 20791
rect 18279 20788 18291 20791
rect 18322 20788 18328 20800
rect 18279 20760 18328 20788
rect 18279 20757 18291 20760
rect 18233 20751 18291 20757
rect 18322 20748 18328 20760
rect 18380 20748 18386 20800
rect 18414 20748 18420 20800
rect 18472 20788 18478 20800
rect 23216 20788 23244 20828
rect 27890 20816 27896 20868
rect 27948 20856 27954 20868
rect 28077 20859 28135 20865
rect 28077 20856 28089 20859
rect 27948 20828 28089 20856
rect 27948 20816 27954 20828
rect 28077 20825 28089 20828
rect 28123 20825 28135 20859
rect 28077 20819 28135 20825
rect 28166 20816 28172 20868
rect 28224 20856 28230 20868
rect 28277 20859 28335 20865
rect 28277 20856 28289 20859
rect 28224 20828 28289 20856
rect 28224 20816 28230 20828
rect 28277 20825 28289 20828
rect 28323 20825 28335 20859
rect 28368 20856 28396 20896
rect 28442 20884 28448 20936
rect 28500 20924 28506 20936
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 28500 20896 29745 20924
rect 28500 20884 28506 20896
rect 29733 20893 29745 20896
rect 29779 20924 29791 20927
rect 31202 20924 31208 20936
rect 29779 20896 31208 20924
rect 29779 20893 29791 20896
rect 29733 20887 29791 20893
rect 31202 20884 31208 20896
rect 31260 20884 31266 20936
rect 32033 20927 32091 20933
rect 32033 20893 32045 20927
rect 32079 20924 32091 20927
rect 32306 20924 32312 20936
rect 32079 20896 32312 20924
rect 32079 20893 32091 20896
rect 32033 20887 32091 20893
rect 32306 20884 32312 20896
rect 32364 20884 32370 20936
rect 32493 20927 32551 20933
rect 32493 20893 32505 20927
rect 32539 20893 32551 20927
rect 32493 20887 32551 20893
rect 31110 20856 31116 20868
rect 28368 20828 31116 20856
rect 28277 20819 28335 20825
rect 31110 20816 31116 20828
rect 31168 20816 31174 20868
rect 31481 20859 31539 20865
rect 31481 20825 31493 20859
rect 31527 20825 31539 20859
rect 31481 20819 31539 20825
rect 18472 20760 23244 20788
rect 18472 20748 18478 20760
rect 27154 20748 27160 20800
rect 27212 20788 27218 20800
rect 28445 20791 28503 20797
rect 28445 20788 28457 20791
rect 27212 20760 28457 20788
rect 27212 20748 27218 20760
rect 28445 20757 28457 20760
rect 28491 20788 28503 20791
rect 28994 20788 29000 20800
rect 28491 20760 29000 20788
rect 28491 20757 28503 20760
rect 28445 20751 28503 20757
rect 28994 20748 29000 20760
rect 29052 20748 29058 20800
rect 30190 20748 30196 20800
rect 30248 20788 30254 20800
rect 31496 20788 31524 20819
rect 31570 20816 31576 20868
rect 31628 20856 31634 20868
rect 32214 20856 32220 20868
rect 31628 20828 32220 20856
rect 31628 20816 31634 20828
rect 32214 20816 32220 20828
rect 32272 20816 32278 20868
rect 32508 20788 32536 20887
rect 30248 20760 32536 20788
rect 32600 20788 32628 20964
rect 32953 20961 32965 20995
rect 32999 20961 33011 20995
rect 32953 20955 33011 20961
rect 35253 20995 35311 21001
rect 35253 20961 35265 20995
rect 35299 20992 35311 20995
rect 42996 20992 43024 21100
rect 43180 21060 43208 21100
rect 43622 21088 43628 21140
rect 43680 21128 43686 21140
rect 46474 21128 46480 21140
rect 43680 21100 46480 21128
rect 43680 21088 43686 21100
rect 46474 21088 46480 21100
rect 46532 21088 46538 21140
rect 45922 21060 45928 21072
rect 43180 21032 45928 21060
rect 45922 21020 45928 21032
rect 45980 21020 45986 21072
rect 35299 20964 43024 20992
rect 45189 20995 45247 21001
rect 35299 20961 35311 20964
rect 35253 20955 35311 20961
rect 45189 20961 45201 20995
rect 45235 20992 45247 20995
rect 46293 20995 46351 21001
rect 46293 20992 46305 20995
rect 45235 20964 46305 20992
rect 45235 20961 45247 20964
rect 45189 20955 45247 20961
rect 46293 20961 46305 20964
rect 46339 20961 46351 20995
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 46293 20955 46351 20961
rect 32968 20924 32996 20955
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 33597 20927 33655 20933
rect 33597 20924 33609 20927
rect 32968 20896 33609 20924
rect 33597 20893 33609 20896
rect 33643 20893 33655 20927
rect 33597 20887 33655 20893
rect 36725 20927 36783 20933
rect 36725 20893 36737 20927
rect 36771 20924 36783 20927
rect 38562 20924 38568 20936
rect 36771 20896 38568 20924
rect 36771 20893 36783 20896
rect 36725 20887 36783 20893
rect 38562 20884 38568 20896
rect 38620 20884 38626 20936
rect 42889 20927 42947 20933
rect 42889 20893 42901 20927
rect 42935 20924 42947 20927
rect 42978 20924 42984 20936
rect 42935 20896 42984 20924
rect 42935 20893 42947 20896
rect 42889 20887 42947 20893
rect 42978 20884 42984 20896
rect 43036 20884 43042 20936
rect 43070 20884 43076 20936
rect 43128 20924 43134 20936
rect 43257 20927 43315 20933
rect 43257 20924 43269 20927
rect 43128 20896 43269 20924
rect 43128 20884 43134 20896
rect 43257 20893 43269 20896
rect 43303 20924 43315 20927
rect 43714 20924 43720 20936
rect 43303 20896 43720 20924
rect 43303 20893 43315 20896
rect 43257 20887 43315 20893
rect 43714 20884 43720 20896
rect 43772 20884 43778 20936
rect 45649 20927 45707 20933
rect 45649 20893 45661 20927
rect 45695 20893 45707 20927
rect 45649 20887 45707 20893
rect 32858 20816 32864 20868
rect 32916 20856 32922 20868
rect 34790 20856 34796 20868
rect 32916 20828 34796 20856
rect 32916 20816 32922 20828
rect 34790 20816 34796 20828
rect 34848 20816 34854 20868
rect 35342 20816 35348 20868
rect 35400 20856 35406 20868
rect 36262 20856 36268 20868
rect 35400 20828 35445 20856
rect 36223 20828 36268 20856
rect 35400 20816 35406 20828
rect 36262 20816 36268 20828
rect 36320 20816 36326 20868
rect 45664 20856 45692 20887
rect 36372 20828 38884 20856
rect 36372 20788 36400 20828
rect 38856 20800 38884 20828
rect 41386 20828 45692 20856
rect 45741 20859 45799 20865
rect 36814 20788 36820 20800
rect 32600 20760 36400 20788
rect 36775 20760 36820 20788
rect 30248 20748 30254 20760
rect 36814 20748 36820 20760
rect 36872 20748 36878 20800
rect 38838 20748 38844 20800
rect 38896 20788 38902 20800
rect 41386 20788 41414 20828
rect 45741 20825 45753 20859
rect 45787 20856 45799 20859
rect 46477 20859 46535 20865
rect 46477 20856 46489 20859
rect 45787 20828 46489 20856
rect 45787 20825 45799 20828
rect 45741 20819 45799 20825
rect 46477 20825 46489 20828
rect 46523 20825 46535 20859
rect 46477 20819 46535 20825
rect 38896 20760 41414 20788
rect 38896 20748 38902 20760
rect 42886 20748 42892 20800
rect 42944 20788 42950 20800
rect 43622 20788 43628 20800
rect 42944 20760 43628 20788
rect 42944 20748 42950 20760
rect 43622 20748 43628 20760
rect 43680 20748 43686 20800
rect 43806 20748 43812 20800
rect 43864 20788 43870 20800
rect 43901 20791 43959 20797
rect 43901 20788 43913 20791
rect 43864 20760 43913 20788
rect 43864 20748 43870 20760
rect 43901 20757 43913 20760
rect 43947 20757 43959 20791
rect 43901 20751 43959 20757
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 3510 20544 3516 20596
rect 3568 20584 3574 20596
rect 3568 20556 6914 20584
rect 3568 20544 3574 20556
rect 6886 20516 6914 20556
rect 10410 20544 10416 20596
rect 10468 20584 10474 20596
rect 10505 20587 10563 20593
rect 10505 20584 10517 20587
rect 10468 20556 10517 20584
rect 10468 20544 10474 20556
rect 10505 20553 10517 20556
rect 10551 20553 10563 20587
rect 10505 20547 10563 20553
rect 12805 20587 12863 20593
rect 12805 20553 12817 20587
rect 12851 20584 12863 20587
rect 12894 20584 12900 20596
rect 12851 20556 12900 20584
rect 12851 20553 12863 20556
rect 12805 20547 12863 20553
rect 12894 20544 12900 20556
rect 12952 20584 12958 20596
rect 13906 20584 13912 20596
rect 12952 20556 13912 20584
rect 12952 20544 12958 20556
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 32214 20584 32220 20596
rect 14016 20556 32220 20584
rect 14016 20516 14044 20556
rect 32214 20544 32220 20556
rect 32272 20544 32278 20596
rect 32398 20584 32404 20596
rect 32359 20556 32404 20584
rect 32398 20544 32404 20556
rect 32456 20544 32462 20596
rect 36630 20584 36636 20596
rect 33428 20556 36636 20584
rect 6886 20488 14044 20516
rect 14093 20519 14151 20525
rect 14093 20485 14105 20519
rect 14139 20485 14151 20519
rect 14093 20479 14151 20485
rect 14309 20519 14367 20525
rect 14309 20485 14321 20519
rect 14355 20516 14367 20519
rect 14826 20516 14832 20528
rect 14355 20488 14832 20516
rect 14355 20485 14367 20488
rect 14309 20479 14367 20485
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20448 10563 20451
rect 11698 20448 11704 20460
rect 10551 20420 11704 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 12802 20448 12808 20460
rect 12763 20420 12808 20448
rect 12802 20408 12808 20420
rect 12860 20408 12866 20460
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20448 13231 20451
rect 13538 20448 13544 20460
rect 13219 20420 13544 20448
rect 13219 20417 13231 20420
rect 13173 20411 13231 20417
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 13265 20383 13323 20389
rect 13265 20349 13277 20383
rect 13311 20349 13323 20383
rect 14108 20380 14136 20479
rect 14826 20476 14832 20488
rect 14884 20516 14890 20528
rect 16853 20519 16911 20525
rect 14884 20488 15516 20516
rect 14884 20476 14890 20488
rect 14458 20408 14464 20460
rect 14516 20448 14522 20460
rect 15013 20451 15071 20457
rect 15013 20448 15025 20451
rect 14516 20420 15025 20448
rect 14516 20408 14522 20420
rect 15013 20417 15025 20420
rect 15059 20417 15071 20451
rect 15013 20411 15071 20417
rect 14366 20380 14372 20392
rect 14108 20352 14372 20380
rect 13265 20343 13323 20349
rect 3510 20272 3516 20324
rect 3568 20312 3574 20324
rect 3568 20284 12848 20312
rect 3568 20272 3574 20284
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 11112 20216 11529 20244
rect 11112 20204 11118 20216
rect 11517 20213 11529 20216
rect 11563 20213 11575 20247
rect 11517 20207 11575 20213
rect 11606 20204 11612 20256
rect 11664 20244 11670 20256
rect 12621 20247 12679 20253
rect 12621 20244 12633 20247
rect 11664 20216 12633 20244
rect 11664 20204 11670 20216
rect 12621 20213 12633 20216
rect 12667 20213 12679 20247
rect 12820 20244 12848 20284
rect 12894 20272 12900 20324
rect 12952 20312 12958 20324
rect 13280 20312 13308 20343
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 15488 20380 15516 20488
rect 16853 20485 16865 20519
rect 16899 20485 16911 20519
rect 16853 20479 16911 20485
rect 17069 20519 17127 20525
rect 17069 20485 17081 20519
rect 17115 20516 17127 20519
rect 17310 20516 17316 20528
rect 17115 20488 17316 20516
rect 17115 20485 17127 20488
rect 17069 20479 17127 20485
rect 15657 20451 15715 20457
rect 15657 20417 15669 20451
rect 15703 20448 15715 20451
rect 16574 20448 16580 20460
rect 15703 20420 16580 20448
rect 15703 20417 15715 20420
rect 15657 20411 15715 20417
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 16868 20448 16896 20479
rect 17310 20476 17316 20488
rect 17368 20516 17374 20528
rect 17494 20516 17500 20528
rect 17368 20488 17500 20516
rect 17368 20476 17374 20488
rect 17494 20476 17500 20488
rect 17552 20476 17558 20528
rect 18322 20516 18328 20528
rect 18283 20488 18328 20516
rect 18322 20476 18328 20488
rect 18380 20476 18386 20528
rect 19978 20516 19984 20528
rect 19939 20488 19984 20516
rect 19978 20476 19984 20488
rect 20036 20476 20042 20528
rect 25314 20476 25320 20528
rect 25372 20516 25378 20528
rect 27338 20516 27344 20528
rect 25372 20488 27344 20516
rect 25372 20476 25378 20488
rect 17402 20448 17408 20460
rect 16868 20420 17408 20448
rect 17402 20408 17408 20420
rect 17460 20408 17466 20460
rect 22002 20448 22008 20460
rect 21963 20420 22008 20448
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 25130 20448 25136 20460
rect 25091 20420 25136 20448
rect 25130 20408 25136 20420
rect 25188 20408 25194 20460
rect 25884 20457 25912 20488
rect 27338 20476 27344 20488
rect 27396 20476 27402 20528
rect 27982 20516 27988 20528
rect 27943 20488 27988 20516
rect 27982 20476 27988 20488
rect 28040 20476 28046 20528
rect 30009 20519 30067 20525
rect 30009 20516 30021 20519
rect 29210 20488 30021 20516
rect 30009 20485 30021 20488
rect 30055 20485 30067 20519
rect 30009 20479 30067 20485
rect 25869 20451 25927 20457
rect 25869 20417 25881 20451
rect 25915 20417 25927 20451
rect 25869 20411 25927 20417
rect 26878 20408 26884 20460
rect 26936 20448 26942 20460
rect 26973 20451 27031 20457
rect 26973 20448 26985 20451
rect 26936 20420 26985 20448
rect 26936 20408 26942 20420
rect 26973 20417 26985 20420
rect 27019 20417 27031 20451
rect 26973 20411 27031 20417
rect 29362 20408 29368 20460
rect 29420 20448 29426 20460
rect 29917 20451 29975 20457
rect 29917 20448 29929 20451
rect 29420 20420 29929 20448
rect 29420 20408 29426 20420
rect 29917 20417 29929 20420
rect 29963 20417 29975 20451
rect 29917 20411 29975 20417
rect 32309 20451 32367 20457
rect 32309 20417 32321 20451
rect 32355 20448 32367 20451
rect 33428 20448 33456 20556
rect 36630 20544 36636 20556
rect 36688 20544 36694 20596
rect 43257 20587 43315 20593
rect 43257 20553 43269 20587
rect 43303 20584 43315 20587
rect 44085 20587 44143 20593
rect 44085 20584 44097 20587
rect 43303 20556 44097 20584
rect 43303 20553 43315 20556
rect 43257 20547 43315 20553
rect 44085 20553 44097 20556
rect 44131 20553 44143 20587
rect 44085 20547 44143 20553
rect 35069 20519 35127 20525
rect 35069 20485 35081 20519
rect 35115 20516 35127 20519
rect 36814 20516 36820 20528
rect 35115 20488 36820 20516
rect 35115 20485 35127 20488
rect 35069 20479 35127 20485
rect 36814 20476 36820 20488
rect 36872 20476 36878 20528
rect 43714 20516 43720 20528
rect 43675 20488 43720 20516
rect 43714 20476 43720 20488
rect 43772 20476 43778 20528
rect 45373 20519 45431 20525
rect 45373 20485 45385 20519
rect 45419 20516 45431 20519
rect 46014 20516 46020 20528
rect 45419 20488 46020 20516
rect 45419 20485 45431 20488
rect 45373 20479 45431 20485
rect 46014 20476 46020 20488
rect 46072 20476 46078 20528
rect 47946 20516 47952 20528
rect 47907 20488 47952 20516
rect 47946 20476 47952 20488
rect 48004 20476 48010 20528
rect 32355 20420 33456 20448
rect 33505 20451 33563 20457
rect 32355 20417 32367 20420
rect 32309 20411 32367 20417
rect 33505 20417 33517 20451
rect 33551 20417 33563 20451
rect 33505 20411 33563 20417
rect 18141 20383 18199 20389
rect 15488 20352 17264 20380
rect 17236 20321 17264 20352
rect 18141 20349 18153 20383
rect 18187 20349 18199 20383
rect 18141 20343 18199 20349
rect 22097 20383 22155 20389
rect 22097 20349 22109 20383
rect 22143 20380 22155 20383
rect 22646 20380 22652 20392
rect 22143 20352 22652 20380
rect 22143 20349 22155 20352
rect 22097 20343 22155 20349
rect 14461 20315 14519 20321
rect 14461 20312 14473 20315
rect 12952 20284 14473 20312
rect 12952 20272 12958 20284
rect 14461 20281 14473 20284
rect 14507 20281 14519 20315
rect 14461 20275 14519 20281
rect 17221 20315 17279 20321
rect 17221 20281 17233 20315
rect 17267 20281 17279 20315
rect 18156 20312 18184 20343
rect 22646 20340 22652 20352
rect 22704 20340 22710 20392
rect 25961 20383 26019 20389
rect 25961 20349 25973 20383
rect 26007 20380 26019 20383
rect 27154 20380 27160 20392
rect 26007 20352 27160 20380
rect 26007 20349 26019 20352
rect 25961 20343 26019 20349
rect 27154 20340 27160 20352
rect 27212 20340 27218 20392
rect 27249 20383 27307 20389
rect 27249 20349 27261 20383
rect 27295 20380 27307 20383
rect 27709 20383 27767 20389
rect 27709 20380 27721 20383
rect 27295 20352 27721 20380
rect 27295 20349 27307 20352
rect 27249 20343 27307 20349
rect 27709 20349 27721 20352
rect 27755 20349 27767 20383
rect 32324 20380 32352 20411
rect 27709 20343 27767 20349
rect 27816 20352 32352 20380
rect 33520 20380 33548 20411
rect 42702 20408 42708 20460
rect 42760 20448 42766 20460
rect 43073 20451 43131 20457
rect 43073 20448 43085 20451
rect 42760 20420 43085 20448
rect 42760 20408 42766 20420
rect 43073 20417 43085 20420
rect 43119 20417 43131 20451
rect 43254 20448 43260 20460
rect 43215 20420 43260 20448
rect 43073 20411 43131 20417
rect 43254 20408 43260 20420
rect 43312 20408 43318 20460
rect 43898 20448 43904 20460
rect 43859 20420 43904 20448
rect 43898 20408 43904 20420
rect 43956 20408 43962 20460
rect 44177 20451 44235 20457
rect 44177 20417 44189 20451
rect 44223 20448 44235 20451
rect 44266 20448 44272 20460
rect 44223 20420 44272 20448
rect 44223 20417 44235 20420
rect 44177 20411 44235 20417
rect 44266 20408 44272 20420
rect 44324 20408 44330 20460
rect 47210 20408 47216 20460
rect 47268 20408 47274 20460
rect 33520 20352 34652 20380
rect 18230 20312 18236 20324
rect 18156 20284 18236 20312
rect 17221 20275 17279 20281
rect 18230 20272 18236 20284
rect 18288 20272 18294 20324
rect 25222 20272 25228 20324
rect 25280 20312 25286 20324
rect 27816 20312 27844 20352
rect 25280 20284 27844 20312
rect 25280 20272 25286 20284
rect 14182 20244 14188 20256
rect 12820 20216 14188 20244
rect 12621 20207 12679 20213
rect 14182 20204 14188 20216
rect 14240 20204 14246 20256
rect 14274 20204 14280 20256
rect 14332 20244 14338 20256
rect 15105 20247 15163 20253
rect 14332 20216 14377 20244
rect 14332 20204 14338 20216
rect 15105 20213 15117 20247
rect 15151 20244 15163 20247
rect 15562 20244 15568 20256
rect 15151 20216 15568 20244
rect 15151 20213 15163 20216
rect 15105 20207 15163 20213
rect 15562 20204 15568 20216
rect 15620 20204 15626 20256
rect 15746 20244 15752 20256
rect 15707 20216 15752 20244
rect 15746 20204 15752 20216
rect 15804 20204 15810 20256
rect 17034 20244 17040 20256
rect 16995 20216 17040 20244
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 22373 20247 22431 20253
rect 22373 20244 22385 20247
rect 22152 20216 22385 20244
rect 22152 20204 22158 20216
rect 22373 20213 22385 20216
rect 22419 20213 22431 20247
rect 22373 20207 22431 20213
rect 25133 20247 25191 20253
rect 25133 20213 25145 20247
rect 25179 20244 25191 20247
rect 25590 20244 25596 20256
rect 25179 20216 25596 20244
rect 25179 20213 25191 20216
rect 25133 20207 25191 20213
rect 25590 20204 25596 20216
rect 25648 20204 25654 20256
rect 25866 20204 25872 20256
rect 25924 20244 25930 20256
rect 26237 20247 26295 20253
rect 26237 20244 26249 20247
rect 25924 20216 26249 20244
rect 25924 20204 25930 20216
rect 26237 20213 26249 20216
rect 26283 20213 26295 20247
rect 29454 20244 29460 20256
rect 29415 20216 29460 20244
rect 26237 20207 26295 20213
rect 29454 20204 29460 20216
rect 29512 20204 29518 20256
rect 33502 20204 33508 20256
rect 33560 20244 33566 20256
rect 33597 20247 33655 20253
rect 33597 20244 33609 20247
rect 33560 20216 33609 20244
rect 33560 20204 33566 20216
rect 33597 20213 33609 20216
rect 33643 20213 33655 20247
rect 34624 20244 34652 20352
rect 34698 20340 34704 20392
rect 34756 20380 34762 20392
rect 34885 20383 34943 20389
rect 34885 20380 34897 20383
rect 34756 20352 34897 20380
rect 34756 20340 34762 20352
rect 34885 20349 34897 20352
rect 34931 20349 34943 20383
rect 34885 20343 34943 20349
rect 35250 20340 35256 20392
rect 35308 20380 35314 20392
rect 35345 20383 35403 20389
rect 35345 20380 35357 20383
rect 35308 20352 35357 20380
rect 35308 20340 35314 20352
rect 35345 20349 35357 20352
rect 35391 20349 35403 20383
rect 35345 20343 35403 20349
rect 43806 20340 43812 20392
rect 43864 20380 43870 20392
rect 45189 20383 45247 20389
rect 45189 20380 45201 20383
rect 43864 20352 45201 20380
rect 43864 20340 43870 20352
rect 45189 20349 45201 20352
rect 45235 20349 45247 20383
rect 45189 20343 45247 20349
rect 45554 20340 45560 20392
rect 45612 20380 45618 20392
rect 45649 20383 45707 20389
rect 45649 20380 45661 20383
rect 45612 20352 45661 20380
rect 45612 20340 45618 20352
rect 45649 20349 45661 20352
rect 45695 20380 45707 20383
rect 47228 20380 47256 20408
rect 45695 20352 47256 20380
rect 45695 20349 45707 20352
rect 45649 20343 45707 20349
rect 36538 20272 36544 20324
rect 36596 20312 36602 20324
rect 48133 20315 48191 20321
rect 48133 20312 48145 20315
rect 36596 20284 48145 20312
rect 36596 20272 36602 20284
rect 48133 20281 48145 20284
rect 48179 20281 48191 20315
rect 48133 20275 48191 20281
rect 38746 20244 38752 20256
rect 34624 20216 38752 20244
rect 33597 20207 33655 20213
rect 38746 20204 38752 20216
rect 38804 20204 38810 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 4982 20000 4988 20052
rect 5040 20040 5046 20052
rect 12805 20043 12863 20049
rect 5040 20012 12388 20040
rect 5040 20000 5046 20012
rect 12360 19972 12388 20012
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 13538 20040 13544 20052
rect 12851 20012 13544 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 14277 20043 14335 20049
rect 14277 20009 14289 20043
rect 14323 20040 14335 20043
rect 14366 20040 14372 20052
rect 14323 20012 14372 20040
rect 14323 20009 14335 20012
rect 14277 20003 14335 20009
rect 14366 20000 14372 20012
rect 14424 20000 14430 20052
rect 14458 20000 14464 20052
rect 14516 20040 14522 20052
rect 16206 20040 16212 20052
rect 14516 20012 16212 20040
rect 14516 20000 14522 20012
rect 16206 20000 16212 20012
rect 16264 20000 16270 20052
rect 27338 20040 27344 20052
rect 22066 20012 27200 20040
rect 27299 20012 27344 20040
rect 22066 19972 22094 20012
rect 12360 19944 22094 19972
rect 22738 19932 22744 19984
rect 22796 19972 22802 19984
rect 27172 19972 27200 20012
rect 27338 20000 27344 20012
rect 27396 20000 27402 20052
rect 28169 20043 28227 20049
rect 28169 20009 28181 20043
rect 28215 20040 28227 20043
rect 28810 20040 28816 20052
rect 28215 20012 28816 20040
rect 28215 20009 28227 20012
rect 28169 20003 28227 20009
rect 28810 20000 28816 20012
rect 28868 20000 28874 20052
rect 30006 20000 30012 20052
rect 30064 20040 30070 20052
rect 36538 20040 36544 20052
rect 30064 20012 36544 20040
rect 30064 20000 30070 20012
rect 36538 20000 36544 20012
rect 36596 20000 36602 20052
rect 45002 20040 45008 20052
rect 44963 20012 45008 20040
rect 45002 20000 45008 20012
rect 45060 20000 45066 20052
rect 46845 20043 46903 20049
rect 46845 20009 46857 20043
rect 46891 20040 46903 20043
rect 47762 20040 47768 20052
rect 46891 20012 47768 20040
rect 46891 20009 46903 20012
rect 46845 20003 46903 20009
rect 47762 20000 47768 20012
rect 47820 20000 47826 20052
rect 31294 19972 31300 19984
rect 22796 19944 25728 19972
rect 27172 19944 31300 19972
rect 22796 19932 22802 19944
rect 14 19864 20 19916
rect 72 19904 78 19916
rect 15746 19904 15752 19916
rect 72 19876 14964 19904
rect 15707 19876 15752 19904
rect 72 19864 78 19876
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 11054 19836 11060 19848
rect 11015 19808 11060 19836
rect 2041 19799 2099 19805
rect 11054 19796 11060 19808
rect 11112 19796 11118 19848
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 13265 19839 13323 19845
rect 13265 19836 13277 19839
rect 12676 19808 13277 19836
rect 12676 19796 12682 19808
rect 13265 19805 13277 19808
rect 13311 19836 13323 19839
rect 13814 19836 13820 19848
rect 13311 19808 13820 19836
rect 13311 19805 13323 19808
rect 13265 19799 13323 19805
rect 13814 19796 13820 19808
rect 13872 19836 13878 19848
rect 14550 19836 14556 19848
rect 13872 19808 14556 19836
rect 13872 19796 13878 19808
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 11333 19771 11391 19777
rect 11333 19737 11345 19771
rect 11379 19768 11391 19771
rect 11606 19768 11612 19780
rect 11379 19740 11612 19768
rect 11379 19737 11391 19740
rect 11333 19731 11391 19737
rect 11606 19728 11612 19740
rect 11664 19728 11670 19780
rect 13357 19771 13415 19777
rect 13357 19768 13369 19771
rect 12558 19740 13369 19768
rect 13357 19737 13369 19740
rect 13403 19737 13415 19771
rect 13357 19731 13415 19737
rect 13538 19728 13544 19780
rect 13596 19768 13602 19780
rect 14093 19771 14151 19777
rect 14093 19768 14105 19771
rect 13596 19740 14105 19768
rect 13596 19728 13602 19740
rect 14093 19737 14105 19740
rect 14139 19737 14151 19771
rect 14093 19731 14151 19737
rect 14182 19728 14188 19780
rect 14240 19768 14246 19780
rect 14936 19768 14964 19876
rect 15746 19864 15752 19876
rect 15804 19864 15810 19916
rect 16945 19907 17003 19913
rect 16945 19873 16957 19907
rect 16991 19873 17003 19907
rect 20073 19907 20131 19913
rect 20073 19904 20085 19907
rect 16945 19867 17003 19873
rect 17052 19876 20085 19904
rect 15378 19796 15384 19848
rect 15436 19836 15442 19848
rect 15565 19839 15623 19845
rect 15565 19836 15577 19839
rect 15436 19808 15577 19836
rect 15436 19796 15442 19808
rect 15565 19805 15577 19808
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 16960 19768 16988 19867
rect 14240 19740 14872 19768
rect 14936 19740 16988 19768
rect 14240 19728 14246 19740
rect 14274 19660 14280 19712
rect 14332 19709 14338 19712
rect 14332 19703 14351 19709
rect 14339 19669 14351 19703
rect 14844 19700 14872 19740
rect 17052 19700 17080 19876
rect 20073 19873 20085 19876
rect 20119 19873 20131 19907
rect 25590 19904 25596 19916
rect 25551 19876 25596 19904
rect 20073 19867 20131 19873
rect 25590 19864 25596 19876
rect 25648 19864 25654 19916
rect 25700 19904 25728 19944
rect 31294 19932 31300 19944
rect 31352 19972 31358 19984
rect 32214 19972 32220 19984
rect 31352 19944 32220 19972
rect 31352 19932 31358 19944
rect 32214 19932 32220 19944
rect 32272 19932 32278 19984
rect 34698 19972 34704 19984
rect 32876 19944 34560 19972
rect 34659 19944 34704 19972
rect 29454 19904 29460 19916
rect 25700 19876 27200 19904
rect 17862 19836 17868 19848
rect 17823 19808 17868 19836
rect 17862 19796 17868 19808
rect 17920 19796 17926 19848
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 19392 19808 19625 19836
rect 19392 19796 19398 19808
rect 19613 19805 19625 19808
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 21450 19796 21456 19848
rect 21508 19836 21514 19848
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 21508 19808 24409 19836
rect 21508 19796 21514 19808
rect 24397 19805 24409 19808
rect 24443 19836 24455 19839
rect 24486 19836 24492 19848
rect 24443 19808 24492 19836
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 26970 19796 26976 19848
rect 27028 19796 27034 19848
rect 19797 19771 19855 19777
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 20438 19768 20444 19780
rect 19843 19740 20444 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 20438 19728 20444 19740
rect 20496 19728 20502 19780
rect 22646 19728 22652 19780
rect 22704 19768 22710 19780
rect 25222 19768 25228 19780
rect 22704 19740 25228 19768
rect 22704 19728 22710 19740
rect 25222 19728 25228 19740
rect 25280 19728 25286 19780
rect 25866 19768 25872 19780
rect 25827 19740 25872 19768
rect 25866 19728 25872 19740
rect 25924 19728 25930 19780
rect 27172 19768 27200 19876
rect 28184 19876 29460 19904
rect 27890 19796 27896 19848
rect 27948 19836 27954 19848
rect 28184 19845 28212 19876
rect 29454 19864 29460 19876
rect 29512 19904 29518 19916
rect 29549 19907 29607 19913
rect 29549 19904 29561 19907
rect 29512 19876 29561 19904
rect 29512 19864 29518 19876
rect 29549 19873 29561 19876
rect 29595 19873 29607 19907
rect 32876 19904 32904 19944
rect 29549 19867 29607 19873
rect 31726 19876 32904 19904
rect 32953 19907 33011 19913
rect 28169 19839 28227 19845
rect 28169 19836 28181 19839
rect 27948 19808 28181 19836
rect 27948 19796 27954 19808
rect 28169 19805 28181 19808
rect 28215 19805 28227 19839
rect 28169 19799 28227 19805
rect 28350 19796 28356 19848
rect 28408 19836 28414 19848
rect 28445 19839 28503 19845
rect 28445 19836 28457 19839
rect 28408 19808 28457 19836
rect 28408 19796 28414 19808
rect 28445 19805 28457 19808
rect 28491 19805 28503 19839
rect 28445 19799 28503 19805
rect 27172 19740 28580 19768
rect 14844 19672 17080 19700
rect 18049 19703 18107 19709
rect 14332 19663 14351 19669
rect 18049 19669 18061 19703
rect 18095 19700 18107 19703
rect 19150 19700 19156 19712
rect 18095 19672 19156 19700
rect 18095 19669 18107 19672
rect 18049 19663 18107 19669
rect 14332 19660 14338 19663
rect 19150 19660 19156 19672
rect 19208 19660 19214 19712
rect 24581 19703 24639 19709
rect 24581 19669 24593 19703
rect 24627 19700 24639 19703
rect 25130 19700 25136 19712
rect 24627 19672 25136 19700
rect 24627 19669 24639 19672
rect 24581 19663 24639 19669
rect 25130 19660 25136 19672
rect 25188 19700 25194 19712
rect 25774 19700 25780 19712
rect 25188 19672 25780 19700
rect 25188 19660 25194 19672
rect 25774 19660 25780 19672
rect 25832 19700 25838 19712
rect 26878 19700 26884 19712
rect 25832 19672 26884 19700
rect 25832 19660 25838 19672
rect 26878 19660 26884 19672
rect 26936 19660 26942 19712
rect 28353 19703 28411 19709
rect 28353 19669 28365 19703
rect 28399 19700 28411 19703
rect 28442 19700 28448 19712
rect 28399 19672 28448 19700
rect 28399 19669 28411 19672
rect 28353 19663 28411 19669
rect 28442 19660 28448 19672
rect 28500 19660 28506 19712
rect 28552 19700 28580 19740
rect 28902 19728 28908 19780
rect 28960 19768 28966 19780
rect 29733 19771 29791 19777
rect 29733 19768 29745 19771
rect 28960 19740 29745 19768
rect 28960 19728 28966 19740
rect 29733 19737 29745 19740
rect 29779 19737 29791 19771
rect 31386 19768 31392 19780
rect 31347 19740 31392 19768
rect 29733 19731 29791 19737
rect 31386 19728 31392 19740
rect 31444 19728 31450 19780
rect 31726 19700 31754 19876
rect 32953 19873 32965 19907
rect 32999 19904 33011 19907
rect 34532 19904 34560 19944
rect 34698 19932 34704 19944
rect 34756 19932 34762 19984
rect 43898 19932 43904 19984
rect 43956 19932 43962 19984
rect 45649 19975 45707 19981
rect 45649 19941 45661 19975
rect 45695 19972 45707 19975
rect 47026 19972 47032 19984
rect 45695 19944 47032 19972
rect 45695 19941 45707 19944
rect 45649 19935 45707 19941
rect 47026 19932 47032 19944
rect 47084 19932 47090 19984
rect 35894 19904 35900 19916
rect 32999 19876 33640 19904
rect 34532 19876 35900 19904
rect 32999 19873 33011 19876
rect 32953 19867 33011 19873
rect 32306 19796 32312 19848
rect 32364 19836 32370 19848
rect 32585 19839 32643 19845
rect 32585 19836 32597 19839
rect 32364 19808 32597 19836
rect 32364 19796 32370 19808
rect 32585 19805 32597 19808
rect 32631 19805 32643 19839
rect 32585 19799 32643 19805
rect 33042 19796 33048 19848
rect 33100 19836 33106 19848
rect 33612 19845 33640 19876
rect 35894 19864 35900 19876
rect 35952 19864 35958 19916
rect 43916 19904 43944 19932
rect 46934 19904 46940 19916
rect 43916 19876 45048 19904
rect 33413 19839 33471 19845
rect 33413 19836 33425 19839
rect 33100 19808 33425 19836
rect 33100 19796 33106 19808
rect 33413 19805 33425 19808
rect 33459 19805 33471 19839
rect 33413 19799 33471 19805
rect 33597 19839 33655 19845
rect 33597 19805 33609 19839
rect 33643 19805 33655 19839
rect 33597 19799 33655 19805
rect 33781 19839 33839 19845
rect 33781 19805 33793 19839
rect 33827 19836 33839 19839
rect 34885 19839 34943 19845
rect 34885 19836 34897 19839
rect 33827 19808 34897 19836
rect 33827 19805 33839 19808
rect 33781 19799 33839 19805
rect 34885 19805 34897 19808
rect 34931 19805 34943 19839
rect 34885 19799 34943 19805
rect 35437 19839 35495 19845
rect 35437 19805 35449 19839
rect 35483 19805 35495 19839
rect 35437 19799 35495 19805
rect 32214 19768 32220 19780
rect 32127 19740 32220 19768
rect 32214 19728 32220 19740
rect 32272 19768 32278 19780
rect 32769 19771 32827 19777
rect 32769 19768 32781 19771
rect 32272 19740 32781 19768
rect 32272 19728 32278 19740
rect 32769 19737 32781 19740
rect 32815 19768 32827 19771
rect 32950 19768 32956 19780
rect 32815 19740 32956 19768
rect 32815 19737 32827 19740
rect 32769 19731 32827 19737
rect 32950 19728 32956 19740
rect 33008 19728 33014 19780
rect 34698 19728 34704 19780
rect 34756 19768 34762 19780
rect 35452 19768 35480 19799
rect 43254 19796 43260 19848
rect 43312 19836 43318 19848
rect 43990 19836 43996 19848
rect 43312 19808 43996 19836
rect 43312 19796 43318 19808
rect 43990 19796 43996 19808
rect 44048 19796 44054 19848
rect 45020 19845 45048 19876
rect 45664 19876 46940 19904
rect 44085 19839 44143 19845
rect 44085 19805 44097 19839
rect 44131 19805 44143 19839
rect 44085 19799 44143 19805
rect 45005 19839 45063 19845
rect 45005 19805 45017 19839
rect 45051 19805 45063 19839
rect 45005 19799 45063 19805
rect 45189 19839 45247 19845
rect 45189 19805 45201 19839
rect 45235 19805 45247 19839
rect 45189 19799 45247 19805
rect 34756 19740 35480 19768
rect 35621 19771 35679 19777
rect 34756 19728 34762 19740
rect 35621 19737 35633 19771
rect 35667 19737 35679 19771
rect 35621 19731 35679 19737
rect 28552 19672 31754 19700
rect 35636 19700 35664 19731
rect 42702 19728 42708 19780
rect 42760 19768 42766 19780
rect 44100 19768 44128 19799
rect 42760 19740 44128 19768
rect 44269 19771 44327 19777
rect 42760 19728 42766 19740
rect 44269 19737 44281 19771
rect 44315 19768 44327 19771
rect 45204 19768 45232 19799
rect 44315 19740 45232 19768
rect 44315 19737 44327 19740
rect 44269 19731 44327 19737
rect 37366 19700 37372 19712
rect 35636 19672 37372 19700
rect 37366 19660 37372 19672
rect 37424 19700 37430 19712
rect 45664 19700 45692 19876
rect 46934 19864 46940 19876
rect 46992 19904 46998 19916
rect 47946 19904 47952 19916
rect 46992 19876 47952 19904
rect 46992 19864 46998 19876
rect 47946 19864 47952 19876
rect 48004 19864 48010 19916
rect 45830 19836 45836 19848
rect 45791 19808 45836 19836
rect 45830 19796 45836 19808
rect 45888 19796 45894 19848
rect 46106 19796 46112 19848
rect 46164 19836 46170 19848
rect 46569 19839 46627 19845
rect 46569 19836 46581 19839
rect 46164 19808 46581 19836
rect 46164 19796 46170 19808
rect 46569 19805 46581 19808
rect 46615 19805 46627 19839
rect 47394 19836 47400 19848
rect 47355 19808 47400 19836
rect 46569 19799 46627 19805
rect 47394 19796 47400 19808
rect 47452 19796 47458 19848
rect 45738 19728 45744 19780
rect 45796 19768 45802 19780
rect 46293 19771 46351 19777
rect 46293 19768 46305 19771
rect 45796 19740 46305 19768
rect 45796 19728 45802 19740
rect 46293 19737 46305 19740
rect 46339 19737 46351 19771
rect 46661 19771 46719 19777
rect 46661 19768 46673 19771
rect 46293 19731 46351 19737
rect 46400 19740 46673 19768
rect 37424 19672 45692 19700
rect 37424 19660 37430 19672
rect 45922 19660 45928 19712
rect 45980 19700 45986 19712
rect 46400 19700 46428 19740
rect 46661 19737 46673 19740
rect 46707 19768 46719 19771
rect 48038 19768 48044 19780
rect 46707 19740 48044 19768
rect 46707 19737 46719 19740
rect 46661 19731 46719 19737
rect 48038 19728 48044 19740
rect 48096 19728 48102 19780
rect 45980 19672 46428 19700
rect 46477 19703 46535 19709
rect 45980 19660 45986 19672
rect 46477 19669 46489 19703
rect 46523 19700 46535 19703
rect 46566 19700 46572 19712
rect 46523 19672 46572 19700
rect 46523 19669 46535 19672
rect 46477 19663 46535 19669
rect 46566 19660 46572 19672
rect 46624 19700 46630 19712
rect 46934 19700 46940 19712
rect 46624 19672 46940 19700
rect 46624 19660 46630 19672
rect 46934 19660 46940 19672
rect 46992 19660 46998 19712
rect 47486 19700 47492 19712
rect 47447 19672 47492 19700
rect 47486 19660 47492 19672
rect 47544 19660 47550 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 13357 19499 13415 19505
rect 13357 19465 13369 19499
rect 13403 19496 13415 19499
rect 14918 19496 14924 19508
rect 13403 19468 14924 19496
rect 13403 19465 13415 19468
rect 13357 19459 13415 19465
rect 14918 19456 14924 19468
rect 14976 19456 14982 19508
rect 20438 19496 20444 19508
rect 20399 19468 20444 19496
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 22830 19456 22836 19508
rect 22888 19496 22894 19508
rect 24486 19496 24492 19508
rect 22888 19468 24348 19496
rect 24447 19468 24492 19496
rect 22888 19456 22894 19468
rect 12894 19428 12900 19440
rect 12855 19400 12900 19428
rect 12894 19388 12900 19400
rect 12952 19388 12958 19440
rect 14366 19428 14372 19440
rect 14016 19400 14372 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 11514 19320 11520 19372
rect 11572 19360 11578 19372
rect 14016 19369 14044 19400
rect 14366 19388 14372 19400
rect 14424 19428 14430 19440
rect 15010 19428 15016 19440
rect 14424 19400 15016 19428
rect 14424 19388 14430 19400
rect 15010 19388 15016 19400
rect 15068 19388 15074 19440
rect 19797 19431 19855 19437
rect 19797 19428 19809 19431
rect 18998 19400 19809 19428
rect 19797 19397 19809 19400
rect 19843 19397 19855 19431
rect 19797 19391 19855 19397
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 11572 19332 12173 19360
rect 11572 19320 11578 19332
rect 12161 19329 12173 19332
rect 12207 19329 12219 19363
rect 12161 19323 12219 19329
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19329 14059 19363
rect 14182 19360 14188 19372
rect 14143 19332 14188 19360
rect 14001 19323 14059 19329
rect 14182 19320 14188 19332
rect 14240 19320 14246 19372
rect 14277 19363 14335 19369
rect 14277 19329 14289 19363
rect 14323 19360 14335 19363
rect 14734 19360 14740 19372
rect 14323 19332 14740 19360
rect 14323 19329 14335 19332
rect 14277 19323 14335 19329
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 14921 19363 14979 19369
rect 14921 19360 14933 19363
rect 14884 19332 14933 19360
rect 14884 19320 14890 19332
rect 14921 19329 14933 19332
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 19150 19320 19156 19372
rect 19208 19360 19214 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19208 19332 19717 19360
rect 19208 19320 19214 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 20349 19363 20407 19369
rect 20349 19329 20361 19363
rect 20395 19360 20407 19363
rect 20993 19363 21051 19369
rect 20993 19360 21005 19363
rect 20395 19332 21005 19360
rect 20395 19329 20407 19332
rect 20349 19323 20407 19329
rect 20993 19329 21005 19332
rect 21039 19360 21051 19363
rect 22646 19360 22652 19372
rect 21039 19332 22652 19360
rect 21039 19329 21051 19332
rect 20993 19323 21051 19329
rect 22646 19320 22652 19332
rect 22704 19320 22710 19372
rect 24118 19320 24124 19372
rect 24176 19320 24182 19372
rect 24320 19360 24348 19468
rect 24486 19456 24492 19468
rect 24544 19456 24550 19508
rect 28261 19499 28319 19505
rect 28261 19465 28273 19499
rect 28307 19465 28319 19499
rect 28902 19496 28908 19508
rect 28863 19468 28908 19496
rect 28261 19459 28319 19465
rect 28276 19428 28304 19459
rect 28902 19456 28908 19468
rect 28960 19456 28966 19508
rect 43898 19456 43904 19508
rect 43956 19496 43962 19508
rect 43993 19499 44051 19505
rect 43993 19496 44005 19499
rect 43956 19468 44005 19496
rect 43956 19456 43962 19468
rect 43993 19465 44005 19468
rect 44039 19465 44051 19499
rect 43993 19459 44051 19465
rect 46014 19456 46020 19508
rect 46072 19496 46078 19508
rect 47673 19499 47731 19505
rect 47673 19496 47685 19499
rect 46072 19468 47685 19496
rect 46072 19456 46078 19468
rect 47673 19465 47685 19468
rect 47719 19465 47731 19499
rect 47673 19459 47731 19465
rect 28994 19428 29000 19440
rect 28276 19400 29000 19428
rect 28994 19388 29000 19400
rect 29052 19428 29058 19440
rect 30282 19428 30288 19440
rect 29052 19400 30288 19428
rect 29052 19388 29058 19400
rect 30282 19388 30288 19400
rect 30340 19388 30346 19440
rect 33502 19428 33508 19440
rect 33463 19400 33508 19428
rect 33502 19388 33508 19400
rect 33560 19388 33566 19440
rect 36630 19388 36636 19440
rect 36688 19428 36694 19440
rect 36688 19400 47624 19428
rect 36688 19388 36694 19400
rect 28077 19363 28135 19369
rect 28077 19360 28089 19363
rect 24320 19332 28089 19360
rect 28077 19329 28089 19332
rect 28123 19329 28135 19363
rect 28077 19323 28135 19329
rect 28258 19320 28264 19372
rect 28316 19360 28322 19372
rect 28813 19363 28871 19369
rect 28813 19360 28825 19363
rect 28316 19332 28825 19360
rect 28316 19320 28322 19332
rect 28813 19329 28825 19332
rect 28859 19360 28871 19363
rect 28902 19360 28908 19372
rect 28859 19332 28908 19360
rect 28859 19329 28871 19332
rect 28813 19323 28871 19329
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 32493 19363 32551 19369
rect 32493 19329 32505 19363
rect 32539 19360 32551 19363
rect 33042 19360 33048 19372
rect 32539 19332 33048 19360
rect 32539 19329 32551 19332
rect 32493 19323 32551 19329
rect 33042 19320 33048 19332
rect 33100 19320 33106 19372
rect 33318 19360 33324 19372
rect 33279 19332 33324 19360
rect 33318 19320 33324 19332
rect 33376 19320 33382 19372
rect 35805 19363 35863 19369
rect 35805 19329 35817 19363
rect 35851 19360 35863 19363
rect 37090 19360 37096 19372
rect 35851 19332 37096 19360
rect 35851 19329 35863 19332
rect 35805 19323 35863 19329
rect 37090 19320 37096 19332
rect 37148 19320 37154 19372
rect 42702 19320 42708 19372
rect 42760 19360 42766 19372
rect 43901 19363 43959 19369
rect 43901 19360 43913 19363
rect 42760 19332 43913 19360
rect 42760 19320 42766 19332
rect 43901 19329 43913 19332
rect 43947 19329 43959 19363
rect 43901 19323 43959 19329
rect 43990 19320 43996 19372
rect 44048 19360 44054 19372
rect 44085 19363 44143 19369
rect 44085 19360 44097 19363
rect 44048 19332 44097 19360
rect 44048 19320 44054 19332
rect 44085 19329 44097 19332
rect 44131 19360 44143 19363
rect 45922 19360 45928 19372
rect 44131 19332 45784 19360
rect 45883 19332 45928 19360
rect 44131 19329 44143 19332
rect 44085 19323 44143 19329
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 13188 19264 14136 19292
rect 13188 19224 13216 19264
rect 6886 19196 13216 19224
rect 13265 19227 13323 19233
rect 3418 19116 3424 19168
rect 3476 19156 3482 19168
rect 6886 19156 6914 19196
rect 13265 19193 13277 19227
rect 13311 19224 13323 19227
rect 13817 19227 13875 19233
rect 13817 19224 13829 19227
rect 13311 19196 13829 19224
rect 13311 19193 13323 19196
rect 13265 19187 13323 19193
rect 13817 19193 13829 19196
rect 13863 19193 13875 19227
rect 14108 19224 14136 19264
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 17497 19295 17555 19301
rect 17497 19292 17509 19295
rect 17276 19264 17509 19292
rect 17276 19252 17282 19264
rect 17497 19261 17509 19264
rect 17543 19261 17555 19295
rect 17770 19292 17776 19304
rect 17731 19264 17776 19292
rect 17497 19255 17555 19261
rect 17770 19252 17776 19264
rect 17828 19252 17834 19304
rect 18230 19252 18236 19304
rect 18288 19292 18294 19304
rect 19245 19295 19303 19301
rect 19245 19292 19257 19295
rect 18288 19264 19257 19292
rect 18288 19252 18294 19264
rect 19245 19261 19257 19264
rect 19291 19261 19303 19295
rect 22738 19292 22744 19304
rect 22699 19264 22744 19292
rect 19245 19255 19303 19261
rect 22738 19252 22744 19264
rect 22796 19252 22802 19304
rect 23017 19295 23075 19301
rect 23017 19261 23029 19295
rect 23063 19292 23075 19295
rect 23658 19292 23664 19304
rect 23063 19264 23664 19292
rect 23063 19261 23075 19264
rect 23017 19255 23075 19261
rect 23658 19252 23664 19264
rect 23716 19252 23722 19304
rect 32582 19292 32588 19304
rect 32543 19264 32588 19292
rect 32582 19252 32588 19264
rect 32640 19252 32646 19304
rect 32861 19295 32919 19301
rect 32861 19261 32873 19295
rect 32907 19292 32919 19295
rect 33336 19292 33364 19320
rect 32907 19264 33364 19292
rect 33781 19295 33839 19301
rect 32907 19261 32919 19264
rect 32861 19255 32919 19261
rect 33781 19261 33793 19295
rect 33827 19261 33839 19295
rect 45756 19292 45784 19332
rect 45922 19320 45928 19332
rect 45980 19320 45986 19372
rect 46106 19320 46112 19372
rect 46164 19360 46170 19372
rect 46293 19363 46351 19369
rect 46293 19360 46305 19363
rect 46164 19332 46305 19360
rect 46164 19320 46170 19332
rect 46293 19329 46305 19332
rect 46339 19329 46351 19363
rect 46566 19360 46572 19372
rect 46527 19332 46572 19360
rect 46293 19323 46351 19329
rect 46566 19320 46572 19332
rect 46624 19320 46630 19372
rect 46658 19320 46664 19372
rect 46716 19320 46722 19372
rect 47596 19369 47624 19400
rect 46845 19363 46903 19369
rect 46845 19329 46857 19363
rect 46891 19329 46903 19363
rect 46845 19323 46903 19329
rect 47581 19363 47639 19369
rect 47581 19329 47593 19363
rect 47627 19329 47639 19363
rect 47581 19323 47639 19329
rect 46676 19292 46704 19320
rect 45756 19264 46704 19292
rect 33781 19255 33839 19261
rect 33796 19224 33824 19255
rect 14108 19196 17264 19224
rect 13817 19187 13875 19193
rect 3476 19128 6914 19156
rect 12345 19159 12403 19165
rect 3476 19116 3482 19128
rect 12345 19125 12357 19159
rect 12391 19156 12403 19159
rect 12802 19156 12808 19168
rect 12391 19128 12808 19156
rect 12391 19125 12403 19128
rect 12345 19119 12403 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 14826 19156 14832 19168
rect 13964 19128 14832 19156
rect 13964 19116 13970 19128
rect 14826 19116 14832 19128
rect 14884 19156 14890 19168
rect 15013 19159 15071 19165
rect 15013 19156 15025 19159
rect 14884 19128 15025 19156
rect 14884 19116 14890 19128
rect 15013 19125 15025 19128
rect 15059 19125 15071 19159
rect 17236 19156 17264 19196
rect 18800 19196 22094 19224
rect 18800 19156 18828 19196
rect 17236 19128 18828 19156
rect 15013 19119 15071 19125
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 21085 19159 21143 19165
rect 21085 19156 21097 19159
rect 20772 19128 21097 19156
rect 20772 19116 20778 19128
rect 21085 19125 21097 19128
rect 21131 19125 21143 19159
rect 22066 19156 22094 19196
rect 24136 19196 33824 19224
rect 24136 19156 24164 19196
rect 45738 19184 45744 19236
rect 45796 19224 45802 19236
rect 46860 19224 46888 19323
rect 45796 19196 46888 19224
rect 45796 19184 45802 19196
rect 35618 19156 35624 19168
rect 22066 19128 24164 19156
rect 35579 19128 35624 19156
rect 21085 19119 21143 19125
rect 35618 19116 35624 19128
rect 35676 19116 35682 19168
rect 45462 19156 45468 19168
rect 45423 19128 45468 19156
rect 45462 19116 45468 19128
rect 45520 19116 45526 19168
rect 46198 19156 46204 19168
rect 46159 19128 46204 19156
rect 46198 19116 46204 19128
rect 46256 19116 46262 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 2225 18915 2283 18921
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 18601 18955 18659 18961
rect 18601 18952 18613 18955
rect 17828 18924 18613 18952
rect 17828 18912 17834 18924
rect 18601 18921 18613 18924
rect 18647 18921 18659 18955
rect 23658 18952 23664 18964
rect 23619 18924 23664 18952
rect 18601 18915 18659 18921
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 30926 18912 30932 18964
rect 30984 18952 30990 18964
rect 31478 18952 31484 18964
rect 30984 18924 31484 18952
rect 30984 18912 30990 18924
rect 31478 18912 31484 18924
rect 31536 18912 31542 18964
rect 32582 18912 32588 18964
rect 32640 18952 32646 18964
rect 33505 18955 33563 18961
rect 33505 18952 33517 18955
rect 32640 18924 33517 18952
rect 32640 18912 32646 18924
rect 33505 18921 33517 18924
rect 33551 18921 33563 18955
rect 33505 18915 33563 18921
rect 6886 18856 22094 18884
rect 1578 18776 1584 18828
rect 1636 18816 1642 18828
rect 6886 18816 6914 18856
rect 1636 18788 6914 18816
rect 1636 18776 1642 18788
rect 15562 18776 15568 18828
rect 15620 18816 15626 18828
rect 15933 18819 15991 18825
rect 15933 18816 15945 18819
rect 15620 18788 15945 18816
rect 15620 18776 15626 18788
rect 15933 18785 15945 18788
rect 15979 18785 15991 18819
rect 17586 18816 17592 18828
rect 15933 18779 15991 18785
rect 17144 18788 17592 18816
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18748 2191 18751
rect 2314 18748 2320 18760
rect 2179 18720 2320 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 2314 18708 2320 18720
rect 2372 18748 2378 18760
rect 6546 18748 6552 18760
rect 2372 18720 6552 18748
rect 2372 18708 2378 18720
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 12802 18708 12808 18760
rect 12860 18748 12866 18760
rect 12989 18751 13047 18757
rect 12989 18748 13001 18751
rect 12860 18720 13001 18748
rect 12860 18708 12866 18720
rect 12989 18717 13001 18720
rect 13035 18717 13047 18751
rect 12989 18711 13047 18717
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 13872 18720 14105 18748
rect 13872 18708 13878 18720
rect 14093 18717 14105 18720
rect 14139 18717 14151 18751
rect 14918 18748 14924 18760
rect 14879 18720 14924 18748
rect 14093 18711 14151 18717
rect 14918 18708 14924 18720
rect 14976 18708 14982 18760
rect 15010 18708 15016 18760
rect 15068 18748 15074 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 15068 18720 15761 18748
rect 15068 18708 15074 18720
rect 15749 18717 15761 18720
rect 15795 18717 15807 18751
rect 15749 18711 15807 18717
rect 17144 18680 17172 18788
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 18104 18788 18153 18816
rect 18104 18776 18110 18788
rect 18141 18785 18153 18788
rect 18187 18785 18199 18819
rect 20714 18816 20720 18828
rect 20675 18788 20720 18816
rect 18141 18779 18199 18785
rect 20714 18776 20720 18788
rect 20772 18776 20778 18828
rect 22066 18816 22094 18856
rect 31110 18844 31116 18896
rect 31168 18884 31174 18896
rect 31662 18884 31668 18896
rect 31168 18856 31668 18884
rect 31168 18844 31174 18856
rect 31662 18844 31668 18856
rect 31720 18844 31726 18896
rect 32861 18887 32919 18893
rect 32861 18853 32873 18887
rect 32907 18884 32919 18887
rect 33042 18884 33048 18896
rect 32907 18856 33048 18884
rect 32907 18853 32919 18856
rect 32861 18847 32919 18853
rect 33042 18844 33048 18856
rect 33100 18844 33106 18896
rect 46106 18884 46112 18896
rect 37108 18856 46112 18884
rect 32309 18819 32367 18825
rect 22066 18788 32260 18816
rect 18230 18748 18236 18760
rect 18191 18720 18236 18748
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 20533 18751 20591 18757
rect 20533 18717 20545 18751
rect 20579 18717 20591 18751
rect 22830 18748 22836 18760
rect 22791 18720 22836 18748
rect 20533 18711 20591 18717
rect 6886 18652 17172 18680
rect 1578 18572 1584 18624
rect 1636 18612 1642 18624
rect 6886 18612 6914 18652
rect 17494 18640 17500 18692
rect 17552 18680 17558 18692
rect 17589 18683 17647 18689
rect 17589 18680 17601 18683
rect 17552 18652 17601 18680
rect 17552 18640 17558 18652
rect 17589 18649 17601 18652
rect 17635 18649 17647 18683
rect 20548 18680 20576 18711
rect 22830 18708 22836 18720
rect 22888 18708 22894 18760
rect 23566 18748 23572 18760
rect 23527 18720 23572 18748
rect 23566 18708 23572 18720
rect 23624 18708 23630 18760
rect 27246 18748 27252 18760
rect 27207 18720 27252 18748
rect 27246 18708 27252 18720
rect 27304 18708 27310 18760
rect 30926 18708 30932 18760
rect 30984 18748 30990 18760
rect 31021 18751 31079 18757
rect 31021 18748 31033 18751
rect 30984 18720 31033 18748
rect 30984 18708 30990 18720
rect 31021 18717 31033 18720
rect 31067 18717 31079 18751
rect 31021 18711 31079 18717
rect 31110 18708 31116 18760
rect 31168 18748 31174 18760
rect 31294 18748 31300 18760
rect 31168 18720 31213 18748
rect 31255 18720 31300 18748
rect 31168 18708 31174 18720
rect 31294 18708 31300 18720
rect 31352 18708 31358 18760
rect 31389 18751 31447 18757
rect 31389 18717 31401 18751
rect 31435 18717 31447 18751
rect 31389 18711 31447 18717
rect 22002 18680 22008 18692
rect 20548 18652 22008 18680
rect 17589 18643 17647 18649
rect 22002 18640 22008 18652
rect 22060 18640 22066 18692
rect 22373 18683 22431 18689
rect 22373 18649 22385 18683
rect 22419 18680 22431 18683
rect 22922 18680 22928 18692
rect 22419 18652 22928 18680
rect 22419 18649 22431 18652
rect 22373 18643 22431 18649
rect 22922 18640 22928 18652
rect 22980 18640 22986 18692
rect 27525 18683 27583 18689
rect 27525 18649 27537 18683
rect 27571 18680 27583 18683
rect 27706 18680 27712 18692
rect 27571 18652 27712 18680
rect 27571 18649 27583 18652
rect 27525 18643 27583 18649
rect 27706 18640 27712 18652
rect 27764 18640 27770 18692
rect 31404 18680 31432 18711
rect 31478 18708 31484 18760
rect 31536 18748 31542 18760
rect 32125 18751 32183 18757
rect 32125 18748 32137 18751
rect 31536 18720 32137 18748
rect 31536 18708 31542 18720
rect 32125 18717 32137 18720
rect 32171 18717 32183 18751
rect 32125 18711 32183 18717
rect 31404 18652 31616 18680
rect 1636 18584 6914 18612
rect 1636 18572 1642 18584
rect 13078 18572 13084 18624
rect 13136 18612 13142 18624
rect 13173 18615 13231 18621
rect 13173 18612 13185 18615
rect 13136 18584 13185 18612
rect 13136 18572 13142 18584
rect 13173 18581 13185 18584
rect 13219 18581 13231 18615
rect 13173 18575 13231 18581
rect 14090 18572 14096 18624
rect 14148 18612 14154 18624
rect 14185 18615 14243 18621
rect 14185 18612 14197 18615
rect 14148 18584 14197 18612
rect 14148 18572 14154 18584
rect 14185 18581 14197 18584
rect 14231 18581 14243 18615
rect 14734 18612 14740 18624
rect 14695 18584 14740 18612
rect 14185 18575 14243 18581
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 23014 18612 23020 18624
rect 22975 18584 23020 18612
rect 23014 18572 23020 18584
rect 23072 18572 23078 18624
rect 31202 18572 31208 18624
rect 31260 18612 31266 18624
rect 31389 18615 31447 18621
rect 31389 18612 31401 18615
rect 31260 18584 31401 18612
rect 31260 18572 31266 18584
rect 31389 18581 31401 18584
rect 31435 18581 31447 18615
rect 31588 18612 31616 18652
rect 31662 18640 31668 18692
rect 31720 18680 31726 18692
rect 31941 18683 31999 18689
rect 31941 18680 31953 18683
rect 31720 18652 31953 18680
rect 31720 18640 31726 18652
rect 31941 18649 31953 18652
rect 31987 18649 31999 18683
rect 32232 18680 32260 18788
rect 32309 18785 32321 18819
rect 32355 18816 32367 18819
rect 32355 18788 33456 18816
rect 32355 18785 32367 18788
rect 32309 18779 32367 18785
rect 32398 18708 32404 18760
rect 32456 18748 32462 18760
rect 32769 18751 32827 18757
rect 32769 18748 32781 18751
rect 32456 18720 32781 18748
rect 32456 18708 32462 18720
rect 32769 18717 32781 18720
rect 32815 18717 32827 18751
rect 32950 18748 32956 18760
rect 32911 18720 32956 18748
rect 32769 18711 32827 18717
rect 32950 18708 32956 18720
rect 33008 18708 33014 18760
rect 33428 18757 33456 18788
rect 33413 18751 33471 18757
rect 33413 18717 33425 18751
rect 33459 18717 33471 18751
rect 33594 18748 33600 18760
rect 33555 18720 33600 18748
rect 33413 18711 33471 18717
rect 33594 18708 33600 18720
rect 33652 18708 33658 18760
rect 37108 18757 37136 18856
rect 46106 18844 46112 18856
rect 46164 18844 46170 18896
rect 42613 18819 42671 18825
rect 42613 18785 42625 18819
rect 42659 18816 42671 18819
rect 43806 18816 43812 18828
rect 42659 18788 43812 18816
rect 42659 18785 42671 18788
rect 42613 18779 42671 18785
rect 43806 18776 43812 18788
rect 43864 18776 43870 18828
rect 45462 18776 45468 18828
rect 45520 18816 45526 18828
rect 46293 18819 46351 18825
rect 46293 18816 46305 18819
rect 45520 18788 46305 18816
rect 45520 18776 45526 18788
rect 46293 18785 46305 18788
rect 46339 18785 46351 18819
rect 46293 18779 46351 18785
rect 46477 18819 46535 18825
rect 46477 18785 46489 18819
rect 46523 18816 46535 18819
rect 47486 18816 47492 18828
rect 46523 18788 47492 18816
rect 46523 18785 46535 18788
rect 46477 18779 46535 18785
rect 47486 18776 47492 18788
rect 47544 18776 47550 18828
rect 48130 18816 48136 18828
rect 48091 18788 48136 18816
rect 48130 18776 48136 18788
rect 48188 18776 48194 18828
rect 37093 18751 37151 18757
rect 37093 18748 37105 18751
rect 36648 18720 37105 18748
rect 36648 18689 36676 18720
rect 37093 18717 37105 18720
rect 37139 18717 37151 18751
rect 37093 18711 37151 18717
rect 37185 18751 37243 18757
rect 37185 18717 37197 18751
rect 37231 18717 37243 18751
rect 37185 18711 37243 18717
rect 37277 18751 37335 18757
rect 37277 18717 37289 18751
rect 37323 18748 37335 18751
rect 37366 18748 37372 18760
rect 37323 18720 37372 18748
rect 37323 18717 37335 18720
rect 37277 18711 37335 18717
rect 36633 18683 36691 18689
rect 36633 18680 36645 18683
rect 32232 18652 36645 18680
rect 31941 18643 31999 18649
rect 36633 18649 36645 18652
rect 36679 18649 36691 18683
rect 36633 18643 36691 18649
rect 36906 18640 36912 18692
rect 36964 18680 36970 18692
rect 37200 18680 37228 18711
rect 37366 18708 37372 18720
rect 37424 18708 37430 18760
rect 45094 18748 45100 18760
rect 44284 18720 44588 18748
rect 45055 18720 45100 18748
rect 42794 18680 42800 18692
rect 36964 18652 41414 18680
rect 42755 18652 42800 18680
rect 36964 18640 36970 18652
rect 32306 18612 32312 18624
rect 31588 18584 32312 18612
rect 31389 18575 31447 18581
rect 32306 18572 32312 18584
rect 32364 18572 32370 18624
rect 37458 18612 37464 18624
rect 37419 18584 37464 18612
rect 37458 18572 37464 18584
rect 37516 18572 37522 18624
rect 41386 18612 41414 18652
rect 42794 18640 42800 18652
rect 42852 18640 42858 18692
rect 44284 18612 44312 18720
rect 44450 18680 44456 18692
rect 44411 18652 44456 18680
rect 44450 18640 44456 18652
rect 44508 18640 44514 18692
rect 44560 18680 44588 18720
rect 45094 18708 45100 18720
rect 45152 18708 45158 18760
rect 45281 18751 45339 18757
rect 45281 18717 45293 18751
rect 45327 18748 45339 18751
rect 45370 18748 45376 18760
rect 45327 18720 45376 18748
rect 45327 18717 45339 18720
rect 45281 18711 45339 18717
rect 45370 18708 45376 18720
rect 45428 18708 45434 18760
rect 45738 18680 45744 18692
rect 44560 18652 45744 18680
rect 45738 18640 45744 18652
rect 45796 18640 45802 18692
rect 41386 18584 44312 18612
rect 44358 18572 44364 18624
rect 44416 18612 44422 18624
rect 45189 18615 45247 18621
rect 45189 18612 45201 18615
rect 44416 18584 45201 18612
rect 44416 18572 44422 18584
rect 45189 18581 45201 18584
rect 45235 18581 45247 18615
rect 45189 18575 45247 18581
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 4614 18368 4620 18420
rect 4672 18408 4678 18420
rect 31294 18408 31300 18420
rect 4672 18380 30328 18408
rect 31255 18380 31300 18408
rect 4672 18368 4678 18380
rect 14090 18300 14096 18352
rect 14148 18300 14154 18352
rect 17218 18340 17224 18352
rect 17179 18312 17224 18340
rect 17218 18300 17224 18312
rect 17276 18300 17282 18352
rect 22554 18300 22560 18352
rect 22612 18300 22618 18352
rect 28810 18340 28816 18352
rect 24964 18312 28816 18340
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 13078 18272 13084 18284
rect 13039 18244 13084 18272
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 17126 18272 17132 18284
rect 17087 18244 17132 18272
rect 17126 18232 17132 18244
rect 17184 18232 17190 18284
rect 17865 18275 17923 18281
rect 17865 18241 17877 18275
rect 17911 18272 17923 18275
rect 17954 18272 17960 18284
rect 17911 18244 17960 18272
rect 17911 18241 17923 18244
rect 17865 18235 17923 18241
rect 17954 18232 17960 18244
rect 18012 18232 18018 18284
rect 18046 18232 18052 18284
rect 18104 18272 18110 18284
rect 21085 18275 21143 18281
rect 18104 18244 18149 18272
rect 18104 18232 18110 18244
rect 21085 18241 21097 18275
rect 21131 18241 21143 18275
rect 21085 18235 21143 18241
rect 13357 18207 13415 18213
rect 13357 18173 13369 18207
rect 13403 18204 13415 18207
rect 14734 18204 14740 18216
rect 13403 18176 14740 18204
rect 13403 18173 13415 18176
rect 13357 18167 13415 18173
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 14829 18207 14887 18213
rect 14829 18173 14841 18207
rect 14875 18204 14887 18207
rect 15010 18204 15016 18216
rect 14875 18176 15016 18204
rect 14875 18173 14887 18176
rect 14829 18167 14887 18173
rect 15010 18164 15016 18176
rect 15068 18164 15074 18216
rect 17862 18068 17868 18080
rect 17823 18040 17868 18068
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 21100 18068 21128 18235
rect 24762 18232 24768 18284
rect 24820 18272 24826 18284
rect 24964 18281 24992 18312
rect 28810 18300 28816 18312
rect 28868 18300 28874 18352
rect 30300 18340 30328 18380
rect 31294 18368 31300 18380
rect 31352 18368 31358 18420
rect 31389 18411 31447 18417
rect 31389 18377 31401 18411
rect 31435 18408 31447 18411
rect 31478 18408 31484 18420
rect 31435 18380 31484 18408
rect 31435 18377 31447 18380
rect 31389 18371 31447 18377
rect 31478 18368 31484 18380
rect 31536 18408 31542 18420
rect 37090 18408 37096 18420
rect 31536 18380 32996 18408
rect 37051 18380 37096 18408
rect 31536 18368 31542 18380
rect 30374 18340 30380 18352
rect 30300 18312 30380 18340
rect 24949 18275 25007 18281
rect 24949 18272 24961 18275
rect 24820 18244 24961 18272
rect 24820 18232 24826 18244
rect 24949 18241 24961 18244
rect 24995 18241 25007 18275
rect 24949 18235 25007 18241
rect 25774 18232 25780 18284
rect 25832 18272 25838 18284
rect 26145 18275 26203 18281
rect 26145 18272 26157 18275
rect 25832 18244 26157 18272
rect 25832 18232 25838 18244
rect 26145 18241 26157 18244
rect 26191 18241 26203 18275
rect 27154 18272 27160 18284
rect 27115 18244 27160 18272
rect 26145 18235 26203 18241
rect 27154 18232 27160 18244
rect 27212 18232 27218 18284
rect 27801 18275 27859 18281
rect 27801 18241 27813 18275
rect 27847 18241 27859 18275
rect 27801 18235 27859 18241
rect 28721 18275 28779 18281
rect 28721 18241 28733 18275
rect 28767 18272 28779 18275
rect 28994 18272 29000 18284
rect 28767 18244 29000 18272
rect 28767 18241 28779 18244
rect 28721 18235 28779 18241
rect 21177 18207 21235 18213
rect 21177 18173 21189 18207
rect 21223 18204 21235 18207
rect 21821 18207 21879 18213
rect 21821 18204 21833 18207
rect 21223 18176 21833 18204
rect 21223 18173 21235 18176
rect 21177 18167 21235 18173
rect 21821 18173 21833 18176
rect 21867 18173 21879 18207
rect 21821 18167 21879 18173
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 22152 18176 22197 18204
rect 22152 18164 22158 18176
rect 22462 18164 22468 18216
rect 22520 18204 22526 18216
rect 23566 18204 23572 18216
rect 22520 18176 23572 18204
rect 22520 18164 22526 18176
rect 23566 18164 23572 18176
rect 23624 18204 23630 18216
rect 26970 18204 26976 18216
rect 23624 18176 26372 18204
rect 26931 18176 26976 18204
rect 23624 18164 23630 18176
rect 26344 18145 26372 18176
rect 26970 18164 26976 18176
rect 27028 18164 27034 18216
rect 27246 18204 27252 18216
rect 27159 18176 27252 18204
rect 26329 18139 26387 18145
rect 26329 18105 26341 18139
rect 26375 18136 26387 18139
rect 27172 18136 27200 18176
rect 27246 18164 27252 18176
rect 27304 18204 27310 18216
rect 27816 18204 27844 18235
rect 28994 18232 29000 18244
rect 29052 18232 29058 18284
rect 30300 18281 30328 18312
rect 30374 18300 30380 18312
rect 30432 18300 30438 18352
rect 31202 18340 31208 18352
rect 31163 18312 31208 18340
rect 31202 18300 31208 18312
rect 31260 18300 31266 18352
rect 31496 18312 32352 18340
rect 30285 18275 30343 18281
rect 30285 18241 30297 18275
rect 30331 18241 30343 18275
rect 30285 18235 30343 18241
rect 30469 18275 30527 18281
rect 30469 18241 30481 18275
rect 30515 18272 30527 18275
rect 30650 18272 30656 18284
rect 30515 18244 30656 18272
rect 30515 18241 30527 18244
rect 30469 18235 30527 18241
rect 30650 18232 30656 18244
rect 30708 18232 30714 18284
rect 31220 18272 31248 18300
rect 31496 18272 31524 18312
rect 31220 18244 31524 18272
rect 31570 18232 31576 18284
rect 31628 18272 31634 18284
rect 32324 18281 32352 18312
rect 32968 18281 32996 18380
rect 37090 18368 37096 18380
rect 37148 18368 37154 18420
rect 37366 18408 37372 18420
rect 37292 18380 37372 18408
rect 34885 18343 34943 18349
rect 34885 18309 34897 18343
rect 34931 18340 34943 18343
rect 35618 18340 35624 18352
rect 34931 18312 35624 18340
rect 34931 18309 34943 18312
rect 34885 18303 34943 18309
rect 35618 18300 35624 18312
rect 35676 18300 35682 18352
rect 32309 18275 32367 18281
rect 31628 18244 31673 18272
rect 31628 18232 31634 18244
rect 32309 18241 32321 18275
rect 32355 18241 32367 18275
rect 32309 18235 32367 18241
rect 32953 18275 33011 18281
rect 32953 18241 32965 18275
rect 32999 18241 33011 18275
rect 32953 18235 33011 18241
rect 33318 18232 33324 18284
rect 33376 18272 33382 18284
rect 34701 18275 34759 18281
rect 34701 18272 34713 18275
rect 33376 18244 34713 18272
rect 33376 18232 33382 18244
rect 34701 18241 34713 18244
rect 34747 18241 34759 18275
rect 34701 18235 34759 18241
rect 36633 18275 36691 18281
rect 36633 18241 36645 18275
rect 36679 18272 36691 18275
rect 37292 18272 37320 18380
rect 37366 18368 37372 18380
rect 37424 18368 37430 18420
rect 42794 18408 42800 18420
rect 42755 18380 42800 18408
rect 42794 18368 42800 18380
rect 42852 18368 42858 18420
rect 45094 18368 45100 18420
rect 45152 18408 45158 18420
rect 47949 18411 48007 18417
rect 47949 18408 47961 18411
rect 45152 18380 47961 18408
rect 45152 18368 45158 18380
rect 47949 18377 47961 18380
rect 47995 18377 48007 18411
rect 47949 18371 48007 18377
rect 37458 18340 37464 18352
rect 37419 18312 37464 18340
rect 37458 18300 37464 18312
rect 37516 18300 37522 18352
rect 37550 18300 37556 18352
rect 37608 18340 37614 18352
rect 41782 18340 41788 18352
rect 37608 18312 41788 18340
rect 37608 18300 37614 18312
rect 41782 18300 41788 18312
rect 41840 18300 41846 18352
rect 45373 18343 45431 18349
rect 45373 18309 45385 18343
rect 45419 18340 45431 18343
rect 46198 18340 46204 18352
rect 45419 18312 46204 18340
rect 45419 18309 45431 18312
rect 45373 18303 45431 18309
rect 46198 18300 46204 18312
rect 46256 18300 46262 18352
rect 47026 18300 47032 18352
rect 47084 18340 47090 18352
rect 47765 18343 47823 18349
rect 47765 18340 47777 18343
rect 47084 18312 47777 18340
rect 47084 18300 47090 18312
rect 47765 18309 47777 18312
rect 47811 18309 47823 18343
rect 47765 18303 47823 18309
rect 44364 18284 44416 18290
rect 42705 18275 42763 18281
rect 42705 18272 42717 18275
rect 36679 18244 37320 18272
rect 39040 18244 42717 18272
rect 36679 18241 36691 18244
rect 36633 18235 36691 18241
rect 27304 18176 27844 18204
rect 27304 18164 27310 18176
rect 31294 18164 31300 18216
rect 31352 18204 31358 18216
rect 32125 18207 32183 18213
rect 32125 18204 32137 18207
rect 31352 18176 32137 18204
rect 31352 18164 31358 18176
rect 32125 18173 32137 18176
rect 32171 18204 32183 18207
rect 33594 18204 33600 18216
rect 32171 18176 33600 18204
rect 32171 18173 32183 18176
rect 32125 18167 32183 18173
rect 33594 18164 33600 18176
rect 33652 18164 33658 18216
rect 35894 18204 35900 18216
rect 35855 18176 35900 18204
rect 35894 18164 35900 18176
rect 35952 18204 35958 18216
rect 37182 18204 37188 18216
rect 35952 18176 37188 18204
rect 35952 18164 35958 18176
rect 37182 18164 37188 18176
rect 37240 18164 37246 18216
rect 37277 18207 37335 18213
rect 37277 18173 37289 18207
rect 37323 18173 37335 18207
rect 37277 18167 37335 18173
rect 26375 18108 27200 18136
rect 27341 18139 27399 18145
rect 26375 18105 26387 18108
rect 26329 18099 26387 18105
rect 27341 18105 27353 18139
rect 27387 18136 27399 18139
rect 27890 18136 27896 18148
rect 27387 18108 27896 18136
rect 27387 18105 27399 18108
rect 27341 18099 27399 18105
rect 27890 18096 27896 18108
rect 27948 18096 27954 18148
rect 31021 18139 31079 18145
rect 31021 18105 31033 18139
rect 31067 18136 31079 18139
rect 34790 18136 34796 18148
rect 31067 18108 34796 18136
rect 31067 18105 31079 18108
rect 31021 18099 31079 18105
rect 34790 18096 34796 18108
rect 34848 18096 34854 18148
rect 37090 18096 37096 18148
rect 37148 18136 37154 18148
rect 37292 18136 37320 18167
rect 37458 18164 37464 18216
rect 37516 18204 37522 18216
rect 37737 18207 37795 18213
rect 37737 18204 37749 18207
rect 37516 18176 37749 18204
rect 37516 18164 37522 18176
rect 37737 18173 37749 18176
rect 37783 18173 37795 18207
rect 37737 18167 37795 18173
rect 38378 18164 38384 18216
rect 38436 18204 38442 18216
rect 39040 18204 39068 18244
rect 42705 18241 42717 18244
rect 42751 18241 42763 18275
rect 42705 18235 42763 18241
rect 46750 18232 46756 18284
rect 46808 18272 46814 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 46808 18244 47593 18272
rect 46808 18232 46814 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47581 18235 47639 18241
rect 44364 18226 44416 18232
rect 43898 18204 43904 18216
rect 38436 18176 39068 18204
rect 41386 18176 43904 18204
rect 38436 18164 38442 18176
rect 37148 18108 37320 18136
rect 37148 18096 37154 18108
rect 22462 18068 22468 18080
rect 21100 18040 22468 18068
rect 22462 18028 22468 18040
rect 22520 18028 22526 18080
rect 22646 18028 22652 18080
rect 22704 18068 22710 18080
rect 23569 18071 23627 18077
rect 23569 18068 23581 18071
rect 22704 18040 23581 18068
rect 22704 18028 22710 18040
rect 23569 18037 23581 18040
rect 23615 18037 23627 18071
rect 23569 18031 23627 18037
rect 24765 18071 24823 18077
rect 24765 18037 24777 18071
rect 24811 18068 24823 18071
rect 24854 18068 24860 18080
rect 24811 18040 24860 18068
rect 24811 18037 24823 18040
rect 24765 18031 24823 18037
rect 24854 18028 24860 18040
rect 24912 18028 24918 18080
rect 27798 18068 27804 18080
rect 27759 18040 27804 18068
rect 27798 18028 27804 18040
rect 27856 18028 27862 18080
rect 28810 18068 28816 18080
rect 28771 18040 28816 18068
rect 28810 18028 28816 18040
rect 28868 18028 28874 18080
rect 30377 18071 30435 18077
rect 30377 18037 30389 18071
rect 30423 18068 30435 18071
rect 31478 18068 31484 18080
rect 30423 18040 31484 18068
rect 30423 18037 30435 18040
rect 30377 18031 30435 18037
rect 31478 18028 31484 18040
rect 31536 18028 31542 18080
rect 32306 18028 32312 18080
rect 32364 18068 32370 18080
rect 32493 18071 32551 18077
rect 32493 18068 32505 18071
rect 32364 18040 32505 18068
rect 32364 18028 32370 18040
rect 32493 18037 32505 18040
rect 32539 18037 32551 18071
rect 33042 18068 33048 18080
rect 33003 18040 33048 18068
rect 32493 18031 32551 18037
rect 33042 18028 33048 18040
rect 33100 18028 33106 18080
rect 36906 18068 36912 18080
rect 36867 18040 36912 18068
rect 36906 18028 36912 18040
rect 36964 18028 36970 18080
rect 37458 18028 37464 18080
rect 37516 18068 37522 18080
rect 41386 18068 41414 18176
rect 43898 18164 43904 18176
rect 43956 18164 43962 18216
rect 44726 18204 44732 18216
rect 44687 18176 44732 18204
rect 44726 18164 44732 18176
rect 44784 18204 44790 18216
rect 45189 18207 45247 18213
rect 45189 18204 45201 18207
rect 44784 18176 45201 18204
rect 44784 18164 44790 18176
rect 45189 18173 45201 18176
rect 45235 18173 45247 18207
rect 45189 18167 45247 18173
rect 45649 18207 45707 18213
rect 45649 18173 45661 18207
rect 45695 18173 45707 18207
rect 45649 18167 45707 18173
rect 41782 18096 41788 18148
rect 41840 18136 41846 18148
rect 45554 18136 45560 18148
rect 41840 18108 45560 18136
rect 41840 18096 41846 18108
rect 45554 18096 45560 18108
rect 45612 18136 45618 18148
rect 45664 18136 45692 18167
rect 45612 18108 45692 18136
rect 45612 18096 45618 18108
rect 37516 18040 41414 18068
rect 37516 18028 37522 18040
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 9766 17864 9772 17876
rect 3108 17836 9772 17864
rect 3108 17824 3114 17836
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 17034 17824 17040 17876
rect 17092 17864 17098 17876
rect 17405 17867 17463 17873
rect 17405 17864 17417 17867
rect 17092 17836 17417 17864
rect 17092 17824 17098 17836
rect 17405 17833 17417 17836
rect 17451 17833 17463 17867
rect 17405 17827 17463 17833
rect 17586 17824 17592 17876
rect 17644 17864 17650 17876
rect 18322 17864 18328 17876
rect 17644 17836 18328 17864
rect 17644 17824 17650 17836
rect 18322 17824 18328 17836
rect 18380 17824 18386 17876
rect 21177 17867 21235 17873
rect 21177 17833 21189 17867
rect 21223 17864 21235 17867
rect 22094 17864 22100 17876
rect 21223 17836 22100 17864
rect 21223 17833 21235 17836
rect 21177 17827 21235 17833
rect 22094 17824 22100 17836
rect 22152 17824 22158 17876
rect 22554 17864 22560 17876
rect 22515 17836 22560 17864
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 26142 17864 26148 17876
rect 25240 17836 26148 17864
rect 17770 17756 17776 17808
rect 17828 17796 17834 17808
rect 18230 17796 18236 17808
rect 17828 17768 18236 17796
rect 17828 17756 17834 17768
rect 18230 17756 18236 17768
rect 18288 17756 18294 17808
rect 22278 17796 22284 17808
rect 20916 17768 22284 17796
rect 20916 17737 20944 17768
rect 22278 17756 22284 17768
rect 22336 17756 22342 17808
rect 18417 17731 18475 17737
rect 18417 17728 18429 17731
rect 15764 17700 18429 17728
rect 12802 17660 12808 17672
rect 12763 17632 12808 17660
rect 12802 17620 12808 17632
rect 12860 17620 12866 17672
rect 13357 17663 13415 17669
rect 13357 17629 13369 17663
rect 13403 17660 13415 17663
rect 13814 17660 13820 17672
rect 13403 17632 13820 17660
rect 13403 17629 13415 17632
rect 13357 17623 13415 17629
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 14826 17620 14832 17672
rect 14884 17660 14890 17672
rect 15764 17669 15792 17700
rect 18417 17697 18429 17700
rect 18463 17697 18475 17731
rect 18417 17691 18475 17697
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17697 20959 17731
rect 22646 17728 22652 17740
rect 20901 17691 20959 17697
rect 22066 17700 22652 17728
rect 15473 17663 15531 17669
rect 15473 17660 15485 17663
rect 14884 17632 15485 17660
rect 14884 17620 14890 17632
rect 15473 17629 15485 17632
rect 15519 17629 15531 17663
rect 15473 17623 15531 17629
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17660 15991 17663
rect 16758 17660 16764 17672
rect 15979 17632 16764 17660
rect 15979 17629 15991 17632
rect 15933 17623 15991 17629
rect 15378 17552 15384 17604
rect 15436 17592 15442 17604
rect 15948 17592 15976 17623
rect 16758 17620 16764 17632
rect 16816 17660 16822 17672
rect 16853 17663 16911 17669
rect 16853 17660 16865 17663
rect 16816 17632 16865 17660
rect 16816 17620 16822 17632
rect 16853 17629 16865 17632
rect 16899 17629 16911 17663
rect 16853 17623 16911 17629
rect 17129 17663 17187 17669
rect 17129 17629 17141 17663
rect 17175 17660 17187 17663
rect 18141 17663 18199 17669
rect 17175 17632 18092 17660
rect 17175 17629 17187 17632
rect 17129 17623 17187 17629
rect 17144 17592 17172 17623
rect 15436 17564 15976 17592
rect 16868 17564 17172 17592
rect 17221 17595 17279 17601
rect 15436 17552 15442 17564
rect 16868 17536 16896 17564
rect 17221 17561 17233 17595
rect 17267 17592 17279 17595
rect 17586 17592 17592 17604
rect 17267 17564 17592 17592
rect 17267 17561 17279 17564
rect 17221 17555 17279 17561
rect 17586 17552 17592 17564
rect 17644 17552 17650 17604
rect 17770 17552 17776 17604
rect 17828 17592 17834 17604
rect 18064 17601 18092 17632
rect 18141 17629 18153 17663
rect 18187 17660 18199 17663
rect 18322 17660 18328 17672
rect 18187 17632 18328 17660
rect 18187 17629 18199 17632
rect 18141 17623 18199 17629
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 20530 17620 20536 17672
rect 20588 17660 20594 17672
rect 20809 17663 20867 17669
rect 20809 17660 20821 17663
rect 20588 17632 20821 17660
rect 20588 17620 20594 17632
rect 20809 17629 20821 17632
rect 20855 17660 20867 17663
rect 22066 17660 22094 17700
rect 22646 17688 22652 17700
rect 22704 17688 22710 17740
rect 24854 17688 24860 17740
rect 24912 17728 24918 17740
rect 25240 17737 25268 17836
rect 26142 17824 26148 17836
rect 26200 17864 26206 17876
rect 26605 17867 26663 17873
rect 26200 17836 26464 17864
rect 26200 17824 26206 17836
rect 25225 17731 25283 17737
rect 25225 17728 25237 17731
rect 24912 17700 25237 17728
rect 24912 17688 24918 17700
rect 25225 17697 25237 17700
rect 25271 17697 25283 17731
rect 25225 17691 25283 17697
rect 25409 17731 25467 17737
rect 25409 17697 25421 17731
rect 25455 17728 25467 17731
rect 25590 17728 25596 17740
rect 25455 17700 25596 17728
rect 25455 17697 25467 17700
rect 25409 17691 25467 17697
rect 25590 17688 25596 17700
rect 25648 17688 25654 17740
rect 20855 17632 22094 17660
rect 22465 17663 22523 17669
rect 20855 17629 20867 17632
rect 20809 17623 20867 17629
rect 22465 17629 22477 17663
rect 22511 17660 22523 17663
rect 23014 17660 23020 17672
rect 22511 17632 23020 17660
rect 22511 17629 22523 17632
rect 22465 17623 22523 17629
rect 23014 17620 23020 17632
rect 23072 17660 23078 17672
rect 23382 17660 23388 17672
rect 23072 17632 23388 17660
rect 23072 17620 23078 17632
rect 23382 17620 23388 17632
rect 23440 17620 23446 17672
rect 23566 17660 23572 17672
rect 23527 17632 23572 17660
rect 23566 17620 23572 17632
rect 23624 17620 23630 17672
rect 26436 17669 26464 17836
rect 26605 17833 26617 17867
rect 26651 17864 26663 17867
rect 27154 17864 27160 17876
rect 26651 17836 27160 17864
rect 26651 17833 26663 17836
rect 26605 17827 26663 17833
rect 27154 17824 27160 17836
rect 27212 17824 27218 17876
rect 28718 17824 28724 17876
rect 28776 17864 28782 17876
rect 28905 17867 28963 17873
rect 28905 17864 28917 17867
rect 28776 17836 28917 17864
rect 28776 17824 28782 17836
rect 28905 17833 28917 17836
rect 28951 17833 28963 17867
rect 28905 17827 28963 17833
rect 31205 17867 31263 17873
rect 31205 17833 31217 17867
rect 31251 17864 31263 17867
rect 31294 17864 31300 17876
rect 31251 17836 31300 17864
rect 31251 17833 31263 17836
rect 31205 17827 31263 17833
rect 31294 17824 31300 17836
rect 31352 17824 31358 17876
rect 34790 17824 34796 17876
rect 34848 17864 34854 17876
rect 37458 17864 37464 17876
rect 34848 17836 37464 17864
rect 34848 17824 34854 17836
rect 37458 17824 37464 17836
rect 37516 17824 37522 17876
rect 44266 17824 44272 17876
rect 44324 17864 44330 17876
rect 45649 17867 45707 17873
rect 45649 17864 45661 17867
rect 44324 17836 45661 17864
rect 44324 17824 44330 17836
rect 45649 17833 45661 17836
rect 45695 17833 45707 17867
rect 45649 17827 45707 17833
rect 35434 17756 35440 17808
rect 35492 17796 35498 17808
rect 44174 17796 44180 17808
rect 35492 17768 44180 17796
rect 35492 17756 35498 17768
rect 44174 17756 44180 17768
rect 44232 17756 44238 17808
rect 27157 17731 27215 17737
rect 27157 17697 27169 17731
rect 27203 17728 27215 17731
rect 27798 17728 27804 17740
rect 27203 17700 27804 17728
rect 27203 17697 27215 17700
rect 27157 17691 27215 17697
rect 27798 17688 27804 17700
rect 27856 17688 27862 17740
rect 30469 17731 30527 17737
rect 30469 17697 30481 17731
rect 30515 17728 30527 17731
rect 31570 17728 31576 17740
rect 30515 17700 31576 17728
rect 30515 17697 30527 17700
rect 30469 17691 30527 17697
rect 31570 17688 31576 17700
rect 31628 17688 31634 17740
rect 32953 17731 33011 17737
rect 32953 17697 32965 17731
rect 32999 17728 33011 17731
rect 37090 17728 37096 17740
rect 32999 17700 37096 17728
rect 32999 17697 33011 17700
rect 32953 17691 33011 17697
rect 37090 17688 37096 17700
rect 37148 17688 37154 17740
rect 43898 17688 43904 17740
rect 43956 17728 43962 17740
rect 45465 17731 45523 17737
rect 45465 17728 45477 17731
rect 43956 17700 45477 17728
rect 43956 17688 43962 17700
rect 45465 17697 45477 17700
rect 45511 17697 45523 17731
rect 45465 17691 45523 17697
rect 46293 17731 46351 17737
rect 46293 17697 46305 17731
rect 46339 17728 46351 17731
rect 47486 17728 47492 17740
rect 46339 17700 47492 17728
rect 46339 17697 46351 17700
rect 46293 17691 46351 17697
rect 47486 17688 47492 17700
rect 47544 17688 47550 17740
rect 25133 17663 25191 17669
rect 25133 17629 25145 17663
rect 25179 17629 25191 17663
rect 25133 17623 25191 17629
rect 25317 17663 25375 17669
rect 25317 17629 25329 17663
rect 25363 17660 25375 17663
rect 26421 17663 26479 17669
rect 25363 17632 26372 17660
rect 25363 17629 25375 17632
rect 25317 17623 25375 17629
rect 17865 17595 17923 17601
rect 17865 17592 17877 17595
rect 17828 17564 17877 17592
rect 17828 17552 17834 17564
rect 17865 17561 17877 17564
rect 17911 17561 17923 17595
rect 17865 17555 17923 17561
rect 18049 17595 18107 17601
rect 18049 17561 18061 17595
rect 18095 17592 18107 17595
rect 19242 17592 19248 17604
rect 18095 17564 19248 17592
rect 18095 17561 18107 17564
rect 18049 17555 18107 17561
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 12805 17527 12863 17533
rect 12805 17524 12817 17527
rect 12676 17496 12817 17524
rect 12676 17484 12682 17496
rect 12805 17493 12817 17496
rect 12851 17493 12863 17527
rect 13446 17524 13452 17536
rect 13407 17496 13452 17524
rect 12805 17487 12863 17493
rect 13446 17484 13452 17496
rect 13504 17484 13510 17536
rect 15286 17524 15292 17536
rect 15247 17496 15292 17524
rect 15286 17484 15292 17496
rect 15344 17484 15350 17536
rect 16850 17484 16856 17536
rect 16908 17484 16914 17536
rect 17037 17527 17095 17533
rect 17037 17493 17049 17527
rect 17083 17524 17095 17527
rect 17880 17524 17908 17555
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 25148 17592 25176 17623
rect 25866 17592 25872 17604
rect 25148 17564 25872 17592
rect 25424 17536 25452 17564
rect 25866 17552 25872 17564
rect 25924 17592 25930 17604
rect 26237 17595 26295 17601
rect 26237 17592 26249 17595
rect 25924 17564 26249 17592
rect 25924 17552 25930 17564
rect 26237 17561 26249 17564
rect 26283 17561 26295 17595
rect 26344 17592 26372 17632
rect 26421 17629 26433 17663
rect 26467 17629 26479 17663
rect 26421 17623 26479 17629
rect 28994 17620 29000 17672
rect 29052 17660 29058 17672
rect 29549 17663 29607 17669
rect 29549 17660 29561 17663
rect 29052 17632 29561 17660
rect 29052 17620 29058 17632
rect 29549 17629 29561 17632
rect 29595 17629 29607 17663
rect 30374 17660 30380 17672
rect 30335 17632 30380 17660
rect 29549 17623 29607 17629
rect 30374 17620 30380 17632
rect 30432 17620 30438 17672
rect 30561 17663 30619 17669
rect 30561 17629 30573 17663
rect 30607 17660 30619 17663
rect 30650 17660 30656 17672
rect 30607 17632 30656 17660
rect 30607 17629 30619 17632
rect 30561 17623 30619 17629
rect 30650 17620 30656 17632
rect 30708 17620 30714 17672
rect 31110 17660 31116 17672
rect 31071 17632 31116 17660
rect 31110 17620 31116 17632
rect 31168 17620 31174 17672
rect 31294 17660 31300 17672
rect 31255 17632 31300 17660
rect 31294 17620 31300 17632
rect 31352 17620 31358 17672
rect 31478 17620 31484 17672
rect 31536 17660 31542 17672
rect 31941 17663 31999 17669
rect 31941 17660 31953 17663
rect 31536 17632 31953 17660
rect 31536 17620 31542 17632
rect 31941 17629 31953 17632
rect 31987 17629 31999 17663
rect 32306 17660 32312 17672
rect 32267 17632 32312 17660
rect 31941 17623 31999 17629
rect 32306 17620 32312 17632
rect 32364 17620 32370 17672
rect 32858 17620 32864 17672
rect 32916 17660 32922 17672
rect 35434 17660 35440 17672
rect 32916 17632 35440 17660
rect 32916 17620 32922 17632
rect 35434 17620 35440 17632
rect 35492 17620 35498 17672
rect 36170 17660 36176 17672
rect 36131 17632 36176 17660
rect 36170 17620 36176 17632
rect 36228 17620 36234 17672
rect 45005 17663 45063 17669
rect 45005 17629 45017 17663
rect 45051 17660 45063 17663
rect 45094 17660 45100 17672
rect 45051 17632 45100 17660
rect 45051 17629 45063 17632
rect 45005 17623 45063 17629
rect 45094 17620 45100 17632
rect 45152 17620 45158 17672
rect 45370 17660 45376 17672
rect 45331 17632 45376 17660
rect 45370 17620 45376 17632
rect 45428 17620 45434 17672
rect 26786 17592 26792 17604
rect 26344 17564 26792 17592
rect 26237 17555 26295 17561
rect 26786 17552 26792 17564
rect 26844 17552 26850 17604
rect 27433 17595 27491 17601
rect 27433 17561 27445 17595
rect 27479 17561 27491 17595
rect 28810 17592 28816 17604
rect 28658 17564 28816 17592
rect 27433 17555 27491 17561
rect 17083 17496 17908 17524
rect 17083 17493 17095 17496
rect 17037 17487 17095 17493
rect 18230 17484 18236 17536
rect 18288 17524 18294 17536
rect 23753 17527 23811 17533
rect 18288 17496 18333 17524
rect 18288 17484 18294 17496
rect 23753 17493 23765 17527
rect 23799 17524 23811 17527
rect 24118 17524 24124 17536
rect 23799 17496 24124 17524
rect 23799 17493 23811 17496
rect 23753 17487 23811 17493
rect 24118 17484 24124 17496
rect 24176 17484 24182 17536
rect 24946 17524 24952 17536
rect 24907 17496 24952 17524
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 25406 17484 25412 17536
rect 25464 17484 25470 17536
rect 27448 17524 27476 17555
rect 28810 17552 28816 17564
rect 28868 17552 28874 17604
rect 30926 17552 30932 17604
rect 30984 17592 30990 17604
rect 31312 17592 31340 17620
rect 30984 17564 31340 17592
rect 35529 17595 35587 17601
rect 30984 17552 30990 17564
rect 35529 17561 35541 17595
rect 35575 17592 35587 17595
rect 36357 17595 36415 17601
rect 36357 17592 36369 17595
rect 35575 17564 36369 17592
rect 35575 17561 35587 17564
rect 35529 17555 35587 17561
rect 36357 17561 36369 17564
rect 36403 17561 36415 17595
rect 36357 17555 36415 17561
rect 38013 17595 38071 17601
rect 38013 17561 38025 17595
rect 38059 17592 38071 17595
rect 46290 17592 46296 17604
rect 38059 17564 46296 17592
rect 38059 17561 38071 17564
rect 38013 17555 38071 17561
rect 46290 17552 46296 17564
rect 46348 17552 46354 17604
rect 46477 17595 46535 17601
rect 46477 17561 46489 17595
rect 46523 17592 46535 17595
rect 46934 17592 46940 17604
rect 46523 17564 46940 17592
rect 46523 17561 46535 17564
rect 46477 17555 46535 17561
rect 46934 17552 46940 17564
rect 46992 17552 46998 17604
rect 48130 17592 48136 17604
rect 48091 17564 48136 17592
rect 48130 17552 48136 17564
rect 48188 17552 48194 17604
rect 27614 17524 27620 17536
rect 27448 17496 27620 17524
rect 27614 17484 27620 17496
rect 27672 17484 27678 17536
rect 29638 17524 29644 17536
rect 29599 17496 29644 17524
rect 29638 17484 29644 17496
rect 29696 17484 29702 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 17129 17323 17187 17329
rect 17129 17289 17141 17323
rect 17175 17320 17187 17323
rect 18046 17320 18052 17332
rect 17175 17292 18052 17320
rect 17175 17289 17187 17292
rect 17129 17283 17187 17289
rect 18046 17280 18052 17292
rect 18104 17280 18110 17332
rect 22925 17323 22983 17329
rect 22925 17289 22937 17323
rect 22971 17320 22983 17323
rect 24762 17320 24768 17332
rect 22971 17292 24768 17320
rect 22971 17289 22983 17292
rect 22925 17283 22983 17289
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 26970 17280 26976 17332
rect 27028 17320 27034 17332
rect 27065 17323 27123 17329
rect 27065 17320 27077 17323
rect 27028 17292 27077 17320
rect 27028 17280 27034 17292
rect 27065 17289 27077 17292
rect 27111 17289 27123 17323
rect 27065 17283 27123 17289
rect 27706 17280 27712 17332
rect 27764 17280 27770 17332
rect 31478 17320 31484 17332
rect 31439 17292 31484 17320
rect 31478 17280 31484 17292
rect 31536 17280 31542 17332
rect 45370 17280 45376 17332
rect 45428 17320 45434 17332
rect 46293 17323 46351 17329
rect 46293 17320 46305 17323
rect 45428 17292 46305 17320
rect 45428 17280 45434 17292
rect 46293 17289 46305 17292
rect 46339 17289 46351 17323
rect 46934 17320 46940 17332
rect 46895 17292 46940 17320
rect 46293 17283 46351 17289
rect 46934 17280 46940 17292
rect 46992 17280 46998 17332
rect 12618 17252 12624 17264
rect 12452 17224 12624 17252
rect 12452 17193 12480 17224
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 13446 17212 13452 17264
rect 13504 17212 13510 17264
rect 16761 17255 16819 17261
rect 16761 17221 16773 17255
rect 16807 17252 16819 17255
rect 16850 17252 16856 17264
rect 16807 17224 16856 17252
rect 16807 17221 16819 17224
rect 16761 17215 16819 17221
rect 16850 17212 16856 17224
rect 16908 17212 16914 17264
rect 16977 17255 17035 17261
rect 16977 17221 16989 17255
rect 17023 17252 17035 17255
rect 17862 17252 17868 17264
rect 17023 17224 17356 17252
rect 17823 17224 17868 17252
rect 17023 17221 17035 17224
rect 16977 17215 17035 17221
rect 12437 17187 12495 17193
rect 12437 17153 12449 17187
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17184 15991 17187
rect 15979 17156 17264 17184
rect 15979 17153 15991 17156
rect 15933 17147 15991 17153
rect 12710 17116 12716 17128
rect 12671 17088 12716 17116
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 12802 17076 12808 17128
rect 12860 17116 12866 17128
rect 15120 17116 15148 17147
rect 17126 17116 17132 17128
rect 12860 17088 17132 17116
rect 12860 17076 12866 17088
rect 17126 17076 17132 17088
rect 17184 17076 17190 17128
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 1452 16952 2053 16980
rect 1452 16940 1458 16952
rect 2041 16949 2053 16952
rect 2087 16949 2099 16983
rect 2041 16943 2099 16949
rect 13354 16940 13360 16992
rect 13412 16980 13418 16992
rect 14182 16980 14188 16992
rect 13412 16952 14188 16980
rect 13412 16940 13418 16952
rect 14182 16940 14188 16952
rect 14240 16940 14246 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 15105 16983 15163 16989
rect 15105 16980 15117 16983
rect 15068 16952 15117 16980
rect 15068 16940 15074 16952
rect 15105 16949 15117 16952
rect 15151 16949 15163 16983
rect 16022 16980 16028 16992
rect 15983 16952 16028 16980
rect 15105 16943 15163 16949
rect 16022 16940 16028 16952
rect 16080 16940 16086 16992
rect 16945 16983 17003 16989
rect 16945 16949 16957 16983
rect 16991 16980 17003 16983
rect 17034 16980 17040 16992
rect 16991 16952 17040 16980
rect 16991 16949 17003 16952
rect 16945 16943 17003 16949
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 17236 16980 17264 17156
rect 17328 17048 17356 17224
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 18874 17212 18880 17264
rect 18932 17212 18938 17264
rect 21821 17255 21879 17261
rect 21821 17221 21833 17255
rect 21867 17252 21879 17255
rect 22186 17252 22192 17264
rect 21867 17224 22192 17252
rect 21867 17221 21879 17224
rect 21821 17215 21879 17221
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 23106 17252 23112 17264
rect 23067 17224 23112 17252
rect 23106 17212 23112 17224
rect 23164 17212 23170 17264
rect 26142 17212 26148 17264
rect 26200 17252 26206 17264
rect 27724 17252 27752 17280
rect 29638 17252 29644 17264
rect 26200 17224 27200 17252
rect 26200 17212 26206 17224
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22097 17187 22155 17193
rect 22097 17153 22109 17187
rect 22143 17184 22155 17187
rect 22278 17184 22284 17196
rect 22143 17156 22284 17184
rect 22143 17153 22155 17156
rect 22097 17147 22155 17153
rect 17402 17076 17408 17128
rect 17460 17116 17466 17128
rect 17589 17119 17647 17125
rect 17589 17116 17601 17119
rect 17460 17088 17601 17116
rect 17460 17076 17466 17088
rect 17589 17085 17601 17088
rect 17635 17085 17647 17119
rect 18230 17116 18236 17128
rect 17589 17079 17647 17085
rect 17696 17088 18236 17116
rect 17696 17048 17724 17088
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 22020 17116 22048 17147
rect 22278 17144 22284 17156
rect 22336 17184 22342 17196
rect 22336 17156 22876 17184
rect 22336 17144 22342 17156
rect 22646 17116 22652 17128
rect 22020 17088 22652 17116
rect 22646 17076 22652 17088
rect 22704 17076 22710 17128
rect 22848 17116 22876 17156
rect 23014 17144 23020 17196
rect 23072 17184 23078 17196
rect 24118 17184 24124 17196
rect 23072 17156 23117 17184
rect 24079 17156 24124 17184
rect 23072 17144 23078 17156
rect 24118 17144 24124 17156
rect 24176 17144 24182 17196
rect 25498 17144 25504 17196
rect 25556 17144 25562 17196
rect 25866 17144 25872 17196
rect 25924 17184 25930 17196
rect 27172 17193 27200 17224
rect 27632 17224 27752 17252
rect 29118 17224 29644 17252
rect 27632 17193 27660 17224
rect 29638 17212 29644 17224
rect 29696 17212 29702 17264
rect 47026 17252 47032 17264
rect 46400 17224 47032 17252
rect 26973 17187 27031 17193
rect 26973 17184 26985 17187
rect 25924 17156 26985 17184
rect 25924 17144 25930 17156
rect 26973 17153 26985 17156
rect 27019 17153 27031 17187
rect 26973 17147 27031 17153
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 27617 17187 27675 17193
rect 27617 17153 27629 17187
rect 27663 17153 27675 17187
rect 27617 17147 27675 17153
rect 31389 17187 31447 17193
rect 31389 17153 31401 17187
rect 31435 17184 31447 17187
rect 31478 17184 31484 17196
rect 31435 17156 31484 17184
rect 31435 17153 31447 17156
rect 31389 17147 31447 17153
rect 31478 17144 31484 17156
rect 31536 17144 31542 17196
rect 31573 17187 31631 17193
rect 31573 17153 31585 17187
rect 31619 17184 31631 17187
rect 33042 17184 33048 17196
rect 31619 17156 33048 17184
rect 31619 17153 31631 17156
rect 31573 17147 31631 17153
rect 33042 17144 33048 17156
rect 33100 17144 33106 17196
rect 37090 17144 37096 17196
rect 37148 17184 37154 17196
rect 46400 17193 46428 17224
rect 47026 17212 47032 17224
rect 47084 17212 47090 17264
rect 47118 17212 47124 17264
rect 47176 17252 47182 17264
rect 47176 17224 47348 17252
rect 47176 17212 47182 17224
rect 43717 17187 43775 17193
rect 43717 17184 43729 17187
rect 37148 17156 43729 17184
rect 37148 17144 37154 17156
rect 43717 17153 43729 17156
rect 43763 17153 43775 17187
rect 43717 17147 43775 17153
rect 46201 17187 46259 17193
rect 46201 17153 46213 17187
rect 46247 17153 46259 17187
rect 46201 17147 46259 17153
rect 46385 17187 46443 17193
rect 46385 17153 46397 17187
rect 46431 17153 46443 17187
rect 46385 17147 46443 17153
rect 46845 17187 46903 17193
rect 46845 17153 46857 17187
rect 46891 17184 46903 17187
rect 47210 17184 47216 17196
rect 46891 17156 47216 17184
rect 46891 17153 46903 17156
rect 46845 17147 46903 17153
rect 24026 17116 24032 17128
rect 22848 17088 24032 17116
rect 24026 17076 24032 17088
rect 24084 17076 24090 17128
rect 24397 17119 24455 17125
rect 24397 17085 24409 17119
rect 24443 17116 24455 17119
rect 25130 17116 25136 17128
rect 24443 17088 25136 17116
rect 24443 17085 24455 17088
rect 24397 17079 24455 17085
rect 25130 17076 25136 17088
rect 25188 17076 25194 17128
rect 27062 17076 27068 17128
rect 27120 17116 27126 17128
rect 27893 17119 27951 17125
rect 27893 17116 27905 17119
rect 27120 17088 27905 17116
rect 27120 17076 27126 17088
rect 27893 17085 27905 17088
rect 27939 17085 27951 17119
rect 27893 17079 27951 17085
rect 29641 17119 29699 17125
rect 29641 17085 29653 17119
rect 29687 17116 29699 17119
rect 36170 17116 36176 17128
rect 29687 17088 36176 17116
rect 29687 17085 29699 17088
rect 29641 17079 29699 17085
rect 17328 17020 17724 17048
rect 22462 17008 22468 17060
rect 22520 17048 22526 17060
rect 22741 17051 22799 17057
rect 22741 17048 22753 17051
rect 22520 17020 22753 17048
rect 22520 17008 22526 17020
rect 22741 17017 22753 17020
rect 22787 17048 22799 17051
rect 23198 17048 23204 17060
rect 22787 17020 23204 17048
rect 22787 17017 22799 17020
rect 22741 17011 22799 17017
rect 23198 17008 23204 17020
rect 23256 17008 23262 17060
rect 19150 16980 19156 16992
rect 17236 16952 19156 16980
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 19242 16940 19248 16992
rect 19300 16980 19306 16992
rect 19337 16983 19395 16989
rect 19337 16980 19349 16983
rect 19300 16952 19349 16980
rect 19300 16940 19306 16952
rect 19337 16949 19349 16952
rect 19383 16949 19395 16983
rect 19337 16943 19395 16949
rect 20990 16940 20996 16992
rect 21048 16980 21054 16992
rect 21821 16983 21879 16989
rect 21821 16980 21833 16983
rect 21048 16952 21833 16980
rect 21048 16940 21054 16952
rect 21821 16949 21833 16952
rect 21867 16949 21879 16983
rect 21821 16943 21879 16949
rect 21910 16940 21916 16992
rect 21968 16980 21974 16992
rect 23293 16983 23351 16989
rect 23293 16980 23305 16983
rect 21968 16952 23305 16980
rect 21968 16940 21974 16952
rect 23293 16949 23305 16952
rect 23339 16949 23351 16983
rect 23293 16943 23351 16949
rect 23934 16940 23940 16992
rect 23992 16980 23998 16992
rect 25590 16980 25596 16992
rect 23992 16952 25596 16980
rect 23992 16940 23998 16952
rect 25590 16940 25596 16952
rect 25648 16980 25654 16992
rect 25869 16983 25927 16989
rect 25869 16980 25881 16983
rect 25648 16952 25881 16980
rect 25648 16940 25654 16952
rect 25869 16949 25881 16952
rect 25915 16949 25927 16983
rect 25869 16943 25927 16949
rect 26786 16940 26792 16992
rect 26844 16980 26850 16992
rect 29656 16980 29684 17079
rect 36170 17076 36176 17088
rect 36228 17076 36234 17128
rect 43898 17116 43904 17128
rect 43859 17088 43904 17116
rect 43898 17076 43904 17088
rect 43956 17076 43962 17128
rect 45370 17116 45376 17128
rect 45331 17088 45376 17116
rect 45370 17076 45376 17088
rect 45428 17076 45434 17128
rect 46216 17116 46244 17147
rect 47210 17144 47216 17156
rect 47268 17144 47274 17196
rect 47320 17184 47348 17224
rect 47581 17187 47639 17193
rect 47581 17184 47593 17187
rect 47320 17156 47593 17184
rect 47581 17153 47593 17156
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 46750 17116 46756 17128
rect 46216 17088 46756 17116
rect 46750 17076 46756 17088
rect 46808 17076 46814 17128
rect 47670 16980 47676 16992
rect 26844 16952 29684 16980
rect 47631 16952 47676 16980
rect 26844 16940 26850 16952
rect 47670 16940 47676 16952
rect 47728 16940 47734 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 12710 16736 12716 16788
rect 12768 16776 12774 16788
rect 12989 16779 13047 16785
rect 12989 16776 13001 16779
rect 12768 16748 13001 16776
rect 12768 16736 12774 16748
rect 12989 16745 13001 16748
rect 13035 16745 13047 16779
rect 16758 16776 16764 16788
rect 16719 16748 16764 16776
rect 12989 16739 13047 16745
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 17402 16776 17408 16788
rect 17363 16748 17408 16776
rect 17402 16736 17408 16748
rect 17460 16736 17466 16788
rect 18230 16736 18236 16788
rect 18288 16776 18294 16788
rect 18325 16779 18383 16785
rect 18325 16776 18337 16779
rect 18288 16748 18337 16776
rect 18288 16736 18294 16748
rect 18325 16745 18337 16748
rect 18371 16745 18383 16779
rect 22646 16776 22652 16788
rect 22607 16748 22652 16776
rect 18325 16739 18383 16745
rect 22646 16736 22652 16748
rect 22704 16736 22710 16788
rect 22833 16779 22891 16785
rect 22833 16745 22845 16779
rect 22879 16776 22891 16779
rect 23014 16776 23020 16788
rect 22879 16748 23020 16776
rect 22879 16745 22891 16748
rect 22833 16739 22891 16745
rect 23014 16736 23020 16748
rect 23072 16736 23078 16788
rect 23934 16776 23940 16788
rect 23308 16748 23940 16776
rect 17310 16668 17316 16720
rect 17368 16708 17374 16720
rect 21910 16708 21916 16720
rect 17368 16680 21916 16708
rect 17368 16668 17374 16680
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 12713 16643 12771 16649
rect 12713 16609 12725 16643
rect 12759 16640 12771 16643
rect 14826 16640 14832 16652
rect 12759 16612 14832 16640
rect 12759 16609 12771 16612
rect 12713 16603 12771 16609
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 15010 16640 15016 16652
rect 14971 16612 15016 16640
rect 15010 16600 15016 16612
rect 15068 16600 15074 16652
rect 15286 16640 15292 16652
rect 15247 16612 15292 16640
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 17034 16600 17040 16652
rect 17092 16640 17098 16652
rect 18322 16640 18328 16652
rect 17092 16612 18328 16640
rect 17092 16600 17098 16612
rect 18322 16600 18328 16612
rect 18380 16600 18386 16652
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16572 12679 16575
rect 13354 16572 13360 16584
rect 12667 16544 13360 16572
rect 12667 16541 12679 16544
rect 12621 16535 12679 16541
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 17126 16532 17132 16584
rect 17184 16572 17190 16584
rect 17221 16575 17279 16581
rect 17221 16572 17233 16575
rect 17184 16544 17233 16572
rect 17184 16532 17190 16544
rect 17221 16541 17233 16544
rect 17267 16541 17279 16575
rect 17221 16535 17279 16541
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 18141 16575 18199 16581
rect 18141 16541 18153 16575
rect 18187 16572 18199 16575
rect 18432 16572 18460 16680
rect 21910 16668 21916 16680
rect 21968 16668 21974 16720
rect 19242 16600 19248 16652
rect 19300 16640 19306 16652
rect 19705 16643 19763 16649
rect 19705 16640 19717 16643
rect 19300 16612 19717 16640
rect 19300 16600 19306 16612
rect 19705 16609 19717 16612
rect 19751 16609 19763 16643
rect 23032 16640 23060 16736
rect 23198 16668 23204 16720
rect 23256 16708 23262 16720
rect 23308 16717 23336 16748
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 24026 16736 24032 16788
rect 24084 16776 24090 16788
rect 25041 16779 25099 16785
rect 25041 16776 25053 16779
rect 24084 16748 25053 16776
rect 24084 16736 24090 16748
rect 25041 16745 25053 16748
rect 25087 16745 25099 16779
rect 25041 16739 25099 16745
rect 25498 16736 25504 16788
rect 25556 16776 25562 16788
rect 25593 16779 25651 16785
rect 25593 16776 25605 16779
rect 25556 16748 25605 16776
rect 25556 16736 25562 16748
rect 25593 16745 25605 16748
rect 25639 16745 25651 16779
rect 27062 16776 27068 16788
rect 27023 16748 27068 16776
rect 25593 16739 25651 16745
rect 27062 16736 27068 16748
rect 27120 16736 27126 16788
rect 27614 16776 27620 16788
rect 27575 16748 27620 16776
rect 27614 16736 27620 16748
rect 27672 16736 27678 16788
rect 43898 16776 43904 16788
rect 43859 16748 43904 16776
rect 43898 16736 43904 16748
rect 43956 16736 43962 16788
rect 47210 16736 47216 16788
rect 47268 16776 47274 16788
rect 47854 16776 47860 16788
rect 47268 16748 47860 16776
rect 47268 16736 47274 16748
rect 47854 16736 47860 16748
rect 47912 16736 47918 16788
rect 23293 16711 23351 16717
rect 23293 16708 23305 16711
rect 23256 16680 23305 16708
rect 23256 16668 23262 16680
rect 23293 16677 23305 16680
rect 23339 16677 23351 16711
rect 23293 16671 23351 16677
rect 23382 16668 23388 16720
rect 23440 16708 23446 16720
rect 23440 16680 25544 16708
rect 23440 16668 23446 16680
rect 23032 16612 23704 16640
rect 19705 16603 19763 16609
rect 23676 16581 23704 16612
rect 23750 16600 23756 16652
rect 23808 16640 23814 16652
rect 23845 16643 23903 16649
rect 23845 16640 23857 16643
rect 23808 16612 23857 16640
rect 23808 16600 23814 16612
rect 23845 16609 23857 16612
rect 23891 16609 23903 16643
rect 23845 16603 23903 16609
rect 23934 16600 23940 16652
rect 23992 16640 23998 16652
rect 24489 16643 24547 16649
rect 24489 16640 24501 16643
rect 23992 16612 24501 16640
rect 23992 16600 23998 16612
rect 24489 16609 24501 16612
rect 24535 16609 24547 16643
rect 24489 16603 24547 16609
rect 24780 16612 25452 16640
rect 23569 16575 23627 16581
rect 23569 16572 23581 16575
rect 18187 16544 18460 16572
rect 21100 16544 23581 16572
rect 18187 16541 18199 16544
rect 18141 16535 18199 16541
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 2130 16504 2136 16516
rect 1627 16476 2136 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 16022 16464 16028 16516
rect 16080 16464 16086 16516
rect 18064 16504 18092 16535
rect 19889 16507 19947 16513
rect 18064 16476 18184 16504
rect 18156 16448 18184 16476
rect 19889 16473 19901 16507
rect 19935 16504 19947 16507
rect 19978 16504 19984 16516
rect 19935 16476 19984 16504
rect 19935 16473 19947 16476
rect 19889 16467 19947 16473
rect 19978 16464 19984 16476
rect 20036 16464 20042 16516
rect 18138 16436 18144 16448
rect 18051 16408 18144 16436
rect 18138 16396 18144 16408
rect 18196 16436 18202 16448
rect 21100 16436 21128 16544
rect 23569 16541 23581 16544
rect 23615 16541 23627 16575
rect 23569 16535 23627 16541
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16541 23719 16575
rect 24673 16575 24731 16581
rect 24673 16572 24685 16575
rect 23661 16535 23719 16541
rect 24412 16544 24685 16572
rect 21545 16507 21603 16513
rect 21545 16473 21557 16507
rect 21591 16504 21603 16507
rect 22278 16504 22284 16516
rect 21591 16476 22284 16504
rect 21591 16473 21603 16476
rect 21545 16467 21603 16473
rect 22278 16464 22284 16476
rect 22336 16464 22342 16516
rect 22465 16507 22523 16513
rect 22465 16473 22477 16507
rect 22511 16473 22523 16507
rect 24412 16504 24440 16544
rect 24673 16541 24685 16544
rect 24719 16572 24731 16575
rect 24780 16572 24808 16612
rect 24719 16544 24808 16572
rect 24719 16541 24731 16544
rect 24673 16535 24731 16541
rect 24854 16532 24860 16584
rect 24912 16532 24918 16584
rect 22465 16467 22523 16473
rect 23400 16476 24440 16504
rect 24765 16507 24823 16513
rect 18196 16408 21128 16436
rect 18196 16396 18202 16408
rect 22186 16396 22192 16448
rect 22244 16436 22250 16448
rect 22480 16436 22508 16467
rect 22244 16408 22508 16436
rect 22675 16439 22733 16445
rect 22244 16396 22250 16408
rect 22675 16405 22687 16439
rect 22721 16436 22733 16439
rect 23400 16436 23428 16476
rect 24765 16473 24777 16507
rect 24811 16504 24823 16507
rect 24872 16504 24900 16532
rect 24811 16476 24900 16504
rect 25424 16504 25452 16612
rect 25516 16581 25544 16680
rect 26881 16643 26939 16649
rect 26881 16609 26893 16643
rect 26927 16640 26939 16643
rect 26970 16640 26976 16652
rect 26927 16612 26976 16640
rect 26927 16609 26939 16612
rect 26881 16603 26939 16609
rect 26970 16600 26976 16612
rect 27028 16600 27034 16652
rect 45646 16640 45652 16652
rect 43824 16612 45652 16640
rect 25501 16575 25559 16581
rect 25501 16541 25513 16575
rect 25547 16541 25559 16575
rect 26786 16572 26792 16584
rect 26747 16544 26792 16572
rect 25501 16535 25559 16541
rect 26786 16532 26792 16544
rect 26844 16532 26850 16584
rect 27801 16575 27859 16581
rect 27801 16541 27813 16575
rect 27847 16572 27859 16575
rect 27890 16572 27896 16584
rect 27847 16544 27896 16572
rect 27847 16541 27859 16544
rect 27801 16535 27859 16541
rect 27890 16532 27896 16544
rect 27948 16532 27954 16584
rect 43824 16581 43852 16612
rect 45646 16600 45652 16612
rect 45704 16600 45710 16652
rect 46293 16643 46351 16649
rect 46293 16609 46305 16643
rect 46339 16640 46351 16643
rect 47762 16640 47768 16652
rect 46339 16612 47768 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47762 16600 47768 16612
rect 47820 16600 47826 16652
rect 43809 16575 43867 16581
rect 43809 16541 43821 16575
rect 43855 16541 43867 16575
rect 43809 16535 43867 16541
rect 26804 16504 26832 16532
rect 25424 16476 26832 16504
rect 46477 16507 46535 16513
rect 24811 16473 24823 16476
rect 24765 16467 24823 16473
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 47670 16504 47676 16516
rect 46523 16476 47676 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 22721 16408 23428 16436
rect 23477 16439 23535 16445
rect 22721 16405 22733 16408
rect 22675 16399 22733 16405
rect 23477 16405 23489 16439
rect 23523 16436 23535 16439
rect 24780 16436 24808 16467
rect 47670 16464 47676 16476
rect 47728 16464 47734 16516
rect 48130 16504 48136 16516
rect 48091 16476 48136 16504
rect 48130 16464 48136 16476
rect 48188 16464 48194 16516
rect 23523 16408 24808 16436
rect 24857 16439 24915 16445
rect 23523 16405 23535 16408
rect 23477 16399 23535 16405
rect 24857 16405 24869 16439
rect 24903 16436 24915 16439
rect 25406 16436 25412 16448
rect 24903 16408 25412 16436
rect 24903 16405 24915 16408
rect 24857 16399 24915 16405
rect 25406 16396 25412 16408
rect 25464 16396 25470 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 18141 16235 18199 16241
rect 18141 16201 18153 16235
rect 18187 16232 18199 16235
rect 18322 16232 18328 16244
rect 18187 16204 18328 16232
rect 18187 16201 18199 16204
rect 18141 16195 18199 16201
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 18785 16235 18843 16241
rect 18785 16201 18797 16235
rect 18831 16232 18843 16235
rect 18874 16232 18880 16244
rect 18831 16204 18880 16232
rect 18831 16201 18843 16204
rect 18785 16195 18843 16201
rect 18874 16192 18880 16204
rect 18932 16192 18938 16244
rect 19889 16235 19947 16241
rect 19889 16201 19901 16235
rect 19935 16232 19947 16235
rect 19978 16232 19984 16244
rect 19935 16204 19984 16232
rect 19935 16201 19947 16204
rect 19889 16195 19947 16201
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 39942 16232 39948 16244
rect 22066 16204 39948 16232
rect 17957 16167 18015 16173
rect 17957 16133 17969 16167
rect 18003 16164 18015 16167
rect 19242 16164 19248 16176
rect 18003 16136 19248 16164
rect 18003 16133 18015 16136
rect 17957 16127 18015 16133
rect 19242 16124 19248 16136
rect 19300 16124 19306 16176
rect 22066 16164 22094 16204
rect 39942 16192 39948 16204
rect 40000 16192 40006 16244
rect 19812 16136 22094 16164
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 2004 16068 2053 16096
rect 2004 16056 2010 16068
rect 2041 16065 2053 16068
rect 2087 16096 2099 16099
rect 15289 16099 15347 16105
rect 2087 16068 6914 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 6886 16028 6914 16068
rect 15289 16065 15301 16099
rect 15335 16065 15347 16099
rect 15289 16059 15347 16065
rect 6886 16000 12434 16028
rect 12406 15960 12434 16000
rect 14274 15988 14280 16040
rect 14332 16028 14338 16040
rect 15304 16028 15332 16059
rect 18230 16056 18236 16108
rect 18288 16096 18294 16108
rect 18288 16068 18333 16096
rect 18288 16056 18294 16068
rect 18414 16056 18420 16108
rect 18472 16096 18478 16108
rect 18693 16099 18751 16105
rect 18693 16096 18705 16099
rect 18472 16068 18705 16096
rect 18472 16056 18478 16068
rect 18693 16065 18705 16068
rect 18739 16096 18751 16099
rect 19150 16096 19156 16108
rect 18739 16068 19156 16096
rect 18739 16065 18751 16068
rect 18693 16059 18751 16065
rect 19150 16056 19156 16068
rect 19208 16056 19214 16108
rect 19812 16105 19840 16136
rect 22554 16124 22560 16176
rect 22612 16124 22618 16176
rect 24026 16124 24032 16176
rect 24084 16164 24090 16176
rect 24397 16167 24455 16173
rect 24397 16164 24409 16167
rect 24084 16136 24409 16164
rect 24084 16124 24090 16136
rect 24397 16133 24409 16136
rect 24443 16133 24455 16167
rect 24397 16127 24455 16133
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16096 21051 16099
rect 21634 16096 21640 16108
rect 21039 16068 21640 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 19812 16028 19840 16059
rect 21634 16056 21640 16068
rect 21692 16056 21698 16108
rect 25501 16099 25559 16105
rect 25501 16096 25513 16099
rect 24872 16068 25513 16096
rect 14332 16000 19840 16028
rect 21085 16031 21143 16037
rect 14332 15988 14338 16000
rect 21085 15997 21097 16031
rect 21131 16028 21143 16031
rect 21821 16031 21879 16037
rect 21821 16028 21833 16031
rect 21131 16000 21833 16028
rect 21131 15997 21143 16000
rect 21085 15991 21143 15997
rect 21821 15997 21833 16000
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 22094 15988 22100 16040
rect 22152 16028 22158 16040
rect 24872 16037 24900 16068
rect 25501 16065 25513 16068
rect 25547 16065 25559 16099
rect 44726 16096 44732 16108
rect 44687 16068 44732 16096
rect 25501 16059 25559 16065
rect 44726 16056 44732 16068
rect 44784 16056 44790 16108
rect 47762 16096 47768 16108
rect 47723 16068 47768 16096
rect 47762 16056 47768 16068
rect 47820 16056 47826 16108
rect 24857 16031 24915 16037
rect 22152 16000 22197 16028
rect 22152 15988 22158 16000
rect 24857 15997 24869 16031
rect 24903 15997 24915 16031
rect 24857 15991 24915 15997
rect 44913 16031 44971 16037
rect 44913 15997 44925 16031
rect 44959 16028 44971 16031
rect 45094 16028 45100 16040
rect 44959 16000 45100 16028
rect 44959 15997 44971 16000
rect 44913 15991 44971 15997
rect 45094 15988 45100 16000
rect 45152 15988 45158 16040
rect 46106 16028 46112 16040
rect 46067 16000 46112 16028
rect 46106 15988 46112 16000
rect 46164 15988 46170 16040
rect 17954 15960 17960 15972
rect 12406 15932 15516 15960
rect 17915 15932 17960 15960
rect 15378 15892 15384 15904
rect 15339 15864 15384 15892
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 15488 15892 15516 15932
rect 17954 15920 17960 15932
rect 18012 15920 18018 15972
rect 24765 15963 24823 15969
rect 24765 15929 24777 15963
rect 24811 15960 24823 15963
rect 24946 15960 24952 15972
rect 24811 15932 24952 15960
rect 24811 15929 24823 15932
rect 24765 15923 24823 15929
rect 24946 15920 24952 15932
rect 25004 15920 25010 15972
rect 25130 15920 25136 15972
rect 25188 15960 25194 15972
rect 25317 15963 25375 15969
rect 25317 15960 25329 15963
rect 25188 15932 25329 15960
rect 25188 15920 25194 15932
rect 25317 15929 25329 15932
rect 25363 15929 25375 15963
rect 25317 15923 25375 15929
rect 20806 15892 20812 15904
rect 15488 15864 20812 15892
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 22186 15852 22192 15904
rect 22244 15892 22250 15904
rect 23569 15895 23627 15901
rect 23569 15892 23581 15895
rect 22244 15864 23581 15892
rect 22244 15852 22250 15864
rect 23569 15861 23581 15864
rect 23615 15861 23627 15895
rect 23569 15855 23627 15861
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 20993 15691 21051 15697
rect 20993 15657 21005 15691
rect 21039 15688 21051 15691
rect 22094 15688 22100 15700
rect 21039 15660 22100 15688
rect 21039 15657 21051 15660
rect 20993 15651 21051 15657
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 22465 15691 22523 15697
rect 22465 15657 22477 15691
rect 22511 15688 22523 15691
rect 22554 15688 22560 15700
rect 22511 15660 22560 15688
rect 22511 15657 22523 15660
rect 22465 15651 22523 15657
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 45094 15688 45100 15700
rect 45055 15660 45100 15688
rect 45094 15648 45100 15660
rect 45152 15648 45158 15700
rect 47486 15648 47492 15700
rect 47544 15688 47550 15700
rect 47673 15691 47731 15697
rect 47673 15688 47685 15691
rect 47544 15660 47685 15688
rect 47544 15648 47550 15660
rect 47673 15657 47685 15660
rect 47719 15657 47731 15691
rect 47673 15651 47731 15657
rect 20530 15620 20536 15632
rect 15212 15592 20536 15620
rect 15212 15561 15240 15592
rect 20530 15580 20536 15592
rect 20588 15580 20594 15632
rect 22278 15580 22284 15632
rect 22336 15620 22342 15632
rect 45554 15620 45560 15632
rect 22336 15592 45560 15620
rect 22336 15580 22342 15592
rect 45554 15580 45560 15592
rect 45612 15580 45618 15632
rect 15197 15555 15255 15561
rect 15197 15521 15209 15555
rect 15243 15521 15255 15555
rect 15378 15552 15384 15564
rect 15339 15524 15384 15552
rect 15197 15515 15255 15521
rect 15378 15512 15384 15524
rect 15436 15512 15442 15564
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 14274 15484 14280 15496
rect 14235 15456 14280 15484
rect 2041 15447 2099 15453
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 18414 15484 18420 15496
rect 18375 15456 18420 15484
rect 18414 15444 18420 15456
rect 18472 15484 18478 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 18472 15456 19257 15484
rect 18472 15444 18478 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 20990 15484 20996 15496
rect 20951 15456 20996 15484
rect 19245 15447 19303 15453
rect 20990 15444 20996 15456
rect 21048 15444 21054 15496
rect 21177 15487 21235 15493
rect 21177 15453 21189 15487
rect 21223 15453 21235 15487
rect 21634 15484 21640 15496
rect 21595 15456 21640 15484
rect 21177 15447 21235 15453
rect 17034 15416 17040 15428
rect 16995 15388 17040 15416
rect 17034 15376 17040 15388
rect 17092 15376 17098 15428
rect 21192 15416 21220 15447
rect 21634 15444 21640 15456
rect 21692 15484 21698 15496
rect 22373 15487 22431 15493
rect 21692 15456 22094 15484
rect 21692 15444 21698 15456
rect 21910 15416 21916 15428
rect 21192 15388 21916 15416
rect 21910 15376 21916 15388
rect 21968 15376 21974 15428
rect 14366 15348 14372 15360
rect 14327 15320 14372 15348
rect 14366 15308 14372 15320
rect 14424 15308 14430 15360
rect 18506 15348 18512 15360
rect 18467 15320 18512 15348
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 19337 15351 19395 15357
rect 19337 15317 19349 15351
rect 19383 15348 19395 15351
rect 19978 15348 19984 15360
rect 19383 15320 19984 15348
rect 19383 15317 19395 15320
rect 19337 15311 19395 15317
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 21818 15348 21824 15360
rect 21779 15320 21824 15348
rect 21818 15308 21824 15320
rect 21876 15308 21882 15360
rect 22066 15348 22094 15456
rect 22373 15453 22385 15487
rect 22419 15484 22431 15487
rect 22830 15484 22836 15496
rect 22419 15456 22836 15484
rect 22419 15453 22431 15456
rect 22373 15447 22431 15453
rect 22830 15444 22836 15456
rect 22888 15444 22894 15496
rect 24857 15487 24915 15493
rect 24857 15453 24869 15487
rect 24903 15484 24915 15487
rect 25774 15484 25780 15496
rect 24903 15456 25780 15484
rect 24903 15453 24915 15456
rect 24857 15447 24915 15453
rect 25774 15444 25780 15456
rect 25832 15444 25838 15496
rect 45005 15487 45063 15493
rect 45005 15453 45017 15487
rect 45051 15484 45063 15487
rect 45646 15484 45652 15496
rect 45051 15456 45652 15484
rect 45051 15453 45063 15456
rect 45005 15447 45063 15453
rect 45646 15444 45652 15456
rect 45704 15444 45710 15496
rect 24394 15348 24400 15360
rect 22066 15320 24400 15348
rect 24394 15308 24400 15320
rect 24452 15348 24458 15360
rect 24949 15351 25007 15357
rect 24949 15348 24961 15351
rect 24452 15320 24961 15348
rect 24452 15308 24458 15320
rect 24949 15317 24961 15320
rect 24995 15317 25007 15351
rect 24949 15311 25007 15317
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 22189 15147 22247 15153
rect 22189 15144 22201 15147
rect 19444 15116 22201 15144
rect 13541 15079 13599 15085
rect 13541 15045 13553 15079
rect 13587 15076 13599 15079
rect 14366 15076 14372 15088
rect 13587 15048 14372 15076
rect 13587 15045 13599 15048
rect 13541 15039 13599 15045
rect 14366 15036 14372 15048
rect 14424 15036 14430 15088
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 13354 15008 13360 15020
rect 13315 14980 13360 15008
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 15654 15008 15660 15020
rect 15615 14980 15660 15008
rect 15654 14968 15660 14980
rect 15712 15008 15718 15020
rect 16574 15008 16580 15020
rect 15712 14980 16580 15008
rect 15712 14968 15718 14980
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 18230 14968 18236 15020
rect 18288 15008 18294 15020
rect 19444 15017 19472 15116
rect 22189 15113 22201 15116
rect 22235 15113 22247 15147
rect 22189 15107 22247 15113
rect 21542 15036 21548 15088
rect 21600 15076 21606 15088
rect 21821 15079 21879 15085
rect 21821 15076 21833 15079
rect 21600 15048 21833 15076
rect 21600 15036 21606 15048
rect 21821 15045 21833 15048
rect 21867 15045 21879 15079
rect 21821 15039 21879 15045
rect 21910 15036 21916 15088
rect 21968 15076 21974 15088
rect 22021 15079 22079 15085
rect 22021 15076 22033 15079
rect 21968 15048 22033 15076
rect 21968 15036 21974 15048
rect 22021 15045 22033 15048
rect 22067 15076 22079 15079
rect 23750 15076 23756 15088
rect 22067 15048 23756 15076
rect 22067 15045 22079 15048
rect 22021 15039 22079 15045
rect 23750 15036 23756 15048
rect 23808 15036 23814 15088
rect 19153 15011 19211 15017
rect 19153 15008 19165 15011
rect 18288 14980 19165 15008
rect 18288 14968 18294 14980
rect 19153 14977 19165 14980
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 14977 19487 15011
rect 19613 15011 19671 15017
rect 19613 15008 19625 15011
rect 19429 14971 19487 14977
rect 19536 14980 19625 15008
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 13817 14943 13875 14949
rect 13817 14909 13829 14943
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 16669 14943 16727 14949
rect 16669 14909 16681 14943
rect 16715 14909 16727 14943
rect 16850 14940 16856 14952
rect 16811 14912 16856 14940
rect 16669 14903 16727 14909
rect 12434 14832 12440 14884
rect 12492 14872 12498 14884
rect 13832 14872 13860 14903
rect 12492 14844 13860 14872
rect 16684 14872 16712 14903
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 18046 14940 18052 14952
rect 18007 14912 18052 14940
rect 18046 14900 18052 14912
rect 18104 14900 18110 14952
rect 19536 14872 19564 14980
rect 19613 14977 19625 14980
rect 19659 14977 19671 15011
rect 22830 15008 22836 15020
rect 22743 14980 22836 15008
rect 19613 14971 19671 14977
rect 22830 14968 22836 14980
rect 22888 15008 22894 15020
rect 23382 15008 23388 15020
rect 22888 14980 23388 15008
rect 22888 14968 22894 14980
rect 23382 14968 23388 14980
rect 23440 14968 23446 15020
rect 45646 14968 45652 15020
rect 45704 15008 45710 15020
rect 46569 15011 46627 15017
rect 46569 15008 46581 15011
rect 45704 14980 46581 15008
rect 45704 14968 45710 14980
rect 46569 14977 46581 14980
rect 46615 14977 46627 15011
rect 46569 14971 46627 14977
rect 20990 14872 20996 14884
rect 16684 14844 20996 14872
rect 12492 14832 12498 14844
rect 20990 14832 20996 14844
rect 21048 14832 21054 14884
rect 15470 14764 15476 14816
rect 15528 14804 15534 14816
rect 15749 14807 15807 14813
rect 15749 14804 15761 14807
rect 15528 14776 15761 14804
rect 15528 14764 15534 14776
rect 15749 14773 15761 14776
rect 15795 14773 15807 14807
rect 15749 14767 15807 14773
rect 18969 14807 19027 14813
rect 18969 14773 18981 14807
rect 19015 14804 19027 14807
rect 19518 14804 19524 14816
rect 19015 14776 19524 14804
rect 19015 14773 19027 14776
rect 18969 14767 19027 14773
rect 19518 14764 19524 14776
rect 19576 14764 19582 14816
rect 22002 14804 22008 14816
rect 21963 14776 22008 14804
rect 22002 14764 22008 14776
rect 22060 14764 22066 14816
rect 22830 14764 22836 14816
rect 22888 14804 22894 14816
rect 22925 14807 22983 14813
rect 22925 14804 22937 14807
rect 22888 14776 22937 14804
rect 22888 14764 22894 14776
rect 22925 14773 22937 14776
rect 22971 14773 22983 14807
rect 22925 14767 22983 14773
rect 46474 14764 46480 14816
rect 46532 14804 46538 14816
rect 46661 14807 46719 14813
rect 46661 14804 46673 14807
rect 46532 14776 46673 14804
rect 46532 14764 46538 14776
rect 46661 14773 46673 14776
rect 46707 14773 46719 14807
rect 46661 14767 46719 14773
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 20990 14600 20996 14612
rect 15304 14572 20576 14600
rect 20951 14572 20996 14600
rect 15304 14473 15332 14572
rect 18230 14532 18236 14544
rect 17880 14504 18236 14532
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14433 15347 14467
rect 15470 14464 15476 14476
rect 15431 14436 15476 14464
rect 15289 14427 15347 14433
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 17880 14473 17908 14504
rect 18230 14492 18236 14504
rect 18288 14492 18294 14544
rect 20548 14532 20576 14572
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 21542 14560 21548 14612
rect 21600 14600 21606 14612
rect 22281 14603 22339 14609
rect 22281 14600 22293 14603
rect 21600 14572 22293 14600
rect 21600 14560 21606 14572
rect 22281 14569 22293 14572
rect 22327 14569 22339 14603
rect 22281 14563 22339 14569
rect 22465 14603 22523 14609
rect 22465 14569 22477 14603
rect 22511 14600 22523 14603
rect 23106 14600 23112 14612
rect 22511 14572 23112 14600
rect 22511 14569 22523 14572
rect 22465 14563 22523 14569
rect 23106 14560 23112 14572
rect 23164 14560 23170 14612
rect 22186 14532 22192 14544
rect 20548 14504 22192 14532
rect 22186 14492 22192 14504
rect 22244 14492 22250 14544
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14433 17923 14467
rect 18138 14464 18144 14476
rect 18099 14436 18144 14464
rect 17865 14427 17923 14433
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 19518 14464 19524 14476
rect 19479 14436 19524 14464
rect 19518 14424 19524 14436
rect 19576 14424 19582 14476
rect 21910 14464 21916 14476
rect 21468 14436 21916 14464
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2682 14396 2688 14408
rect 2179 14368 2688 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 14274 14356 14280 14408
rect 14332 14396 14338 14408
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 14332 14368 14657 14396
rect 14332 14356 14338 14368
rect 14645 14365 14657 14368
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 17773 14399 17831 14405
rect 17773 14365 17785 14399
rect 17819 14396 17831 14399
rect 18230 14396 18236 14408
rect 17819 14368 18236 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 21468 14405 21496 14436
rect 21910 14424 21916 14436
rect 21968 14424 21974 14476
rect 23569 14467 23627 14473
rect 23569 14433 23581 14467
rect 23615 14464 23627 14467
rect 23750 14464 23756 14476
rect 23615 14436 23756 14464
rect 23615 14433 23627 14436
rect 23569 14427 23627 14433
rect 23750 14424 23756 14436
rect 23808 14424 23814 14476
rect 23845 14467 23903 14473
rect 23845 14433 23857 14467
rect 23891 14464 23903 14467
rect 24673 14467 24731 14473
rect 24673 14464 24685 14467
rect 23891 14436 24685 14464
rect 23891 14433 23903 14436
rect 23845 14427 23903 14433
rect 24673 14433 24685 14436
rect 24719 14433 24731 14467
rect 24673 14427 24731 14433
rect 19245 14399 19303 14405
rect 19245 14365 19257 14399
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 21453 14399 21511 14405
rect 21453 14365 21465 14399
rect 21499 14365 21511 14399
rect 21453 14359 21511 14365
rect 21637 14399 21695 14405
rect 21637 14365 21649 14399
rect 21683 14396 21695 14399
rect 22002 14396 22008 14408
rect 21683 14368 22008 14396
rect 21683 14365 21695 14368
rect 21637 14359 21695 14365
rect 17126 14328 17132 14340
rect 17087 14300 17132 14328
rect 17126 14288 17132 14300
rect 17184 14288 17190 14340
rect 19260 14328 19288 14359
rect 22002 14356 22008 14368
rect 22060 14396 22066 14408
rect 23477 14399 23535 14405
rect 23477 14396 23489 14399
rect 22060 14368 23489 14396
rect 22060 14356 22066 14368
rect 19426 14328 19432 14340
rect 19260 14300 19432 14328
rect 19426 14288 19432 14300
rect 19484 14288 19490 14340
rect 19978 14288 19984 14340
rect 20036 14288 20042 14340
rect 20990 14288 20996 14340
rect 21048 14328 21054 14340
rect 22296 14337 22324 14368
rect 23477 14365 23489 14368
rect 23523 14365 23535 14399
rect 23477 14359 23535 14365
rect 22097 14331 22155 14337
rect 22097 14328 22109 14331
rect 21048 14300 22109 14328
rect 21048 14288 21054 14300
rect 22097 14297 22109 14300
rect 22143 14297 22155 14331
rect 22296 14331 22355 14337
rect 22296 14300 22309 14331
rect 22097 14291 22155 14297
rect 22297 14297 22309 14300
rect 22343 14297 22355 14331
rect 22297 14291 22355 14297
rect 14737 14263 14795 14269
rect 14737 14229 14749 14263
rect 14783 14260 14795 14263
rect 15194 14260 15200 14272
rect 14783 14232 15200 14260
rect 14783 14229 14795 14232
rect 14737 14223 14795 14229
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 21634 14260 21640 14272
rect 21595 14232 21640 14260
rect 21634 14220 21640 14232
rect 21692 14220 21698 14272
rect 23492 14260 23520 14359
rect 24302 14356 24308 14408
rect 24360 14396 24366 14408
rect 24397 14399 24455 14405
rect 24397 14396 24409 14399
rect 24360 14368 24409 14396
rect 24360 14356 24366 14368
rect 24397 14365 24409 14368
rect 24443 14365 24455 14399
rect 24397 14359 24455 14365
rect 31205 14399 31263 14405
rect 31205 14365 31217 14399
rect 31251 14396 31263 14399
rect 32858 14396 32864 14408
rect 31251 14368 32864 14396
rect 31251 14365 31263 14368
rect 31205 14359 31263 14365
rect 32858 14356 32864 14368
rect 32916 14356 32922 14408
rect 45002 14396 45008 14408
rect 44963 14368 45008 14396
rect 45002 14356 45008 14368
rect 45060 14356 45066 14408
rect 25130 14288 25136 14340
rect 25188 14288 25194 14340
rect 45186 14328 45192 14340
rect 45147 14300 45192 14328
rect 45186 14288 45192 14300
rect 45244 14288 45250 14340
rect 46842 14328 46848 14340
rect 46803 14300 46848 14328
rect 46842 14288 46848 14300
rect 46900 14288 46906 14340
rect 26145 14263 26203 14269
rect 26145 14260 26157 14263
rect 23492 14232 26157 14260
rect 26145 14229 26157 14232
rect 26191 14260 26203 14263
rect 30374 14260 30380 14272
rect 26191 14232 30380 14260
rect 26191 14229 26203 14232
rect 26145 14223 26203 14229
rect 30374 14220 30380 14232
rect 30432 14220 30438 14272
rect 30558 14220 30564 14272
rect 30616 14260 30622 14272
rect 31297 14263 31355 14269
rect 31297 14260 31309 14263
rect 30616 14232 31309 14260
rect 30616 14220 30622 14232
rect 31297 14229 31309 14232
rect 31343 14229 31355 14263
rect 31297 14223 31355 14229
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 16850 14056 16856 14068
rect 15611 14028 16856 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 21542 14016 21548 14068
rect 21600 14056 21606 14068
rect 23569 14059 23627 14065
rect 23569 14056 23581 14059
rect 21600 14028 23581 14056
rect 21600 14016 21606 14028
rect 23569 14025 23581 14028
rect 23615 14025 23627 14059
rect 24302 14056 24308 14068
rect 24263 14028 24308 14056
rect 23569 14019 23627 14025
rect 24302 14016 24308 14028
rect 24360 14016 24366 14068
rect 25041 14059 25099 14065
rect 25041 14025 25053 14059
rect 25087 14056 25099 14059
rect 25130 14056 25136 14068
rect 25087 14028 25136 14056
rect 25087 14025 25099 14028
rect 25041 14019 25099 14025
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 45186 14056 45192 14068
rect 45147 14028 45192 14056
rect 45186 14016 45192 14028
rect 45244 14016 45250 14068
rect 17865 13991 17923 13997
rect 17865 13957 17877 13991
rect 17911 13988 17923 13991
rect 18138 13988 18144 14000
rect 17911 13960 18144 13988
rect 17911 13957 17923 13960
rect 17865 13951 17923 13957
rect 18138 13948 18144 13960
rect 18196 13948 18202 14000
rect 18506 13948 18512 14000
rect 18564 13948 18570 14000
rect 22830 13948 22836 14000
rect 22888 13948 22894 14000
rect 23382 13948 23388 14000
rect 23440 13988 23446 14000
rect 23440 13960 24992 13988
rect 23440 13948 23446 13960
rect 15473 13923 15531 13929
rect 15473 13889 15485 13923
rect 15519 13920 15531 13923
rect 15654 13920 15660 13932
rect 15519 13892 15660 13920
rect 15519 13889 15531 13892
rect 15473 13883 15531 13889
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 21818 13920 21824 13932
rect 21779 13892 21824 13920
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 24305 13923 24363 13929
rect 24305 13889 24317 13923
rect 24351 13920 24363 13923
rect 24394 13920 24400 13932
rect 24351 13892 24400 13920
rect 24351 13889 24363 13892
rect 24305 13883 24363 13889
rect 24394 13880 24400 13892
rect 24452 13880 24458 13932
rect 24964 13929 24992 13960
rect 24949 13923 25007 13929
rect 24949 13889 24961 13923
rect 24995 13889 25007 13923
rect 24949 13883 25007 13889
rect 44174 13880 44180 13932
rect 44232 13920 44238 13932
rect 45097 13923 45155 13929
rect 45097 13920 45109 13923
rect 44232 13892 45109 13920
rect 44232 13880 44238 13892
rect 45097 13889 45109 13892
rect 45143 13889 45155 13923
rect 45097 13883 45155 13889
rect 17589 13855 17647 13861
rect 17589 13821 17601 13855
rect 17635 13852 17647 13855
rect 17954 13852 17960 13864
rect 17635 13824 17960 13852
rect 17635 13821 17647 13824
rect 17589 13815 17647 13821
rect 17954 13812 17960 13824
rect 18012 13812 18018 13864
rect 18230 13812 18236 13864
rect 18288 13852 18294 13864
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 18288 13824 19625 13852
rect 18288 13812 18294 13824
rect 19613 13821 19625 13824
rect 19659 13852 19671 13855
rect 45002 13852 45008 13864
rect 19659 13824 45008 13852
rect 19659 13821 19671 13824
rect 19613 13815 19671 13821
rect 45002 13812 45008 13824
rect 45060 13812 45066 13864
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 15930 13784 15936 13796
rect 3476 13756 15936 13784
rect 3476 13744 3482 13756
rect 15930 13744 15936 13756
rect 15988 13744 15994 13796
rect 21818 13676 21824 13728
rect 21876 13716 21882 13728
rect 22078 13719 22136 13725
rect 22078 13716 22090 13719
rect 21876 13688 22090 13716
rect 21876 13676 21882 13688
rect 22078 13685 22090 13688
rect 22124 13685 22136 13719
rect 47762 13716 47768 13728
rect 47723 13688 47768 13716
rect 22078 13679 22136 13685
rect 47762 13676 47768 13688
rect 47820 13676 47826 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 17954 13512 17960 13524
rect 17915 13484 17960 13512
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 19426 13512 19432 13524
rect 19387 13484 19432 13512
rect 19426 13472 19432 13484
rect 19484 13472 19490 13524
rect 21818 13512 21824 13524
rect 21779 13484 21824 13512
rect 21818 13472 21824 13484
rect 21876 13472 21882 13524
rect 14642 13404 14648 13456
rect 14700 13444 14706 13456
rect 24394 13444 24400 13456
rect 14700 13416 15516 13444
rect 14700 13404 14706 13416
rect 15194 13376 15200 13388
rect 15155 13348 15200 13376
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 15488 13385 15516 13416
rect 19444 13416 24400 13444
rect 15473 13379 15531 13385
rect 15473 13345 15485 13379
rect 15519 13345 15531 13379
rect 15473 13339 15531 13345
rect 19444 13317 19472 13416
rect 24394 13404 24400 13416
rect 24452 13404 24458 13456
rect 47762 13444 47768 13456
rect 46308 13416 47768 13444
rect 21634 13376 21640 13388
rect 21595 13348 21640 13376
rect 21634 13336 21640 13348
rect 21692 13336 21698 13388
rect 30374 13376 30380 13388
rect 30335 13348 30380 13376
rect 30374 13336 30380 13348
rect 30432 13336 30438 13388
rect 30558 13376 30564 13388
rect 30519 13348 30564 13376
rect 30558 13336 30564 13348
rect 30616 13336 30622 13388
rect 46308 13385 46336 13416
rect 47762 13404 47768 13416
rect 47820 13404 47826 13456
rect 46293 13379 46351 13385
rect 46293 13345 46305 13379
rect 46339 13345 46351 13379
rect 46474 13376 46480 13388
rect 46435 13348 46480 13376
rect 46293 13339 46351 13345
rect 46474 13336 46480 13348
rect 46532 13336 46538 13388
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 18141 13311 18199 13317
rect 18141 13277 18153 13311
rect 18187 13308 18199 13311
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 18187 13280 19441 13308
rect 18187 13277 18199 13280
rect 18141 13271 18199 13277
rect 19429 13277 19441 13280
rect 19475 13277 19487 13311
rect 21542 13308 21548 13320
rect 21455 13280 21548 13308
rect 19429 13271 19487 13277
rect 15028 13240 15056 13271
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 21560 13240 21588 13268
rect 32214 13240 32220 13252
rect 15028 13212 21588 13240
rect 32175 13212 32220 13240
rect 32214 13200 32220 13212
rect 32272 13200 32278 13252
rect 48130 13240 48136 13252
rect 48091 13212 48136 13240
rect 48130 13200 48136 13212
rect 48188 13200 48194 13252
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 30466 12628 30472 12640
rect 1627 12600 30472 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 30466 12588 30472 12600
rect 30524 12588 30530 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 46290 12180 46296 12232
rect 46348 12220 46354 12232
rect 47673 12223 47731 12229
rect 47673 12220 47685 12223
rect 46348 12192 47685 12220
rect 46348 12180 46354 12192
rect 47673 12189 47685 12192
rect 47719 12189 47731 12223
rect 47673 12183 47731 12189
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 22462 11812 22468 11824
rect 22112 11784 22468 11812
rect 22112 11753 22140 11784
rect 22462 11772 22468 11784
rect 22520 11772 22526 11824
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 22278 11676 22284 11688
rect 22239 11648 22284 11676
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 23934 11676 23940 11688
rect 23895 11648 23940 11676
rect 23934 11636 23940 11648
rect 23992 11636 23998 11688
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 22278 11336 22284 11348
rect 22239 11308 22284 11336
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 46290 11200 46296 11212
rect 46251 11172 46296 11200
rect 46290 11160 46296 11172
rect 46348 11160 46354 11212
rect 22186 11132 22192 11144
rect 22147 11104 22192 11132
rect 22186 11092 22192 11104
rect 22244 11132 22250 11144
rect 38838 11132 38844 11144
rect 22244 11104 38844 11132
rect 22244 11092 22250 11104
rect 38838 11092 38844 11104
rect 38896 11092 38902 11144
rect 46014 11024 46020 11076
rect 46072 11064 46078 11076
rect 46477 11067 46535 11073
rect 46477 11064 46489 11067
rect 46072 11036 46489 11064
rect 46072 11024 46078 11036
rect 46477 11033 46489 11036
rect 46523 11033 46535 11067
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 46477 11027 46535 11033
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 12434 10996 12440 11008
rect 3200 10968 12440 10996
rect 3200 10956 3206 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 47118 10616 47124 10668
rect 47176 10656 47182 10668
rect 47486 10656 47492 10668
rect 47176 10628 47492 10656
rect 47176 10616 47182 10628
rect 47486 10616 47492 10628
rect 47544 10656 47550 10668
rect 47581 10659 47639 10665
rect 47581 10656 47593 10659
rect 47544 10628 47593 10656
rect 47544 10616 47550 10628
rect 47581 10625 47593 10628
rect 47627 10625 47639 10659
rect 47581 10619 47639 10625
rect 46290 10412 46296 10464
rect 46348 10452 46354 10464
rect 47029 10455 47087 10461
rect 47029 10452 47041 10455
rect 46348 10424 47041 10452
rect 46348 10412 46354 10424
rect 47029 10421 47041 10424
rect 47075 10421 47087 10455
rect 47670 10452 47676 10464
rect 47631 10424 47676 10452
rect 47029 10415 47087 10421
rect 47670 10412 47676 10424
rect 47728 10412 47734 10464
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 46477 10115 46535 10121
rect 46477 10081 46489 10115
rect 46523 10112 46535 10115
rect 47670 10112 47676 10124
rect 46523 10084 47676 10112
rect 46523 10081 46535 10084
rect 46477 10075 46535 10081
rect 47670 10072 47676 10084
rect 47728 10072 47734 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 47854 9568 47860 9580
rect 47815 9540 47860 9568
rect 47854 9528 47860 9540
rect 47912 9528 47918 9580
rect 48041 9435 48099 9441
rect 48041 9401 48053 9435
rect 48087 9432 48099 9435
rect 48222 9432 48228 9444
rect 48087 9404 48228 9432
rect 48087 9401 48099 9404
rect 48041 9395 48099 9401
rect 48222 9392 48228 9404
rect 48280 9392 48286 9444
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 47762 8888 47768 8900
rect 47723 8860 47768 8888
rect 47762 8848 47768 8860
rect 47820 8848 47826 8900
rect 28534 8780 28540 8832
rect 28592 8820 28598 8832
rect 47857 8823 47915 8829
rect 47857 8820 47869 8823
rect 28592 8792 47869 8820
rect 28592 8780 28598 8792
rect 47857 8789 47869 8792
rect 47903 8789 47915 8823
rect 47857 8783 47915 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 46934 8480 46940 8492
rect 46895 8452 46940 8480
rect 46934 8440 46940 8452
rect 46992 8440 46998 8492
rect 46753 8347 46811 8353
rect 46753 8313 46765 8347
rect 46799 8344 46811 8347
rect 47118 8344 47124 8356
rect 46799 8316 47124 8344
rect 46799 8313 46811 8316
rect 46753 8307 46811 8313
rect 47118 8304 47124 8316
rect 47176 8304 47182 8356
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 18046 8276 18052 8288
rect 3200 8248 18052 8276
rect 3200 8236 3206 8248
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 46477 7939 46535 7945
rect 46477 7905 46489 7939
rect 46523 7936 46535 7939
rect 46750 7936 46756 7948
rect 46523 7908 46756 7936
rect 46523 7905 46535 7908
rect 46477 7899 46535 7905
rect 46750 7896 46756 7908
rect 46808 7936 46814 7948
rect 47305 7939 47363 7945
rect 47305 7936 47317 7939
rect 46808 7908 47317 7936
rect 46808 7896 46814 7908
rect 47305 7905 47317 7908
rect 47351 7905 47363 7939
rect 47305 7899 47363 7905
rect 45462 7800 45468 7812
rect 45423 7772 45468 7800
rect 45462 7760 45468 7772
rect 45520 7760 45526 7812
rect 45554 7760 45560 7812
rect 45612 7800 45618 7812
rect 47026 7800 47032 7812
rect 45612 7772 45657 7800
rect 46987 7772 47032 7800
rect 45612 7760 45618 7772
rect 47026 7760 47032 7772
rect 47084 7760 47090 7812
rect 47118 7760 47124 7812
rect 47176 7800 47182 7812
rect 47176 7772 47221 7800
rect 47176 7760 47182 7772
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 46661 7531 46719 7537
rect 46661 7497 46673 7531
rect 46707 7528 46719 7531
rect 46934 7528 46940 7540
rect 46707 7500 46940 7528
rect 46707 7497 46719 7500
rect 46661 7491 46719 7497
rect 46934 7488 46940 7500
rect 46992 7488 46998 7540
rect 47026 7488 47032 7540
rect 47084 7528 47090 7540
rect 47949 7531 48007 7537
rect 47949 7528 47961 7531
rect 47084 7500 47961 7528
rect 47084 7488 47090 7500
rect 47949 7497 47961 7500
rect 47995 7497 48007 7531
rect 47949 7491 48007 7497
rect 45554 7352 45560 7404
rect 45612 7392 45618 7404
rect 46198 7392 46204 7404
rect 45612 7364 46204 7392
rect 45612 7352 45618 7364
rect 46198 7352 46204 7364
rect 46256 7352 46262 7404
rect 48130 7392 48136 7404
rect 48091 7364 48136 7392
rect 48130 7352 48136 7364
rect 48188 7352 48194 7404
rect 2038 7216 2044 7268
rect 2096 7256 2102 7268
rect 2096 7228 45554 7256
rect 2096 7216 2102 7228
rect 45526 7188 45554 7228
rect 45925 7191 45983 7197
rect 45925 7188 45937 7191
rect 45526 7160 45937 7188
rect 45925 7157 45937 7160
rect 45971 7188 45983 7191
rect 46293 7191 46351 7197
rect 46293 7188 46305 7191
rect 45971 7160 46305 7188
rect 45971 7157 45983 7160
rect 45925 7151 45983 7157
rect 46293 7157 46305 7160
rect 46339 7157 46351 7191
rect 46293 7151 46351 7157
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 17126 6848 17132 6860
rect 3476 6820 17132 6848
rect 3476 6808 3482 6820
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 47302 6848 47308 6860
rect 47263 6820 47308 6848
rect 47302 6808 47308 6820
rect 47360 6808 47366 6860
rect 47210 6740 47216 6792
rect 47268 6780 47274 6792
rect 47581 6783 47639 6789
rect 47581 6780 47593 6783
rect 47268 6752 47593 6780
rect 47268 6740 47274 6752
rect 47581 6749 47593 6752
rect 47627 6749 47639 6783
rect 47581 6743 47639 6749
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 46658 6400 46664 6452
rect 46716 6440 46722 6452
rect 48041 6443 48099 6449
rect 48041 6440 48053 6443
rect 46716 6412 48053 6440
rect 46716 6400 46722 6412
rect 48041 6409 48053 6412
rect 48087 6409 48099 6443
rect 48041 6403 48099 6409
rect 47946 6304 47952 6316
rect 47907 6276 47952 6304
rect 47946 6264 47952 6276
rect 48004 6264 48010 6316
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 41693 5763 41751 5769
rect 41693 5760 41705 5763
rect 4028 5732 41705 5760
rect 4028 5720 4034 5732
rect 41693 5729 41705 5732
rect 41739 5760 41751 5763
rect 42153 5763 42211 5769
rect 42153 5760 42165 5763
rect 41739 5732 42165 5760
rect 41739 5729 41751 5732
rect 41693 5723 41751 5729
rect 42153 5729 42165 5732
rect 42199 5729 42211 5763
rect 43162 5760 43168 5772
rect 43123 5732 43168 5760
rect 42153 5723 42211 5729
rect 43162 5720 43168 5732
rect 43220 5720 43226 5772
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 36725 5695 36783 5701
rect 36725 5692 36737 5695
rect 6696 5664 36737 5692
rect 6696 5652 6702 5664
rect 36725 5661 36737 5664
rect 36771 5661 36783 5695
rect 36725 5655 36783 5661
rect 36740 5624 36768 5655
rect 37185 5627 37243 5633
rect 37185 5624 37197 5627
rect 36740 5596 37197 5624
rect 37185 5593 37197 5596
rect 37231 5593 37243 5627
rect 37185 5587 37243 5593
rect 37274 5584 37280 5636
rect 37332 5624 37338 5636
rect 38197 5627 38255 5633
rect 37332 5596 37377 5624
rect 37332 5584 37338 5596
rect 38197 5593 38209 5627
rect 38243 5624 38255 5627
rect 38470 5624 38476 5636
rect 38243 5596 38476 5624
rect 38243 5593 38255 5596
rect 38197 5587 38255 5593
rect 38470 5584 38476 5596
rect 38528 5584 38534 5636
rect 42242 5584 42248 5636
rect 42300 5624 42306 5636
rect 42300 5596 42345 5624
rect 42300 5584 42306 5596
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 42242 5312 42248 5364
rect 42300 5352 42306 5364
rect 42429 5355 42487 5361
rect 42429 5352 42441 5355
rect 42300 5324 42441 5352
rect 42300 5312 42306 5324
rect 42429 5321 42441 5324
rect 42475 5321 42487 5355
rect 42429 5315 42487 5321
rect 45922 5312 45928 5364
rect 45980 5352 45986 5364
rect 48041 5355 48099 5361
rect 48041 5352 48053 5355
rect 45980 5324 48053 5352
rect 45980 5312 45986 5324
rect 48041 5321 48053 5324
rect 48087 5321 48099 5355
rect 48041 5315 48099 5321
rect 37734 5284 37740 5296
rect 37695 5256 37740 5284
rect 37734 5244 37740 5256
rect 37792 5244 37798 5296
rect 39761 5219 39819 5225
rect 39761 5185 39773 5219
rect 39807 5185 39819 5219
rect 40402 5216 40408 5228
rect 40363 5188 40408 5216
rect 39761 5179 39819 5185
rect 37642 5148 37648 5160
rect 37603 5120 37648 5148
rect 37642 5108 37648 5120
rect 37700 5108 37706 5160
rect 38470 5148 38476 5160
rect 38431 5120 38476 5148
rect 38470 5108 38476 5120
rect 38528 5108 38534 5160
rect 39776 5148 39804 5179
rect 40402 5176 40408 5188
rect 40460 5176 40466 5228
rect 42613 5219 42671 5225
rect 42613 5185 42625 5219
rect 42659 5216 42671 5219
rect 42886 5216 42892 5228
rect 42659 5188 42892 5216
rect 42659 5185 42671 5188
rect 42613 5179 42671 5185
rect 42886 5176 42892 5188
rect 42944 5176 42950 5228
rect 47857 5219 47915 5225
rect 47857 5185 47869 5219
rect 47903 5216 47915 5219
rect 48314 5216 48320 5228
rect 47903 5188 48320 5216
rect 47903 5185 47915 5188
rect 47857 5179 47915 5185
rect 48314 5176 48320 5188
rect 48372 5176 48378 5228
rect 41230 5148 41236 5160
rect 39776 5120 41236 5148
rect 41230 5108 41236 5120
rect 41288 5108 41294 5160
rect 39114 4972 39120 5024
rect 39172 5012 39178 5024
rect 39853 5015 39911 5021
rect 39853 5012 39865 5015
rect 39172 4984 39865 5012
rect 39172 4972 39178 4984
rect 39853 4981 39865 4984
rect 39899 4981 39911 5015
rect 39853 4975 39911 4981
rect 39942 4972 39948 5024
rect 40000 5012 40006 5024
rect 40497 5015 40555 5021
rect 40497 5012 40509 5015
rect 40000 4984 40509 5012
rect 40000 4972 40006 4984
rect 40497 4981 40509 4984
rect 40543 4981 40555 5015
rect 40497 4975 40555 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 37093 4811 37151 4817
rect 37093 4777 37105 4811
rect 37139 4808 37151 4811
rect 37274 4808 37280 4820
rect 37139 4780 37280 4808
rect 37139 4777 37151 4780
rect 37093 4771 37151 4777
rect 37274 4768 37280 4780
rect 37332 4768 37338 4820
rect 39209 4811 39267 4817
rect 39209 4777 39221 4811
rect 39255 4808 39267 4811
rect 40402 4808 40408 4820
rect 39255 4780 40408 4808
rect 39255 4777 39267 4780
rect 39209 4771 39267 4777
rect 40402 4768 40408 4780
rect 40460 4768 40466 4820
rect 41506 4700 41512 4752
rect 41564 4740 41570 4752
rect 45462 4740 45468 4752
rect 41564 4712 45468 4740
rect 41564 4700 41570 4712
rect 39942 4672 39948 4684
rect 39903 4644 39948 4672
rect 39942 4632 39948 4644
rect 40000 4632 40006 4684
rect 41782 4672 41788 4684
rect 41743 4644 41788 4672
rect 41782 4632 41788 4644
rect 41840 4632 41846 4684
rect 42628 4681 42656 4712
rect 45462 4700 45468 4712
rect 45520 4700 45526 4752
rect 46198 4700 46204 4752
rect 46256 4740 46262 4752
rect 46256 4712 47624 4740
rect 46256 4700 46262 4712
rect 42613 4675 42671 4681
rect 42613 4641 42625 4675
rect 42659 4641 42671 4675
rect 43162 4672 43168 4684
rect 43123 4644 43168 4672
rect 42613 4635 42671 4641
rect 43162 4632 43168 4644
rect 43220 4632 43226 4684
rect 47394 4672 47400 4684
rect 46676 4644 47400 4672
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 18325 4607 18383 4613
rect 18325 4604 18337 4607
rect 18104 4576 18337 4604
rect 18104 4564 18110 4576
rect 18325 4573 18337 4576
rect 18371 4573 18383 4607
rect 18325 4567 18383 4573
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4604 20683 4607
rect 21910 4604 21916 4616
rect 20671 4576 21916 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 21910 4564 21916 4576
rect 21968 4564 21974 4616
rect 37274 4604 37280 4616
rect 37235 4576 37280 4604
rect 37274 4564 37280 4576
rect 37332 4564 37338 4616
rect 39114 4604 39120 4616
rect 39075 4576 39120 4604
rect 39114 4564 39120 4576
rect 39172 4564 39178 4616
rect 46676 4613 46704 4644
rect 47394 4632 47400 4644
rect 47452 4632 47458 4684
rect 47596 4681 47624 4712
rect 47581 4675 47639 4681
rect 47581 4641 47593 4675
rect 47627 4641 47639 4675
rect 47581 4635 47639 4641
rect 46661 4607 46719 4613
rect 46661 4573 46673 4607
rect 46707 4573 46719 4607
rect 46661 4567 46719 4573
rect 46842 4564 46848 4616
rect 46900 4604 46906 4616
rect 47305 4607 47363 4613
rect 47305 4604 47317 4607
rect 46900 4576 47317 4604
rect 46900 4564 46906 4576
rect 47305 4573 47317 4576
rect 47351 4573 47363 4607
rect 47305 4567 47363 4573
rect 40126 4536 40132 4548
rect 40087 4508 40132 4536
rect 40126 4496 40132 4508
rect 40184 4496 40190 4548
rect 42705 4539 42763 4545
rect 42705 4505 42717 4539
rect 42751 4505 42763 4539
rect 42705 4499 42763 4505
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 14369 4471 14427 4477
rect 14369 4468 14381 4471
rect 14240 4440 14381 4468
rect 14240 4428 14246 4440
rect 14369 4437 14381 4440
rect 14415 4437 14427 4471
rect 14369 4431 14427 4437
rect 18230 4428 18236 4480
rect 18288 4468 18294 4480
rect 18417 4471 18475 4477
rect 18417 4468 18429 4471
rect 18288 4440 18429 4468
rect 18288 4428 18294 4440
rect 18417 4437 18429 4440
rect 18463 4437 18475 4471
rect 18417 4431 18475 4437
rect 20717 4471 20775 4477
rect 20717 4437 20729 4471
rect 20763 4468 20775 4471
rect 22370 4468 22376 4480
rect 20763 4440 22376 4468
rect 20763 4437 20775 4440
rect 20717 4431 20775 4437
rect 22370 4428 22376 4440
rect 22428 4428 22434 4480
rect 42518 4428 42524 4480
rect 42576 4468 42582 4480
rect 42720 4468 42748 4499
rect 42576 4440 42748 4468
rect 42576 4428 42582 4440
rect 46474 4428 46480 4480
rect 46532 4468 46538 4480
rect 46753 4471 46811 4477
rect 46753 4468 46765 4471
rect 46532 4440 46765 4468
rect 46532 4428 46538 4440
rect 46753 4437 46765 4440
rect 46799 4437 46811 4471
rect 46753 4431 46811 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 37274 4224 37280 4276
rect 37332 4264 37338 4276
rect 37737 4267 37795 4273
rect 37737 4264 37749 4267
rect 37332 4236 37749 4264
rect 37332 4224 37338 4236
rect 37737 4233 37749 4236
rect 37783 4233 37795 4267
rect 37737 4227 37795 4233
rect 27154 4196 27160 4208
rect 7116 4168 7328 4196
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2958 3952 2964 4004
rect 3016 3992 3022 4004
rect 7116 3992 7144 4168
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7300 4128 7328 4168
rect 15028 4168 15332 4196
rect 11790 4128 11796 4140
rect 7300 4100 11796 4128
rect 7193 4091 7251 4097
rect 7208 4060 7236 4091
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4128 11943 4131
rect 12802 4128 12808 4140
rect 11931 4100 12808 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 13265 4131 13323 4137
rect 13265 4128 13277 4131
rect 13044 4100 13277 4128
rect 13044 4088 13050 4100
rect 13265 4097 13277 4100
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4128 13415 4131
rect 13909 4131 13967 4137
rect 13909 4128 13921 4131
rect 13403 4100 13921 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 13909 4097 13921 4100
rect 13955 4097 13967 4131
rect 13909 4091 13967 4097
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4128 14059 4131
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14047 4100 14565 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 15028 4060 15056 4168
rect 15194 4128 15200 4140
rect 15155 4100 15200 4128
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 15304 4128 15332 4168
rect 21744 4168 22876 4196
rect 15304 4100 15516 4128
rect 7208 4032 15056 4060
rect 3016 3964 7144 3992
rect 3016 3952 3022 3964
rect 10410 3952 10416 4004
rect 10468 3992 10474 4004
rect 15010 3992 15016 4004
rect 10468 3964 15016 3992
rect 10468 3952 10474 3964
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 15488 3992 15516 4100
rect 15562 4088 15568 4140
rect 15620 4128 15626 4140
rect 15841 4131 15899 4137
rect 15841 4128 15853 4131
rect 15620 4100 15853 4128
rect 15620 4088 15626 4100
rect 15841 4097 15853 4100
rect 15887 4097 15899 4131
rect 16666 4128 16672 4140
rect 16627 4100 16672 4128
rect 15841 4091 15899 4097
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 16114 4020 16120 4072
rect 16172 4060 16178 4072
rect 17328 4060 17356 4091
rect 17586 4088 17592 4140
rect 17644 4128 17650 4140
rect 17957 4131 18015 4137
rect 17957 4128 17969 4131
rect 17644 4100 17969 4128
rect 17644 4088 17650 4100
rect 17957 4097 17969 4100
rect 18003 4097 18015 4131
rect 17957 4091 18015 4097
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 19242 4128 19248 4140
rect 19203 4100 19248 4128
rect 18601 4091 18659 4097
rect 16172 4032 17356 4060
rect 16172 4020 16178 4032
rect 17402 4020 17408 4072
rect 17460 4060 17466 4072
rect 18616 4060 18644 4091
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 20070 4128 20076 4140
rect 19935 4100 20076 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 20533 4131 20591 4137
rect 20533 4097 20545 4131
rect 20579 4128 20591 4131
rect 20806 4128 20812 4140
rect 20579 4100 20812 4128
rect 20579 4097 20591 4100
rect 20533 4091 20591 4097
rect 20806 4088 20812 4100
rect 20864 4088 20870 4140
rect 17460 4032 18644 4060
rect 17460 4020 17466 4032
rect 18782 4020 18788 4072
rect 18840 4060 18846 4072
rect 21744 4060 21772 4168
rect 21821 4131 21879 4137
rect 21821 4097 21833 4131
rect 21867 4097 21879 4131
rect 21821 4091 21879 4097
rect 21913 4131 21971 4137
rect 21913 4097 21925 4131
rect 21959 4128 21971 4131
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 21959 4100 22753 4128
rect 21959 4097 21971 4100
rect 21913 4091 21971 4097
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 22848 4128 22876 4168
rect 24044 4168 24256 4196
rect 27115 4168 27160 4196
rect 24044 4128 24072 4168
rect 22848 4100 24072 4128
rect 24121 4131 24179 4137
rect 22741 4091 22799 4097
rect 24121 4097 24133 4131
rect 24167 4097 24179 4131
rect 24228 4128 24256 4168
rect 27154 4156 27160 4168
rect 27212 4156 27218 4208
rect 37642 4196 37648 4208
rect 30944 4168 31340 4196
rect 24765 4131 24823 4137
rect 24765 4128 24777 4131
rect 24228 4100 24777 4128
rect 24121 4091 24179 4097
rect 24765 4097 24777 4100
rect 24811 4128 24823 4131
rect 25682 4128 25688 4140
rect 24811 4100 25688 4128
rect 24811 4097 24823 4100
rect 24765 4091 24823 4097
rect 18840 4032 21772 4060
rect 21836 4060 21864 4091
rect 22554 4060 22560 4072
rect 21836 4032 22560 4060
rect 18840 4020 18846 4032
rect 22554 4020 22560 4032
rect 22612 4020 22618 4072
rect 22186 3992 22192 4004
rect 15488 3964 22192 3992
rect 22186 3952 22192 3964
rect 22244 3952 22250 4004
rect 24136 3992 24164 4091
rect 25682 4088 25688 4100
rect 25740 4088 25746 4140
rect 30944 4128 30972 4168
rect 27908 4100 30972 4128
rect 24302 4020 24308 4072
rect 24360 4060 24366 4072
rect 27065 4063 27123 4069
rect 27065 4060 27077 4063
rect 24360 4032 27077 4060
rect 24360 4020 24366 4032
rect 27065 4029 27077 4032
rect 27111 4060 27123 4063
rect 27908 4060 27936 4100
rect 31018 4088 31024 4140
rect 31076 4128 31082 4140
rect 31312 4128 31340 4168
rect 37200 4168 37648 4196
rect 31570 4128 31576 4140
rect 31076 4100 31248 4128
rect 31312 4100 31576 4128
rect 31076 4088 31082 4100
rect 28074 4060 28080 4072
rect 27111 4032 27936 4060
rect 27987 4032 28080 4060
rect 27111 4029 27123 4032
rect 27065 4023 27123 4029
rect 28074 4020 28080 4032
rect 28132 4060 28138 4072
rect 31110 4060 31116 4072
rect 28132 4032 31116 4060
rect 28132 4020 28138 4032
rect 31110 4020 31116 4032
rect 31168 4020 31174 4072
rect 31220 4060 31248 4100
rect 31570 4088 31576 4100
rect 31628 4128 31634 4140
rect 37200 4128 37228 4168
rect 37642 4156 37648 4168
rect 37700 4196 37706 4208
rect 40310 4196 40316 4208
rect 37700 4168 39252 4196
rect 40271 4168 40316 4196
rect 37700 4156 37706 4168
rect 31628 4100 37228 4128
rect 37277 4131 37335 4137
rect 31628 4088 31634 4100
rect 37277 4097 37289 4131
rect 37323 4128 37335 4131
rect 37734 4128 37740 4140
rect 37323 4100 37740 4128
rect 37323 4097 37335 4100
rect 37277 4091 37335 4097
rect 37734 4088 37740 4100
rect 37792 4128 37798 4140
rect 38194 4128 38200 4140
rect 37792 4100 38200 4128
rect 37792 4088 37798 4100
rect 38194 4088 38200 4100
rect 38252 4088 38258 4140
rect 39224 4137 39252 4168
rect 40310 4156 40316 4168
rect 40368 4156 40374 4208
rect 46658 4196 46664 4208
rect 46619 4168 46664 4196
rect 46658 4156 46664 4168
rect 46716 4156 46722 4208
rect 47762 4196 47768 4208
rect 47723 4168 47768 4196
rect 47762 4156 47768 4168
rect 47820 4156 47826 4208
rect 39209 4131 39267 4137
rect 39209 4097 39221 4131
rect 39255 4128 39267 4131
rect 39298 4128 39304 4140
rect 39255 4100 39304 4128
rect 39255 4097 39267 4100
rect 39209 4091 39267 4097
rect 39298 4088 39304 4100
rect 39356 4088 39362 4140
rect 39393 4131 39451 4137
rect 39393 4097 39405 4131
rect 39439 4128 39451 4131
rect 40034 4128 40040 4140
rect 39439 4100 40040 4128
rect 39439 4097 39451 4100
rect 39393 4091 39451 4097
rect 40034 4088 40040 4100
rect 40092 4128 40098 4140
rect 40497 4131 40555 4137
rect 40497 4128 40509 4131
rect 40092 4100 40509 4128
rect 40092 4088 40098 4100
rect 40497 4097 40509 4100
rect 40543 4097 40555 4131
rect 40497 4091 40555 4097
rect 41141 4131 41199 4137
rect 41141 4097 41153 4131
rect 41187 4097 41199 4131
rect 41141 4091 41199 4097
rect 36538 4060 36544 4072
rect 31220 4032 36544 4060
rect 36538 4020 36544 4032
rect 36596 4020 36602 4072
rect 39853 4063 39911 4069
rect 39853 4029 39865 4063
rect 39899 4060 39911 4063
rect 41156 4060 41184 4091
rect 41230 4088 41236 4140
rect 41288 4128 41294 4140
rect 42429 4131 42487 4137
rect 41288 4100 41333 4128
rect 41288 4088 41294 4100
rect 42429 4097 42441 4131
rect 42475 4128 42487 4131
rect 42518 4128 42524 4140
rect 42475 4100 42524 4128
rect 42475 4097 42487 4100
rect 42429 4091 42487 4097
rect 42518 4088 42524 4100
rect 42576 4088 42582 4140
rect 42886 4060 42892 4072
rect 39899 4032 41184 4060
rect 42847 4032 42892 4060
rect 39899 4029 39911 4032
rect 39853 4023 39911 4029
rect 42886 4020 42892 4032
rect 42944 4020 42950 4072
rect 28810 3992 28816 4004
rect 24136 3964 28816 3992
rect 28810 3952 28816 3964
rect 28868 3952 28874 4004
rect 46845 3995 46903 4001
rect 46845 3992 46857 3995
rect 31726 3964 46857 3992
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1636 3896 2145 3924
rect 1636 3884 1642 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2866 3924 2872 3936
rect 2827 3896 2872 3924
rect 2133 3887 2191 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 7285 3927 7343 3933
rect 7285 3893 7297 3927
rect 7331 3924 7343 3927
rect 7374 3924 7380 3936
rect 7331 3896 7380 3924
rect 7331 3893 7343 3896
rect 7285 3887 7343 3893
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 11977 3927 12035 3933
rect 11977 3924 11989 3927
rect 11296 3896 11989 3924
rect 11296 3884 11302 3896
rect 11977 3893 11989 3896
rect 12023 3893 12035 3927
rect 11977 3887 12035 3893
rect 12066 3884 12072 3936
rect 12124 3924 12130 3936
rect 14550 3924 14556 3936
rect 12124 3896 14556 3924
rect 12124 3884 12130 3896
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14645 3927 14703 3933
rect 14645 3893 14657 3927
rect 14691 3924 14703 3927
rect 14734 3924 14740 3936
rect 14691 3896 14740 3924
rect 14691 3893 14703 3896
rect 14645 3887 14703 3893
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 15286 3924 15292 3936
rect 15247 3896 15292 3924
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 15378 3884 15384 3936
rect 15436 3924 15442 3936
rect 15933 3927 15991 3933
rect 15933 3924 15945 3927
rect 15436 3896 15945 3924
rect 15436 3884 15442 3896
rect 15933 3893 15945 3896
rect 15979 3893 15991 3927
rect 15933 3887 15991 3893
rect 16022 3884 16028 3936
rect 16080 3924 16086 3936
rect 16761 3927 16819 3933
rect 16761 3924 16773 3927
rect 16080 3896 16773 3924
rect 16080 3884 16086 3896
rect 16761 3893 16773 3896
rect 16807 3893 16819 3927
rect 16761 3887 16819 3893
rect 16850 3884 16856 3936
rect 16908 3924 16914 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 16908 3896 17417 3924
rect 16908 3884 16914 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 17405 3887 17463 3893
rect 17494 3884 17500 3936
rect 17552 3924 17558 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17552 3896 18061 3924
rect 17552 3884 17558 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18690 3924 18696 3936
rect 18651 3896 18696 3924
rect 18049 3887 18107 3893
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 19334 3924 19340 3936
rect 19295 3896 19340 3924
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 19981 3927 20039 3933
rect 19981 3893 19993 3927
rect 20027 3924 20039 3927
rect 20530 3924 20536 3936
rect 20027 3896 20536 3924
rect 20027 3893 20039 3896
rect 19981 3887 20039 3893
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 20625 3927 20683 3933
rect 20625 3893 20637 3927
rect 20671 3924 20683 3927
rect 21818 3924 21824 3936
rect 20671 3896 21824 3924
rect 20671 3893 20683 3896
rect 20625 3887 20683 3893
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 22830 3924 22836 3936
rect 22791 3896 22836 3924
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 23382 3884 23388 3936
rect 23440 3924 23446 3936
rect 24213 3927 24271 3933
rect 24213 3924 24225 3927
rect 23440 3896 24225 3924
rect 23440 3884 23446 3896
rect 24213 3893 24225 3896
rect 24259 3893 24271 3927
rect 24854 3924 24860 3936
rect 24815 3896 24860 3924
rect 24213 3887 24271 3893
rect 24854 3884 24860 3896
rect 24912 3884 24918 3936
rect 25590 3924 25596 3936
rect 25551 3896 25596 3924
rect 25590 3884 25596 3896
rect 25648 3884 25654 3936
rect 25958 3884 25964 3936
rect 26016 3924 26022 3936
rect 31726 3924 31754 3964
rect 46845 3961 46857 3964
rect 46891 3961 46903 3995
rect 46845 3955 46903 3961
rect 37366 3924 37372 3936
rect 26016 3896 31754 3924
rect 37327 3896 37372 3924
rect 26016 3884 26022 3896
rect 37366 3884 37372 3896
rect 37424 3884 37430 3936
rect 40218 3884 40224 3936
rect 40276 3924 40282 3936
rect 40681 3927 40739 3933
rect 40681 3924 40693 3927
rect 40276 3896 40693 3924
rect 40276 3884 40282 3896
rect 40681 3893 40693 3896
rect 40727 3893 40739 3927
rect 40681 3887 40739 3893
rect 41414 3884 41420 3936
rect 41472 3924 41478 3936
rect 42521 3927 42579 3933
rect 42521 3924 42533 3927
rect 41472 3896 42533 3924
rect 41472 3884 41478 3896
rect 42521 3893 42533 3896
rect 42567 3893 42579 3927
rect 42521 3887 42579 3893
rect 46109 3927 46167 3933
rect 46109 3893 46121 3927
rect 46155 3924 46167 3927
rect 46290 3924 46296 3936
rect 46155 3896 46296 3924
rect 46155 3893 46167 3896
rect 46109 3887 46167 3893
rect 46290 3884 46296 3896
rect 46348 3884 46354 3936
rect 47854 3924 47860 3936
rect 47815 3896 47860 3924
rect 47854 3884 47860 3896
rect 47912 3884 47918 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 44450 3720 44456 3732
rect 3936 3692 44456 3720
rect 3936 3680 3942 3692
rect 44450 3680 44456 3692
rect 44508 3680 44514 3732
rect 6546 3612 6552 3664
rect 6604 3652 6610 3664
rect 6604 3624 14136 3652
rect 6604 3612 6610 3624
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 1820 3556 3985 3584
rect 1820 3544 1826 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 3973 3547 4031 3553
rect 2682 3516 2688 3528
rect 2643 3488 2688 3516
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 6178 3516 6184 3528
rect 6139 3488 6184 3516
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 6656 3525 6684 3624
rect 11238 3584 11244 3596
rect 11199 3556 11244 3584
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11514 3584 11520 3596
rect 11475 3556 11520 3584
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 7190 3476 7196 3528
rect 7248 3516 7254 3528
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 7248 3488 7481 3516
rect 7248 3476 7254 3488
rect 7469 3485 7481 3488
rect 7515 3485 7527 3519
rect 10410 3516 10416 3528
rect 7469 3479 7527 3485
rect 9324 3488 9536 3516
rect 10371 3488 10416 3516
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 1857 3451 1915 3457
rect 1857 3448 1869 3451
rect 1360 3420 1869 3448
rect 1360 3408 1366 3420
rect 1857 3417 1869 3420
rect 1903 3417 1915 3451
rect 1857 3411 1915 3417
rect 2225 3451 2283 3457
rect 2225 3417 2237 3451
rect 2271 3448 2283 3451
rect 9324 3448 9352 3488
rect 2271 3420 9352 3448
rect 9401 3451 9459 3457
rect 2271 3417 2283 3420
rect 2225 3411 2283 3417
rect 9401 3417 9413 3451
rect 9447 3417 9459 3451
rect 9508 3448 9536 3488
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 11020 3488 11069 3516
rect 11020 3476 11026 3488
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13630 3516 13636 3528
rect 13587 3488 13636 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 14108 3525 14136 3624
rect 14274 3612 14280 3664
rect 14332 3652 14338 3664
rect 14829 3655 14887 3661
rect 14829 3652 14841 3655
rect 14332 3624 14841 3652
rect 14332 3612 14338 3624
rect 14829 3621 14841 3624
rect 14875 3621 14887 3655
rect 14829 3615 14887 3621
rect 15473 3655 15531 3661
rect 15473 3621 15485 3655
rect 15519 3652 15531 3655
rect 16666 3652 16672 3664
rect 15519 3624 16672 3652
rect 15519 3621 15531 3624
rect 15473 3615 15531 3621
rect 16666 3612 16672 3624
rect 16724 3612 16730 3664
rect 17402 3652 17408 3664
rect 17363 3624 17408 3652
rect 17402 3612 17408 3624
rect 17460 3612 17466 3664
rect 18046 3652 18052 3664
rect 18007 3624 18052 3652
rect 18046 3612 18052 3624
rect 18104 3612 18110 3664
rect 18138 3612 18144 3664
rect 18196 3652 18202 3664
rect 22646 3652 22652 3664
rect 18196 3624 22652 3652
rect 18196 3612 18202 3624
rect 22646 3612 22652 3624
rect 22704 3612 22710 3664
rect 22741 3655 22799 3661
rect 22741 3621 22753 3655
rect 22787 3652 22799 3655
rect 24302 3652 24308 3664
rect 22787 3624 24308 3652
rect 22787 3621 22799 3624
rect 22741 3615 22799 3621
rect 24302 3612 24308 3624
rect 24360 3612 24366 3664
rect 25590 3652 25596 3664
rect 24688 3624 25596 3652
rect 16114 3584 16120 3596
rect 16075 3556 16120 3584
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 22278 3584 22284 3596
rect 16592 3556 22284 3584
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3485 14151 3519
rect 14734 3516 14740 3528
rect 14695 3488 14740 3516
rect 14093 3479 14151 3485
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 15378 3516 15384 3528
rect 15068 3488 15240 3516
rect 15339 3488 15384 3516
rect 15068 3476 15074 3488
rect 9508 3420 11744 3448
rect 9401 3411 9459 3417
rect 2774 3380 2780 3392
rect 2735 3352 2780 3380
rect 2774 3340 2780 3352
rect 2832 3340 2838 3392
rect 6730 3380 6736 3392
rect 6691 3352 6736 3380
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 9416 3380 9444 3411
rect 8444 3352 9444 3380
rect 9677 3383 9735 3389
rect 8444 3340 8450 3352
rect 9677 3349 9689 3383
rect 9723 3380 9735 3383
rect 10318 3380 10324 3392
rect 9723 3352 10324 3380
rect 9723 3349 9735 3352
rect 9677 3343 9735 3349
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 10502 3380 10508 3392
rect 10463 3352 10508 3380
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 10870 3340 10876 3392
rect 10928 3380 10934 3392
rect 11514 3380 11520 3392
rect 10928 3352 11520 3380
rect 10928 3340 10934 3352
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 11716 3380 11744 3420
rect 12406 3420 14320 3448
rect 12406 3380 12434 3420
rect 11716 3352 12434 3380
rect 13814 3340 13820 3392
rect 13872 3380 13878 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 13872 3352 14197 3380
rect 13872 3340 13878 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14292 3380 14320 3420
rect 14366 3408 14372 3460
rect 14424 3448 14430 3460
rect 15102 3448 15108 3460
rect 14424 3420 15108 3448
rect 14424 3408 14430 3420
rect 15102 3408 15108 3420
rect 15160 3408 15166 3460
rect 15212 3448 15240 3488
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 16022 3516 16028 3528
rect 15983 3488 16028 3516
rect 16022 3476 16028 3488
rect 16080 3476 16086 3528
rect 16592 3448 16620 3556
rect 22278 3544 22284 3556
rect 22336 3544 22342 3596
rect 24688 3593 24716 3624
rect 25590 3612 25596 3624
rect 25648 3612 25654 3664
rect 25682 3612 25688 3664
rect 25740 3652 25746 3664
rect 36998 3652 37004 3664
rect 25740 3624 37004 3652
rect 25740 3612 25746 3624
rect 36998 3612 37004 3624
rect 37056 3612 37062 3664
rect 40037 3655 40095 3661
rect 40037 3621 40049 3655
rect 40083 3652 40095 3655
rect 40126 3652 40132 3664
rect 40083 3624 40132 3652
rect 40083 3621 40095 3624
rect 40037 3615 40095 3621
rect 40126 3612 40132 3624
rect 40184 3612 40190 3664
rect 47854 3652 47860 3664
rect 41386 3624 47860 3652
rect 24673 3587 24731 3593
rect 24673 3553 24685 3587
rect 24719 3553 24731 3587
rect 24854 3584 24860 3596
rect 24815 3556 24860 3584
rect 24673 3547 24731 3553
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 25130 3584 25136 3596
rect 25091 3556 25136 3584
rect 25130 3544 25136 3556
rect 25188 3544 25194 3596
rect 25222 3544 25228 3596
rect 25280 3584 25286 3596
rect 25280 3556 28994 3584
rect 25280 3544 25286 3556
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3516 16727 3519
rect 16850 3516 16856 3528
rect 16715 3488 16856 3516
rect 16715 3485 16727 3488
rect 16669 3479 16727 3485
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3516 17371 3519
rect 17494 3516 17500 3528
rect 17359 3488 17500 3516
rect 17359 3485 17371 3488
rect 17313 3479 17371 3485
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3516 18015 3519
rect 18690 3516 18696 3528
rect 18003 3488 18696 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 15212 3420 16620 3448
rect 16761 3451 16819 3457
rect 16761 3417 16773 3451
rect 16807 3448 16819 3451
rect 17586 3448 17592 3460
rect 16807 3420 17592 3448
rect 16807 3417 16819 3420
rect 16761 3411 16819 3417
rect 17586 3408 17592 3420
rect 17644 3408 17650 3460
rect 17770 3408 17776 3460
rect 17828 3448 17834 3460
rect 18782 3448 18788 3460
rect 17828 3420 18788 3448
rect 17828 3408 17834 3420
rect 18782 3408 18788 3420
rect 18840 3408 18846 3460
rect 19444 3448 19472 3479
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 20254 3516 20260 3528
rect 19576 3488 19621 3516
rect 20215 3488 20260 3516
rect 19576 3476 19582 3488
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 20530 3476 20536 3528
rect 20588 3516 20594 3528
rect 20717 3519 20775 3525
rect 20717 3516 20729 3519
rect 20588 3488 20729 3516
rect 20588 3476 20594 3488
rect 20717 3485 20729 3488
rect 20763 3485 20775 3519
rect 20717 3479 20775 3485
rect 20806 3476 20812 3528
rect 20864 3516 20870 3528
rect 22005 3519 22063 3525
rect 20864 3488 20909 3516
rect 20864 3476 20870 3488
rect 22005 3485 22017 3519
rect 22051 3516 22063 3519
rect 22094 3516 22100 3528
rect 22051 3488 22100 3516
rect 22051 3485 22063 3488
rect 22005 3479 22063 3485
rect 22094 3476 22100 3488
rect 22152 3476 22158 3528
rect 22830 3516 22836 3528
rect 22791 3488 22836 3516
rect 22830 3476 22836 3488
rect 22888 3476 22894 3528
rect 23198 3476 23204 3528
rect 23256 3516 23262 3528
rect 23661 3519 23719 3525
rect 23661 3516 23673 3519
rect 23256 3488 23673 3516
rect 23256 3476 23262 3488
rect 23661 3485 23673 3488
rect 23707 3485 23719 3519
rect 23661 3479 23719 3485
rect 27157 3519 27215 3525
rect 27157 3485 27169 3519
rect 27203 3516 27215 3519
rect 27430 3516 27436 3528
rect 27203 3488 27436 3516
rect 27203 3485 27215 3488
rect 27157 3479 27215 3485
rect 27430 3476 27436 3488
rect 27488 3476 27494 3528
rect 28966 3516 28994 3556
rect 30926 3544 30932 3596
rect 30984 3584 30990 3596
rect 32214 3584 32220 3596
rect 30984 3556 32220 3584
rect 30984 3544 30990 3556
rect 32214 3544 32220 3556
rect 32272 3544 32278 3596
rect 32950 3544 32956 3596
rect 33008 3584 33014 3596
rect 33873 3587 33931 3593
rect 33873 3584 33885 3587
rect 33008 3556 33885 3584
rect 33008 3544 33014 3556
rect 33873 3553 33885 3556
rect 33919 3553 33931 3587
rect 33873 3547 33931 3553
rect 36538 3544 36544 3596
rect 36596 3584 36602 3596
rect 41386 3584 41414 3624
rect 47854 3612 47860 3624
rect 47912 3612 47918 3664
rect 41782 3584 41788 3596
rect 36596 3556 41414 3584
rect 41743 3556 41788 3584
rect 36596 3544 36602 3556
rect 41782 3544 41788 3556
rect 41840 3544 41846 3596
rect 42426 3544 42432 3596
rect 42484 3584 42490 3596
rect 44177 3587 44235 3593
rect 44177 3584 44189 3587
rect 42484 3556 44189 3584
rect 42484 3544 42490 3556
rect 44177 3553 44189 3556
rect 44223 3553 44235 3587
rect 46290 3584 46296 3596
rect 46251 3556 46296 3584
rect 44177 3547 44235 3553
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 46474 3584 46480 3596
rect 46435 3556 46480 3584
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 31294 3516 31300 3528
rect 28966 3488 31300 3516
rect 31294 3476 31300 3488
rect 31352 3476 31358 3528
rect 33045 3519 33103 3525
rect 33045 3516 33057 3519
rect 31680 3488 33057 3516
rect 26602 3448 26608 3460
rect 19444 3420 26608 3448
rect 26602 3408 26608 3420
rect 26660 3408 26666 3460
rect 26786 3408 26792 3460
rect 26844 3448 26850 3460
rect 31680 3448 31708 3488
rect 33045 3485 33057 3488
rect 33091 3516 33103 3519
rect 38286 3516 38292 3528
rect 33091 3488 38292 3516
rect 33091 3485 33103 3488
rect 33045 3479 33103 3485
rect 38286 3476 38292 3488
rect 38344 3476 38350 3528
rect 40218 3516 40224 3528
rect 40179 3488 40224 3516
rect 40218 3476 40224 3488
rect 40276 3476 40282 3528
rect 41046 3516 41052 3528
rect 41007 3488 41052 3516
rect 41046 3476 41052 3488
rect 41104 3476 41110 3528
rect 43349 3519 43407 3525
rect 43349 3485 43361 3519
rect 43395 3485 43407 3519
rect 45186 3516 45192 3528
rect 45147 3488 45192 3516
rect 43349 3479 43407 3485
rect 26844 3420 31708 3448
rect 32968 3420 33272 3448
rect 26844 3408 26850 3420
rect 25222 3380 25228 3392
rect 14292 3352 25228 3380
rect 14185 3343 14243 3349
rect 25222 3340 25228 3352
rect 25280 3340 25286 3392
rect 26878 3340 26884 3392
rect 26936 3380 26942 3392
rect 26973 3383 27031 3389
rect 26973 3380 26985 3383
rect 26936 3352 26985 3380
rect 26936 3340 26942 3352
rect 26973 3349 26985 3352
rect 27019 3349 27031 3383
rect 26973 3343 27031 3349
rect 31478 3340 31484 3392
rect 31536 3380 31542 3392
rect 32968 3380 32996 3420
rect 33134 3380 33140 3392
rect 31536 3352 32996 3380
rect 33095 3352 33140 3380
rect 31536 3340 31542 3352
rect 33134 3340 33140 3352
rect 33192 3340 33198 3392
rect 33244 3380 33272 3420
rect 39850 3408 39856 3460
rect 39908 3448 39914 3460
rect 41233 3451 41291 3457
rect 41233 3448 41245 3451
rect 39908 3420 41245 3448
rect 39908 3408 39914 3420
rect 41233 3417 41245 3420
rect 41279 3417 41291 3451
rect 41233 3411 41291 3417
rect 41322 3408 41328 3460
rect 41380 3448 41386 3460
rect 43364 3448 43392 3479
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 45649 3519 45707 3525
rect 45649 3485 45661 3519
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 41380 3420 43392 3448
rect 45664 3448 45692 3479
rect 47486 3448 47492 3460
rect 45664 3420 47492 3448
rect 41380 3408 41386 3420
rect 47486 3408 47492 3420
rect 47544 3408 47550 3460
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 42334 3380 42340 3392
rect 33244 3352 42340 3380
rect 42334 3340 42340 3352
rect 42392 3340 42398 3392
rect 42610 3340 42616 3392
rect 42668 3380 42674 3392
rect 43441 3383 43499 3389
rect 43441 3380 43453 3383
rect 42668 3352 43453 3380
rect 42668 3340 42674 3352
rect 43441 3349 43453 3352
rect 43487 3349 43499 3383
rect 43441 3343 43499 3349
rect 45370 3340 45376 3392
rect 45428 3380 45434 3392
rect 45741 3383 45799 3389
rect 45741 3380 45753 3383
rect 45428 3352 45753 3380
rect 45428 3340 45434 3352
rect 45741 3349 45753 3352
rect 45787 3349 45799 3383
rect 45741 3343 45799 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 12986 3176 12992 3188
rect 2740 3148 11744 3176
rect 12947 3148 12992 3176
rect 2740 3136 2746 3148
rect 1949 3111 2007 3117
rect 1949 3077 1961 3111
rect 1995 3108 2007 3111
rect 2774 3108 2780 3120
rect 1995 3080 2780 3108
rect 1995 3077 2007 3080
rect 1949 3071 2007 3077
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 7374 3108 7380 3120
rect 7335 3080 7380 3108
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 11716 3108 11744 3148
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13648 3148 13952 3176
rect 13648 3108 13676 3148
rect 13814 3108 13820 3120
rect 11716 3080 13676 3108
rect 13775 3080 13820 3108
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 13924 3108 13952 3148
rect 14550 3136 14556 3188
rect 14608 3176 14614 3188
rect 17034 3176 17040 3188
rect 14608 3148 17040 3176
rect 14608 3136 14614 3148
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 18230 3136 18236 3188
rect 18288 3136 18294 3188
rect 18325 3179 18383 3185
rect 18325 3145 18337 3179
rect 18371 3176 18383 3179
rect 19242 3176 19248 3188
rect 18371 3148 19248 3176
rect 18371 3145 18383 3148
rect 18325 3139 18383 3145
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 20530 3176 20536 3188
rect 19352 3148 20536 3176
rect 17770 3108 17776 3120
rect 13924 3080 17776 3108
rect 17770 3068 17776 3080
rect 17828 3068 17834 3120
rect 18248 3055 18276 3136
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 7190 3040 7196 3052
rect 7151 3012 7196 3040
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 10962 3040 10968 3052
rect 10923 3012 10968 3040
rect 10962 3000 10968 3012
rect 11020 3000 11026 3052
rect 12069 3043 12127 3049
rect 12069 3009 12081 3043
rect 12115 3009 12127 3043
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 12069 3003 12127 3009
rect 12452 3012 12909 3040
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 716 2944 2237 2972
rect 716 2932 722 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 7742 2972 7748 2984
rect 7703 2944 7748 2972
rect 2225 2935 2283 2941
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 11974 2972 11980 2984
rect 11935 2944 11980 2972
rect 11974 2932 11980 2944
rect 12032 2932 12038 2984
rect 6454 2864 6460 2916
rect 6512 2904 6518 2916
rect 8202 2904 8208 2916
rect 6512 2876 8208 2904
rect 6512 2864 6518 2876
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 12084 2904 12112 3003
rect 12452 2981 12480 3012
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 13630 3040 13636 3052
rect 13591 3012 13636 3040
rect 12897 3003 12955 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 18241 3049 18299 3055
rect 15028 3012 15332 3040
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12802 2932 12808 2984
rect 12860 2972 12866 2984
rect 15028 2972 15056 3012
rect 12860 2944 15056 2972
rect 12860 2932 12866 2944
rect 15102 2932 15108 2984
rect 15160 2972 15166 2984
rect 15304 2972 15332 3012
rect 18241 3015 18253 3049
rect 18287 3015 18299 3049
rect 19352 3040 19380 3148
rect 20530 3136 20536 3148
rect 20588 3136 20594 3188
rect 21910 3176 21916 3188
rect 21871 3148 21916 3176
rect 21910 3136 21916 3148
rect 21968 3136 21974 3188
rect 22554 3176 22560 3188
rect 22515 3148 22560 3176
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 27062 3176 27068 3188
rect 23032 3148 27068 3176
rect 19518 3068 19524 3120
rect 19576 3108 19582 3120
rect 19576 3080 19621 3108
rect 19576 3068 19582 3080
rect 19702 3068 19708 3120
rect 19760 3108 19766 3120
rect 22922 3108 22928 3120
rect 19760 3080 22928 3108
rect 19760 3068 19766 3080
rect 22922 3068 22928 3080
rect 22980 3068 22986 3120
rect 18241 3009 18299 3015
rect 18340 3012 19380 3040
rect 15160 2944 15205 2972
rect 15304 2956 18276 2972
rect 18340 2956 18368 3012
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 21177 3043 21235 3049
rect 21177 3040 21189 3043
rect 20772 3012 21189 3040
rect 20772 3000 20778 3012
rect 21177 3009 21189 3012
rect 21223 3009 21235 3043
rect 21818 3040 21824 3052
rect 21779 3012 21824 3040
rect 21177 3003 21235 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 22370 3000 22376 3052
rect 22428 3040 22434 3052
rect 22473 3043 22531 3049
rect 22473 3040 22485 3043
rect 22428 3012 22485 3040
rect 22428 3000 22434 3012
rect 22473 3009 22485 3012
rect 22519 3009 22531 3043
rect 23032 3040 23060 3148
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 39850 3176 39856 3188
rect 30760 3148 36584 3176
rect 39811 3148 39856 3176
rect 23382 3108 23388 3120
rect 23343 3080 23388 3108
rect 23382 3068 23388 3080
rect 23440 3068 23446 3120
rect 23474 3068 23480 3120
rect 23532 3108 23538 3120
rect 26050 3108 26056 3120
rect 23532 3080 26056 3108
rect 23532 3068 23538 3080
rect 26050 3068 26056 3080
rect 26108 3068 26114 3120
rect 26878 3068 26884 3120
rect 26936 3108 26942 3120
rect 27157 3111 27215 3117
rect 27157 3108 27169 3111
rect 26936 3080 27169 3108
rect 26936 3068 26942 3080
rect 27157 3077 27169 3080
rect 27203 3077 27215 3111
rect 28074 3108 28080 3120
rect 28035 3080 28080 3108
rect 27157 3071 27215 3077
rect 28074 3068 28080 3080
rect 28132 3068 28138 3120
rect 28626 3068 28632 3120
rect 28684 3108 28690 3120
rect 30760 3108 30788 3148
rect 33134 3108 33140 3120
rect 28684 3080 30788 3108
rect 33095 3080 33140 3108
rect 28684 3068 28690 3080
rect 33134 3068 33140 3080
rect 33192 3068 33198 3120
rect 36556 3108 36584 3148
rect 39850 3136 39856 3148
rect 39908 3136 39914 3188
rect 41046 3136 41052 3188
rect 41104 3176 41110 3188
rect 41141 3179 41199 3185
rect 41141 3176 41153 3179
rect 41104 3148 41153 3176
rect 41104 3136 41110 3148
rect 41141 3145 41153 3148
rect 41187 3145 41199 3179
rect 41141 3139 41199 3145
rect 42610 3108 42616 3120
rect 36556 3080 41920 3108
rect 42571 3080 42616 3108
rect 23198 3040 23204 3052
rect 22473 3003 22531 3009
rect 22572 3012 23060 3040
rect 23159 3012 23204 3040
rect 15304 2944 18368 2956
rect 15160 2932 15166 2944
rect 18248 2928 18368 2944
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 19383 2944 19564 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 18138 2904 18144 2916
rect 12084 2876 18144 2904
rect 18138 2864 18144 2876
rect 18196 2864 18202 2916
rect 19536 2904 19564 2944
rect 20162 2932 20168 2984
rect 20220 2972 20226 2984
rect 22572 2972 22600 3012
rect 23198 3000 23204 3012
rect 23256 3000 23262 3052
rect 26237 3043 26295 3049
rect 26237 3009 26249 3043
rect 26283 3040 26295 3043
rect 26418 3040 26424 3052
rect 26283 3012 26424 3040
rect 26283 3009 26295 3012
rect 26237 3003 26295 3009
rect 26418 3000 26424 3012
rect 26476 3000 26482 3052
rect 32950 3040 32956 3052
rect 32911 3012 32956 3040
rect 32950 3000 32956 3012
rect 33008 3000 33014 3052
rect 39393 3043 39451 3049
rect 39393 3009 39405 3043
rect 39439 3040 39451 3043
rect 39942 3040 39948 3052
rect 39439 3012 39948 3040
rect 39439 3009 39451 3012
rect 39393 3003 39451 3009
rect 39942 3000 39948 3012
rect 40000 3000 40006 3052
rect 40037 3043 40095 3049
rect 40037 3009 40049 3043
rect 40083 3040 40095 3043
rect 40586 3040 40592 3052
rect 40083 3012 40592 3040
rect 40083 3009 40095 3012
rect 40037 3003 40095 3009
rect 40586 3000 40592 3012
rect 40644 3000 40650 3052
rect 41230 3000 41236 3052
rect 41288 3040 41294 3052
rect 41785 3043 41843 3049
rect 41785 3040 41797 3043
rect 41288 3012 41797 3040
rect 41288 3000 41294 3012
rect 41785 3009 41797 3012
rect 41831 3009 41843 3043
rect 41785 3003 41843 3009
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 20220 2944 22600 2972
rect 22756 2944 23673 2972
rect 20220 2932 20226 2944
rect 20254 2904 20260 2916
rect 19536 2876 20260 2904
rect 20254 2864 20260 2876
rect 20312 2864 20318 2916
rect 22002 2904 22008 2916
rect 20364 2876 22008 2904
rect 9766 2836 9772 2848
rect 9727 2808 9772 2836
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 10318 2796 10324 2848
rect 10376 2836 10382 2848
rect 20364 2836 20392 2876
rect 22002 2864 22008 2876
rect 22060 2864 22066 2916
rect 22554 2864 22560 2916
rect 22612 2904 22618 2916
rect 22756 2904 22784 2944
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 27065 2975 27123 2981
rect 27065 2972 27077 2975
rect 23661 2935 23719 2941
rect 25148 2944 27077 2972
rect 22612 2876 22784 2904
rect 22612 2864 22618 2876
rect 23474 2864 23480 2916
rect 23532 2904 23538 2916
rect 25148 2904 25176 2944
rect 27065 2941 27077 2944
rect 27111 2941 27123 2975
rect 27065 2935 27123 2941
rect 27154 2932 27160 2984
rect 27212 2972 27218 2984
rect 32214 2972 32220 2984
rect 27212 2944 32220 2972
rect 27212 2932 27218 2944
rect 32214 2932 32220 2944
rect 32272 2932 32278 2984
rect 33502 2972 33508 2984
rect 33463 2944 33508 2972
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 39298 2932 39304 2984
rect 39356 2972 39362 2984
rect 40497 2975 40555 2981
rect 40497 2972 40509 2975
rect 39356 2944 40509 2972
rect 39356 2932 39362 2944
rect 40497 2941 40509 2944
rect 40543 2941 40555 2975
rect 40678 2972 40684 2984
rect 40639 2944 40684 2972
rect 40497 2935 40555 2941
rect 38378 2904 38384 2916
rect 23532 2876 25176 2904
rect 26206 2876 38384 2904
rect 23532 2864 23538 2876
rect 10376 2808 20392 2836
rect 10376 2796 10382 2808
rect 20530 2796 20536 2848
rect 20588 2836 20594 2848
rect 26206 2836 26234 2876
rect 38378 2864 38384 2876
rect 38436 2864 38442 2916
rect 39209 2907 39267 2913
rect 39209 2873 39221 2907
rect 39255 2904 39267 2907
rect 40034 2904 40040 2916
rect 39255 2876 40040 2904
rect 39255 2873 39267 2876
rect 39209 2867 39267 2873
rect 40034 2864 40040 2876
rect 40092 2864 40098 2916
rect 40512 2904 40540 2935
rect 40678 2932 40684 2944
rect 40736 2972 40742 2984
rect 40736 2944 41644 2972
rect 40736 2932 40742 2944
rect 41506 2904 41512 2916
rect 40512 2876 41512 2904
rect 41506 2864 41512 2876
rect 41564 2864 41570 2916
rect 41616 2913 41644 2944
rect 41601 2907 41659 2913
rect 41601 2873 41613 2907
rect 41647 2873 41659 2907
rect 41892 2904 41920 3080
rect 42610 3068 42616 3080
rect 42668 3068 42674 3120
rect 45370 3108 45376 3120
rect 45331 3080 45376 3108
rect 45370 3068 45376 3080
rect 45428 3068 45434 3120
rect 42426 3040 42432 3052
rect 42387 3012 42432 3040
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 46750 3000 46756 3052
rect 46808 3040 46814 3052
rect 47765 3043 47823 3049
rect 47765 3040 47777 3043
rect 46808 3012 47777 3040
rect 46808 3000 46814 3012
rect 47765 3009 47777 3012
rect 47811 3009 47823 3043
rect 47765 3003 47823 3009
rect 43162 2972 43168 2984
rect 43123 2944 43168 2972
rect 43162 2932 43168 2944
rect 43220 2932 43226 2984
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 47949 2907 48007 2913
rect 47949 2904 47961 2907
rect 41892 2876 47961 2904
rect 41601 2867 41659 2873
rect 47949 2873 47961 2876
rect 47995 2873 48007 2907
rect 47949 2867 48007 2873
rect 20588 2808 26234 2836
rect 26329 2839 26387 2845
rect 20588 2796 20594 2808
rect 26329 2805 26341 2839
rect 26375 2836 26387 2839
rect 30650 2836 30656 2848
rect 26375 2808 30656 2836
rect 26375 2805 26387 2808
rect 26329 2799 26387 2805
rect 30650 2796 30656 2808
rect 30708 2796 30714 2848
rect 38286 2796 38292 2848
rect 38344 2836 38350 2848
rect 41322 2836 41328 2848
rect 38344 2808 41328 2836
rect 38344 2796 38350 2808
rect 41322 2796 41328 2808
rect 41380 2796 41386 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 3973 2635 4031 2641
rect 3973 2601 3985 2635
rect 4019 2632 4031 2635
rect 14277 2635 14335 2641
rect 4019 2604 9996 2632
rect 4019 2601 4031 2604
rect 3973 2595 4031 2601
rect 2866 2564 2872 2576
rect 1412 2536 2872 2564
rect 1412 2505 1440 2536
rect 2866 2524 2872 2536
rect 2924 2524 2930 2576
rect 9030 2524 9036 2576
rect 9088 2564 9094 2576
rect 9088 2536 9904 2564
rect 9088 2524 9094 2536
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1397 2459 1455 2465
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 2832 2468 2877 2496
rect 2832 2456 2838 2468
rect 6178 2456 6184 2508
rect 6236 2496 6242 2508
rect 6549 2499 6607 2505
rect 6549 2496 6561 2499
rect 6236 2468 6561 2496
rect 6236 2456 6242 2468
rect 6549 2465 6561 2468
rect 6595 2465 6607 2499
rect 6730 2496 6736 2508
rect 6691 2468 6736 2496
rect 6549 2459 6607 2465
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 7098 2496 7104 2508
rect 7059 2468 7104 2496
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 9125 2499 9183 2505
rect 9125 2465 9137 2499
rect 9171 2496 9183 2499
rect 9766 2496 9772 2508
rect 9171 2468 9772 2496
rect 9171 2465 9183 2468
rect 9125 2459 9183 2465
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 9876 2505 9904 2536
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2465 9919 2499
rect 9968 2496 9996 2604
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 15194 2632 15200 2644
rect 14323 2604 15200 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 19337 2635 19395 2641
rect 16546 2604 19288 2632
rect 10042 2524 10048 2576
rect 10100 2564 10106 2576
rect 16546 2564 16574 2604
rect 10100 2536 16574 2564
rect 10100 2524 10106 2536
rect 16758 2496 16764 2508
rect 9968 2468 16764 2496
rect 9861 2459 9919 2465
rect 16758 2456 16764 2468
rect 16816 2456 16822 2508
rect 19260 2496 19288 2604
rect 19337 2601 19349 2635
rect 19383 2632 19395 2635
rect 20070 2632 20076 2644
rect 19383 2604 20076 2632
rect 19383 2601 19395 2604
rect 19337 2595 19395 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 20901 2635 20959 2641
rect 20901 2632 20913 2635
rect 20496 2604 20913 2632
rect 20496 2592 20502 2604
rect 20901 2601 20913 2604
rect 20947 2601 20959 2635
rect 20901 2595 20959 2601
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 22373 2635 22431 2641
rect 22373 2632 22385 2635
rect 22152 2604 22385 2632
rect 22152 2592 22158 2604
rect 22373 2601 22385 2604
rect 22419 2601 22431 2635
rect 22373 2595 22431 2601
rect 23385 2635 23443 2641
rect 23385 2601 23397 2635
rect 23431 2632 23443 2635
rect 23474 2632 23480 2644
rect 23431 2604 23480 2632
rect 23431 2601 23443 2604
rect 23385 2595 23443 2601
rect 23474 2592 23480 2604
rect 23532 2592 23538 2644
rect 27249 2635 27307 2641
rect 27249 2601 27261 2635
rect 27295 2601 27307 2635
rect 27430 2632 27436 2644
rect 27391 2604 27436 2632
rect 27249 2595 27307 2601
rect 25038 2564 25044 2576
rect 24999 2536 25044 2564
rect 25038 2524 25044 2536
rect 25096 2524 25102 2576
rect 27264 2564 27292 2595
rect 27430 2592 27436 2604
rect 27488 2592 27494 2644
rect 35342 2592 35348 2644
rect 35400 2632 35406 2644
rect 35400 2604 35664 2632
rect 35400 2592 35406 2604
rect 35529 2567 35587 2573
rect 35529 2564 35541 2567
rect 27264 2536 35541 2564
rect 35529 2533 35541 2536
rect 35575 2533 35587 2567
rect 35636 2564 35664 2604
rect 35894 2592 35900 2644
rect 35952 2632 35958 2644
rect 39209 2635 39267 2641
rect 39209 2632 39221 2635
rect 35952 2604 39221 2632
rect 35952 2592 35958 2604
rect 39209 2601 39221 2604
rect 39255 2601 39267 2635
rect 40310 2632 40316 2644
rect 40271 2604 40316 2632
rect 39209 2595 39267 2601
rect 40310 2592 40316 2604
rect 40368 2592 40374 2644
rect 40586 2632 40592 2644
rect 40547 2604 40592 2632
rect 40586 2592 40592 2604
rect 40644 2592 40650 2644
rect 48038 2632 48044 2644
rect 47999 2604 48044 2632
rect 48038 2592 48044 2604
rect 48096 2592 48102 2644
rect 36449 2567 36507 2573
rect 36449 2564 36461 2567
rect 35636 2536 36461 2564
rect 35529 2527 35587 2533
rect 36449 2533 36461 2536
rect 36495 2533 36507 2567
rect 36449 2527 36507 2533
rect 38289 2567 38347 2573
rect 38289 2533 38301 2567
rect 38335 2533 38347 2567
rect 38289 2527 38347 2533
rect 41325 2567 41383 2573
rect 41325 2533 41337 2567
rect 41371 2564 41383 2567
rect 41874 2564 41880 2576
rect 41371 2536 41880 2564
rect 41371 2533 41383 2536
rect 41325 2527 41383 2533
rect 23934 2496 23940 2508
rect 19260 2468 23940 2496
rect 23934 2456 23940 2468
rect 23992 2456 23998 2508
rect 26421 2499 26479 2505
rect 26421 2465 26433 2499
rect 26467 2496 26479 2499
rect 27982 2496 27988 2508
rect 26467 2468 27988 2496
rect 26467 2465 26479 2468
rect 26421 2459 26479 2465
rect 27982 2456 27988 2468
rect 28040 2456 28046 2508
rect 32674 2456 32680 2508
rect 32732 2496 32738 2508
rect 35894 2496 35900 2508
rect 32732 2468 35900 2496
rect 32732 2456 32738 2468
rect 35894 2456 35900 2468
rect 35952 2456 35958 2508
rect 38304 2496 38332 2527
rect 41874 2524 41880 2536
rect 41932 2524 41938 2576
rect 36004 2468 38332 2496
rect 40313 2499 40371 2505
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3160 2400 3801 2428
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 3160 2360 3188 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5224 2400 5457 2428
rect 5224 2388 5230 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 14182 2428 14188 2440
rect 14143 2400 14188 2428
rect 5445 2391 5503 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2428 14887 2431
rect 15286 2428 15292 2440
rect 14875 2400 15292 2428
rect 14875 2397 14887 2400
rect 14829 2391 14887 2397
rect 15286 2388 15292 2400
rect 15344 2388 15350 2440
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16172 2400 16681 2428
rect 16172 2388 16178 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2428 19303 2431
rect 19334 2428 19340 2440
rect 19291 2400 19340 2428
rect 19291 2397 19303 2400
rect 19245 2391 19303 2397
rect 19334 2388 19340 2400
rect 19392 2388 19398 2440
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23256 2400 23581 2428
rect 23256 2388 23262 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 26970 2428 26976 2440
rect 26931 2400 26976 2428
rect 23569 2391 23627 2397
rect 26970 2388 26976 2400
rect 27028 2388 27034 2440
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 28408 2400 28457 2428
rect 28408 2388 28414 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29696 2400 29929 2428
rect 29696 2388 29702 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 2648 2332 3188 2360
rect 9309 2363 9367 2369
rect 2648 2320 2654 2332
rect 9309 2329 9321 2363
rect 9355 2360 9367 2363
rect 10502 2360 10508 2372
rect 9355 2332 10508 2360
rect 9355 2329 9367 2332
rect 9309 2323 9367 2329
rect 10502 2320 10508 2332
rect 10560 2320 10566 2372
rect 15470 2320 15476 2372
rect 15528 2360 15534 2372
rect 15657 2363 15715 2369
rect 15657 2360 15669 2363
rect 15528 2332 15669 2360
rect 15528 2320 15534 2332
rect 15657 2329 15669 2332
rect 15703 2329 15715 2363
rect 15657 2323 15715 2329
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 20809 2363 20867 2369
rect 20809 2360 20821 2363
rect 20680 2332 20821 2360
rect 20680 2320 20686 2332
rect 20809 2329 20821 2332
rect 20855 2329 20867 2363
rect 20809 2323 20867 2329
rect 21910 2320 21916 2372
rect 21968 2360 21974 2372
rect 22281 2363 22339 2369
rect 22281 2360 22293 2363
rect 21968 2332 22293 2360
rect 21968 2320 21974 2332
rect 22281 2329 22293 2332
rect 22327 2329 22339 2363
rect 22281 2323 22339 2329
rect 24486 2320 24492 2372
rect 24544 2360 24550 2372
rect 24857 2363 24915 2369
rect 24857 2360 24869 2363
rect 24544 2332 24869 2360
rect 24544 2320 24550 2332
rect 24857 2329 24869 2332
rect 24903 2329 24915 2363
rect 24857 2323 24915 2329
rect 26237 2363 26295 2369
rect 26237 2329 26249 2363
rect 26283 2360 26295 2363
rect 27062 2360 27068 2372
rect 26283 2332 27068 2360
rect 26283 2329 26295 2332
rect 26237 2323 26295 2329
rect 27062 2320 27068 2332
rect 27120 2320 27126 2372
rect 5261 2295 5319 2301
rect 5261 2261 5273 2295
rect 5307 2292 5319 2295
rect 11974 2292 11980 2304
rect 5307 2264 11980 2292
rect 5307 2261 5319 2264
rect 5261 2255 5319 2261
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 14921 2295 14979 2301
rect 14921 2261 14933 2295
rect 14967 2292 14979 2295
rect 15562 2292 15568 2304
rect 14967 2264 15568 2292
rect 14967 2261 14979 2264
rect 14921 2255 14979 2261
rect 15562 2252 15568 2264
rect 15620 2252 15626 2304
rect 15746 2292 15752 2304
rect 15707 2264 15752 2292
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2292 16911 2295
rect 21726 2292 21732 2304
rect 16899 2264 21732 2292
rect 16899 2261 16911 2264
rect 16853 2255 16911 2261
rect 21726 2252 21732 2264
rect 21784 2252 21790 2304
rect 27338 2252 27344 2304
rect 27396 2292 27402 2304
rect 28629 2295 28687 2301
rect 28629 2292 28641 2295
rect 27396 2264 28641 2292
rect 27396 2252 27402 2264
rect 28629 2261 28641 2264
rect 28675 2261 28687 2295
rect 29730 2292 29736 2304
rect 29691 2264 29736 2292
rect 28629 2255 28687 2261
rect 29730 2252 29736 2264
rect 29788 2252 29794 2304
rect 32490 2252 32496 2304
rect 32548 2292 32554 2304
rect 36004 2292 36032 2468
rect 40313 2465 40325 2499
rect 40359 2496 40371 2499
rect 40678 2496 40684 2508
rect 40359 2468 40684 2496
rect 40359 2465 40371 2468
rect 40313 2459 40371 2465
rect 40678 2456 40684 2468
rect 40736 2456 40742 2508
rect 42518 2456 42524 2508
rect 42576 2496 42582 2508
rect 46477 2499 46535 2505
rect 46477 2496 46489 2499
rect 42576 2468 46489 2496
rect 42576 2456 42582 2468
rect 46477 2465 46489 2468
rect 46523 2465 46535 2499
rect 46477 2459 46535 2465
rect 38010 2388 38016 2440
rect 38068 2428 38074 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 38068 2400 38117 2428
rect 38068 2388 38074 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 38194 2388 38200 2440
rect 38252 2428 38258 2440
rect 40034 2428 40040 2440
rect 38252 2400 39436 2428
rect 39995 2400 40040 2428
rect 38252 2388 38258 2400
rect 36078 2320 36084 2372
rect 36136 2360 36142 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 36136 2332 36277 2360
rect 36136 2320 36142 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 36265 2323 36323 2329
rect 39117 2363 39175 2369
rect 39117 2329 39129 2363
rect 39163 2360 39175 2363
rect 39298 2360 39304 2372
rect 39163 2332 39304 2360
rect 39163 2329 39175 2332
rect 39117 2323 39175 2329
rect 39298 2320 39304 2332
rect 39356 2320 39362 2372
rect 39408 2360 39436 2400
rect 40034 2388 40040 2400
rect 40092 2388 40098 2440
rect 40586 2388 40592 2440
rect 40644 2428 40650 2440
rect 41141 2431 41199 2437
rect 41141 2428 41153 2431
rect 40644 2400 41153 2428
rect 40644 2388 40650 2400
rect 41141 2397 41153 2400
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 43625 2431 43683 2437
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43806 2428 43812 2440
rect 43671 2400 43812 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 43901 2431 43959 2437
rect 43901 2397 43913 2431
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 46201 2431 46259 2437
rect 46201 2397 46213 2431
rect 46247 2428 46259 2431
rect 47026 2428 47032 2440
rect 46247 2400 47032 2428
rect 46247 2397 46259 2400
rect 46201 2391 46259 2397
rect 43916 2360 43944 2391
rect 47026 2388 47032 2400
rect 47084 2388 47090 2440
rect 39408 2332 43944 2360
rect 45373 2363 45431 2369
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46382 2360 46388 2372
rect 45419 2332 46388 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46382 2320 46388 2332
rect 46440 2320 46446 2372
rect 47765 2363 47823 2369
rect 47765 2329 47777 2363
rect 47811 2360 47823 2363
rect 48038 2360 48044 2372
rect 47811 2332 48044 2360
rect 47811 2329 47823 2332
rect 47765 2323 47823 2329
rect 48038 2320 48044 2332
rect 48096 2320 48102 2372
rect 45462 2292 45468 2304
rect 32548 2264 36032 2292
rect 45423 2264 45468 2292
rect 32548 2252 32554 2264
rect 45462 2252 45468 2264
rect 45520 2252 45526 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 4062 2048 4068 2100
rect 4120 2088 4126 2100
rect 10042 2088 10048 2100
rect 4120 2060 10048 2088
rect 4120 2048 4126 2060
rect 10042 2048 10048 2060
rect 10100 2048 10106 2100
rect 21174 1980 21180 2032
rect 21232 2020 21238 2032
rect 45462 2020 45468 2032
rect 21232 1992 45468 2020
rect 21232 1980 21238 1992
rect 45462 1980 45468 1992
rect 45520 1980 45526 2032
rect 15746 1912 15752 1964
rect 15804 1952 15810 1964
rect 37366 1952 37372 1964
rect 15804 1924 37372 1952
rect 15804 1912 15810 1924
rect 37366 1912 37372 1924
rect 37424 1912 37430 1964
rect 29730 1844 29736 1896
rect 29788 1884 29794 1896
rect 41414 1884 41420 1896
rect 29788 1856 41420 1884
rect 29788 1844 29794 1856
rect 41414 1844 41420 1856
rect 41472 1844 41478 1896
<< via1 >>
rect 18604 47404 18656 47456
rect 22560 47404 22612 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 17224 47200 17276 47252
rect 20812 47200 20864 47252
rect 22560 47200 22612 47252
rect 12256 47064 12308 47116
rect 19248 47064 19300 47116
rect 30104 47132 30156 47184
rect 34796 47132 34848 47184
rect 47400 47132 47452 47184
rect 30748 47107 30800 47116
rect 30748 47073 30757 47107
rect 30757 47073 30791 47107
rect 30791 47073 30800 47107
rect 30748 47064 30800 47073
rect 1952 46996 2004 47048
rect 3240 46996 3292 47048
rect 4712 47039 4764 47048
rect 4712 47005 4721 47039
rect 4721 47005 4755 47039
rect 4755 47005 4764 47039
rect 4712 46996 4764 47005
rect 5816 46996 5868 47048
rect 7288 47039 7340 47048
rect 7288 47005 7297 47039
rect 7297 47005 7331 47039
rect 7331 47005 7340 47039
rect 7288 46996 7340 47005
rect 9036 46996 9088 47048
rect 2044 46971 2096 46980
rect 2044 46937 2053 46971
rect 2053 46937 2087 46971
rect 2087 46937 2096 46971
rect 2044 46928 2096 46937
rect 4068 46971 4120 46980
rect 2596 46860 2648 46912
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 4988 46971 5040 46980
rect 4988 46937 4997 46971
rect 4997 46937 5031 46971
rect 5031 46937 5040 46971
rect 4988 46928 5040 46937
rect 6644 46971 6696 46980
rect 6644 46937 6653 46971
rect 6653 46937 6687 46971
rect 6687 46937 6696 46971
rect 6644 46928 6696 46937
rect 9496 46928 9548 46980
rect 7472 46903 7524 46912
rect 7472 46869 7481 46903
rect 7481 46869 7515 46903
rect 7515 46869 7524 46903
rect 7472 46860 7524 46869
rect 12900 46860 12952 46912
rect 14188 46996 14240 47048
rect 16488 46996 16540 47048
rect 20168 46996 20220 47048
rect 20996 47039 21048 47048
rect 20996 47005 21005 47039
rect 21005 47005 21039 47039
rect 21039 47005 21048 47039
rect 20996 46996 21048 47005
rect 22008 47039 22060 47048
rect 22008 47005 22017 47039
rect 22017 47005 22051 47039
rect 22051 47005 22060 47039
rect 22008 46996 22060 47005
rect 24860 47039 24912 47048
rect 15016 46928 15068 46980
rect 18696 46860 18748 46912
rect 20536 46928 20588 46980
rect 24860 47005 24869 47039
rect 24869 47005 24903 47039
rect 24903 47005 24912 47039
rect 24860 46996 24912 47005
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 30840 46996 30892 47048
rect 38108 46996 38160 47048
rect 41512 47039 41564 47048
rect 41512 47005 41521 47039
rect 41521 47005 41555 47039
rect 41555 47005 41564 47039
rect 41512 46996 41564 47005
rect 42708 47039 42760 47048
rect 42708 47005 42717 47039
rect 42717 47005 42751 47039
rect 42751 47005 42760 47039
rect 42708 46996 42760 47005
rect 44456 47064 44508 47116
rect 48320 47064 48372 47116
rect 43812 46996 43864 47048
rect 45100 46996 45152 47048
rect 47676 46996 47728 47048
rect 19984 46860 20036 46912
rect 34612 46928 34664 46980
rect 39304 46860 39356 46912
rect 40408 46928 40460 46980
rect 43352 46928 43404 46980
rect 45376 46971 45428 46980
rect 45376 46937 45385 46971
rect 45385 46937 45419 46971
rect 45419 46937 45428 46971
rect 45376 46928 45428 46937
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 1860 46631 1912 46640
rect 1860 46597 1869 46631
rect 1869 46597 1903 46631
rect 1903 46597 1912 46631
rect 1860 46588 1912 46597
rect 3884 46588 3936 46640
rect 22008 46588 22060 46640
rect 24860 46588 24912 46640
rect 38108 46563 38160 46572
rect 38108 46529 38117 46563
rect 38117 46529 38151 46563
rect 38151 46529 38160 46563
rect 38108 46520 38160 46529
rect 41512 46520 41564 46572
rect 47952 46563 48004 46572
rect 47952 46529 47961 46563
rect 47961 46529 47995 46563
rect 47995 46529 48004 46563
rect 47952 46520 48004 46529
rect 3976 46495 4028 46504
rect 3976 46461 3985 46495
rect 3985 46461 4019 46495
rect 4019 46461 4028 46495
rect 3976 46452 4028 46461
rect 5172 46452 5224 46504
rect 11888 46452 11940 46504
rect 13544 46452 13596 46504
rect 14188 46452 14240 46504
rect 14280 46495 14332 46504
rect 14280 46461 14289 46495
rect 14289 46461 14323 46495
rect 14323 46461 14332 46495
rect 14280 46452 14332 46461
rect 19892 46452 19944 46504
rect 20628 46495 20680 46504
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 25136 46495 25188 46504
rect 25136 46461 25145 46495
rect 25145 46461 25179 46495
rect 25179 46461 25188 46495
rect 25136 46452 25188 46461
rect 32220 46495 32272 46504
rect 32220 46461 32229 46495
rect 32229 46461 32263 46495
rect 32263 46461 32272 46495
rect 32220 46452 32272 46461
rect 32404 46495 32456 46504
rect 32404 46461 32413 46495
rect 32413 46461 32447 46495
rect 32447 46461 32456 46495
rect 32404 46452 32456 46461
rect 38292 46495 38344 46504
rect 32312 46384 32364 46436
rect 38292 46461 38301 46495
rect 38301 46461 38335 46495
rect 38335 46461 38344 46495
rect 38292 46452 38344 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 42616 46495 42668 46504
rect 42616 46461 42625 46495
rect 42625 46461 42659 46495
rect 42659 46461 42668 46495
rect 42616 46452 42668 46461
rect 45192 46495 45244 46504
rect 41880 46384 41932 46436
rect 45192 46461 45201 46495
rect 45201 46461 45235 46495
rect 45235 46461 45244 46495
rect 45192 46452 45244 46461
rect 45652 46452 45704 46504
rect 46848 46495 46900 46504
rect 46848 46461 46857 46495
rect 46857 46461 46891 46495
rect 46891 46461 46900 46495
rect 46848 46452 46900 46461
rect 2136 46359 2188 46368
rect 2136 46325 2145 46359
rect 2145 46325 2179 46359
rect 2179 46325 2188 46359
rect 2136 46316 2188 46325
rect 10968 46316 11020 46368
rect 41052 46316 41104 46368
rect 48044 46359 48096 46368
rect 48044 46325 48053 46359
rect 48053 46325 48087 46359
rect 48087 46325 48096 46359
rect 48044 46316 48096 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3976 46112 4028 46164
rect 5172 46155 5224 46164
rect 5172 46121 5181 46155
rect 5181 46121 5215 46155
rect 5215 46121 5224 46155
rect 5172 46112 5224 46121
rect 13544 46155 13596 46164
rect 13544 46121 13553 46155
rect 13553 46121 13587 46155
rect 13587 46121 13596 46155
rect 13544 46112 13596 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 19892 46155 19944 46164
rect 19892 46121 19901 46155
rect 19901 46121 19935 46155
rect 19935 46121 19944 46155
rect 19892 46112 19944 46121
rect 24768 46112 24820 46164
rect 32220 46112 32272 46164
rect 38292 46155 38344 46164
rect 38292 46121 38301 46155
rect 38301 46121 38335 46155
rect 38335 46121 38344 46155
rect 38292 46112 38344 46121
rect 11612 45976 11664 46028
rect 20996 45976 21048 46028
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 25780 46019 25832 46028
rect 25780 45985 25789 46019
rect 25789 45985 25823 46019
rect 25823 45985 25832 46019
rect 25780 45976 25832 45985
rect 41052 46019 41104 46028
rect 41052 45985 41061 46019
rect 41061 45985 41095 46019
rect 41095 45985 41104 46019
rect 41052 45976 41104 45985
rect 42524 46019 42576 46028
rect 42524 45985 42533 46019
rect 42533 45985 42567 46019
rect 42567 45985 42576 46019
rect 42524 45976 42576 45985
rect 1768 45908 1820 45960
rect 11980 45951 12032 45960
rect 11980 45917 11989 45951
rect 11989 45917 12023 45951
rect 12023 45917 12032 45951
rect 11980 45908 12032 45917
rect 14096 45951 14148 45960
rect 14096 45917 14105 45951
rect 14105 45917 14139 45951
rect 14139 45917 14148 45951
rect 14096 45908 14148 45917
rect 20260 45908 20312 45960
rect 25228 45951 25280 45960
rect 20996 45883 21048 45892
rect 20996 45849 21005 45883
rect 21005 45849 21039 45883
rect 21039 45849 21048 45883
rect 20996 45840 21048 45849
rect 24492 45772 24544 45824
rect 25228 45917 25237 45951
rect 25237 45917 25271 45951
rect 25271 45917 25280 45951
rect 25228 45908 25280 45917
rect 38200 45951 38252 45960
rect 38200 45917 38209 45951
rect 38209 45917 38243 45951
rect 38243 45917 38252 45951
rect 38200 45908 38252 45917
rect 46848 46112 46900 46164
rect 47584 46044 47636 46096
rect 47032 46019 47084 46028
rect 47032 45985 47041 46019
rect 47041 45985 47075 46019
rect 47075 45985 47084 46019
rect 47032 45976 47084 45985
rect 45744 45908 45796 45960
rect 45836 45908 45888 45960
rect 25412 45883 25464 45892
rect 25412 45849 25421 45883
rect 25421 45849 25455 45883
rect 25455 45849 25464 45883
rect 25412 45840 25464 45849
rect 41236 45883 41288 45892
rect 41236 45849 41245 45883
rect 41245 45849 41279 45883
rect 41279 45849 41288 45883
rect 41236 45840 41288 45849
rect 38200 45772 38252 45824
rect 43444 45815 43496 45824
rect 43444 45781 43453 45815
rect 43453 45781 43487 45815
rect 43487 45781 43496 45815
rect 43444 45772 43496 45781
rect 45468 45772 45520 45824
rect 46020 45772 46072 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 11888 45611 11940 45620
rect 11888 45577 11897 45611
rect 11897 45577 11931 45611
rect 11931 45577 11940 45611
rect 11888 45568 11940 45577
rect 20996 45611 21048 45620
rect 20996 45577 21005 45611
rect 21005 45577 21039 45611
rect 21039 45577 21048 45611
rect 20996 45568 21048 45577
rect 32404 45568 32456 45620
rect 41236 45568 41288 45620
rect 42616 45568 42668 45620
rect 46388 45568 46440 45620
rect 43444 45500 43496 45552
rect 44824 45500 44876 45552
rect 1768 45475 1820 45484
rect 1768 45441 1777 45475
rect 1777 45441 1811 45475
rect 1811 45441 1820 45475
rect 1768 45432 1820 45441
rect 20904 45475 20956 45484
rect 20904 45441 20913 45475
rect 20913 45441 20947 45475
rect 20947 45441 20956 45475
rect 20904 45432 20956 45441
rect 25228 45432 25280 45484
rect 38752 45432 38804 45484
rect 40224 45432 40276 45484
rect 42708 45475 42760 45484
rect 2320 45364 2372 45416
rect 2780 45407 2832 45416
rect 2780 45373 2789 45407
rect 2789 45373 2823 45407
rect 2823 45373 2832 45407
rect 2780 45364 2832 45373
rect 42708 45441 42717 45475
rect 42717 45441 42751 45475
rect 42751 45441 42760 45475
rect 42708 45432 42760 45441
rect 43168 45407 43220 45416
rect 43168 45373 43177 45407
rect 43177 45373 43211 45407
rect 43211 45373 43220 45407
rect 43168 45364 43220 45373
rect 45008 45407 45060 45416
rect 45008 45373 45017 45407
rect 45017 45373 45051 45407
rect 45051 45373 45060 45407
rect 45008 45364 45060 45373
rect 45560 45407 45612 45416
rect 43260 45296 43312 45348
rect 45560 45373 45569 45407
rect 45569 45373 45603 45407
rect 45603 45373 45612 45407
rect 45560 45364 45612 45373
rect 46756 45228 46808 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 2320 45067 2372 45076
rect 2320 45033 2329 45067
rect 2329 45033 2363 45067
rect 2363 45033 2372 45067
rect 2320 45024 2372 45033
rect 25412 45067 25464 45076
rect 25412 45033 25421 45067
rect 25421 45033 25455 45067
rect 25455 45033 25464 45067
rect 25412 45024 25464 45033
rect 43260 45067 43312 45076
rect 43260 45033 43269 45067
rect 43269 45033 43303 45067
rect 43303 45033 43312 45067
rect 43260 45024 43312 45033
rect 45008 45024 45060 45076
rect 45192 45067 45244 45076
rect 45192 45033 45201 45067
rect 45201 45033 45235 45067
rect 45235 45033 45244 45067
rect 45192 45024 45244 45033
rect 45652 45024 45704 45076
rect 47032 44888 47084 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 3792 44820 3844 44872
rect 25320 44863 25372 44872
rect 25320 44829 25329 44863
rect 25329 44829 25363 44863
rect 25363 44829 25372 44863
rect 25320 44820 25372 44829
rect 43168 44863 43220 44872
rect 43168 44829 43177 44863
rect 43177 44829 43211 44863
rect 43211 44829 43220 44863
rect 43168 44820 43220 44829
rect 45560 44820 45612 44872
rect 47676 44752 47728 44804
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 45376 44480 45428 44532
rect 47676 44523 47728 44532
rect 47676 44489 47685 44523
rect 47685 44489 47719 44523
rect 47719 44489 47728 44523
rect 47676 44480 47728 44489
rect 45100 44387 45152 44396
rect 45100 44353 45109 44387
rect 45109 44353 45143 44387
rect 45143 44353 45152 44387
rect 45100 44344 45152 44353
rect 45836 44344 45888 44396
rect 46204 44387 46256 44396
rect 46204 44353 46213 44387
rect 46213 44353 46247 44387
rect 46247 44353 46256 44387
rect 46204 44344 46256 44353
rect 38660 44319 38712 44328
rect 38660 44285 38669 44319
rect 38669 44285 38703 44319
rect 38703 44285 38712 44319
rect 38660 44276 38712 44285
rect 38844 44319 38896 44328
rect 38844 44285 38853 44319
rect 38853 44285 38887 44319
rect 38887 44285 38896 44319
rect 38844 44276 38896 44285
rect 40040 44319 40092 44328
rect 40040 44285 40049 44319
rect 40049 44285 40083 44319
rect 40083 44285 40092 44319
rect 40040 44276 40092 44285
rect 46940 44183 46992 44192
rect 46940 44149 46949 44183
rect 46949 44149 46983 44183
rect 46983 44149 46992 44183
rect 46940 44140 46992 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 38844 43979 38896 43988
rect 38844 43945 38853 43979
rect 38853 43945 38887 43979
rect 38887 43945 38896 43979
rect 38844 43936 38896 43945
rect 46940 43800 46992 43852
rect 48228 43800 48280 43852
rect 25780 43732 25832 43784
rect 25320 43664 25372 43716
rect 38936 43732 38988 43784
rect 38660 43596 38712 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 47032 43299 47084 43308
rect 47032 43265 47041 43299
rect 47041 43265 47075 43299
rect 47075 43265 47084 43299
rect 47032 43256 47084 43265
rect 1676 43231 1728 43240
rect 1676 43197 1685 43231
rect 1685 43197 1719 43231
rect 1719 43197 1728 43231
rect 1676 43188 1728 43197
rect 47768 43095 47820 43104
rect 47768 43061 47777 43095
rect 47777 43061 47811 43095
rect 47811 43061 47820 43095
rect 47768 43052 47820 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 47768 42712 47820 42764
rect 46940 42576 46992 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 46940 42347 46992 42356
rect 46940 42313 46949 42347
rect 46949 42313 46983 42347
rect 46983 42313 46992 42347
rect 46940 42304 46992 42313
rect 46572 42168 46624 42220
rect 46848 42211 46900 42220
rect 46848 42177 46857 42211
rect 46857 42177 46891 42211
rect 46891 42177 46900 42211
rect 46848 42168 46900 42177
rect 47584 42211 47636 42220
rect 47584 42177 47593 42211
rect 47593 42177 47627 42211
rect 47627 42177 47636 42211
rect 47584 42168 47636 42177
rect 1400 41964 1452 42016
rect 46480 41964 46532 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 46480 41667 46532 41676
rect 46480 41633 46489 41667
rect 46489 41633 46523 41667
rect 46523 41633 46532 41667
rect 46480 41624 46532 41633
rect 48136 41599 48188 41608
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 48136 41565 48145 41599
rect 48145 41565 48179 41599
rect 48179 41565 48188 41599
rect 48136 41556 48188 41565
rect 47676 41488 47728 41540
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 14096 41080 14148 41132
rect 47952 41123 48004 41132
rect 47952 41089 47961 41123
rect 47961 41089 47995 41123
rect 47995 41089 48004 41123
rect 47952 41080 48004 41089
rect 47492 40876 47544 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47676 40715 47728 40724
rect 47676 40681 47685 40715
rect 47685 40681 47719 40715
rect 47719 40681 47728 40715
rect 47676 40672 47728 40681
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 1952 40375 2004 40384
rect 1952 40341 1961 40375
rect 1961 40341 1995 40375
rect 1995 40341 2004 40375
rect 1952 40332 2004 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 46756 40035 46808 40044
rect 46756 40001 46765 40035
rect 46765 40001 46799 40035
rect 46799 40001 46808 40035
rect 46756 39992 46808 40001
rect 46480 39788 46532 39840
rect 47768 39831 47820 39840
rect 47768 39797 47777 39831
rect 47777 39797 47811 39831
rect 47811 39797 47820 39831
rect 47768 39788 47820 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 20352 39448 20404 39500
rect 47768 39516 47820 39568
rect 46480 39491 46532 39500
rect 46480 39457 46489 39491
rect 46489 39457 46523 39491
rect 46523 39457 46532 39491
rect 46480 39448 46532 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 22100 39244 22152 39296
rect 24584 39312 24636 39364
rect 46020 39244 46072 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 24584 39083 24636 39092
rect 24584 39049 24593 39083
rect 24593 39049 24627 39083
rect 24627 39049 24636 39083
rect 24584 39040 24636 39049
rect 20812 38972 20864 39024
rect 22100 39015 22152 39024
rect 22100 38981 22109 39015
rect 22109 38981 22143 39015
rect 22143 38981 22152 39015
rect 22100 38972 22152 38981
rect 22560 38972 22612 39024
rect 20352 38904 20404 38956
rect 20536 38836 20588 38888
rect 24676 38904 24728 38956
rect 24124 38879 24176 38888
rect 24124 38845 24133 38879
rect 24133 38845 24167 38879
rect 24167 38845 24176 38879
rect 24124 38836 24176 38845
rect 19064 38700 19116 38752
rect 38660 38700 38712 38752
rect 47860 38947 47912 38956
rect 47860 38913 47869 38947
rect 47869 38913 47903 38947
rect 47903 38913 47912 38947
rect 47860 38904 47912 38913
rect 39856 38836 39908 38888
rect 46204 38836 46256 38888
rect 41144 38768 41196 38820
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 9496 38360 9548 38412
rect 21364 38496 21416 38548
rect 22560 38496 22612 38548
rect 38936 38496 38988 38548
rect 46756 38496 46808 38548
rect 18144 38428 18196 38480
rect 19248 38335 19300 38344
rect 19248 38301 19257 38335
rect 19257 38301 19291 38335
rect 19291 38301 19300 38335
rect 19248 38292 19300 38301
rect 22836 38292 22888 38344
rect 26976 38360 27028 38412
rect 40684 38403 40736 38412
rect 40684 38369 40693 38403
rect 40693 38369 40727 38403
rect 40727 38369 40736 38403
rect 40684 38360 40736 38369
rect 43168 38360 43220 38412
rect 24492 38292 24544 38344
rect 38660 38335 38712 38344
rect 38660 38301 38669 38335
rect 38669 38301 38703 38335
rect 38703 38301 38712 38335
rect 38660 38292 38712 38301
rect 46296 38335 46348 38344
rect 46296 38301 46305 38335
rect 46305 38301 46339 38335
rect 46339 38301 46348 38335
rect 46296 38292 46348 38301
rect 23204 38224 23256 38276
rect 19340 38199 19392 38208
rect 19340 38165 19349 38199
rect 19349 38165 19383 38199
rect 19383 38165 19392 38199
rect 19340 38156 19392 38165
rect 20812 38199 20864 38208
rect 20812 38165 20821 38199
rect 20821 38165 20855 38199
rect 20855 38165 20864 38199
rect 20812 38156 20864 38165
rect 24492 38199 24544 38208
rect 24492 38165 24501 38199
rect 24501 38165 24535 38199
rect 24535 38165 24544 38199
rect 24492 38156 24544 38165
rect 46848 38224 46900 38276
rect 48136 38267 48188 38276
rect 48136 38233 48145 38267
rect 48145 38233 48179 38267
rect 48179 38233 48188 38267
rect 48136 38224 48188 38233
rect 47308 38156 47360 38208
rect 47584 38156 47636 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 17224 37816 17276 37868
rect 22376 37952 22428 38004
rect 46848 37995 46900 38004
rect 19800 37927 19852 37936
rect 19800 37893 19809 37927
rect 19809 37893 19843 37927
rect 19843 37893 19852 37927
rect 19800 37884 19852 37893
rect 20812 37884 20864 37936
rect 24492 37884 24544 37936
rect 46848 37961 46857 37995
rect 46857 37961 46891 37995
rect 46891 37961 46900 37995
rect 46848 37952 46900 37961
rect 19432 37748 19484 37800
rect 20536 37748 20588 37800
rect 26976 37859 27028 37868
rect 26976 37825 26985 37859
rect 26985 37825 27019 37859
rect 27019 37825 27028 37859
rect 26976 37816 27028 37825
rect 30656 37816 30708 37868
rect 38660 37884 38712 37936
rect 39948 37884 40000 37936
rect 40224 37927 40276 37936
rect 40224 37893 40233 37927
rect 40233 37893 40267 37927
rect 40267 37893 40276 37927
rect 40224 37884 40276 37893
rect 46296 37884 46348 37936
rect 38752 37859 38804 37868
rect 38752 37825 38761 37859
rect 38761 37825 38795 37859
rect 38795 37825 38804 37859
rect 38752 37816 38804 37825
rect 46756 37859 46808 37868
rect 46756 37825 46765 37859
rect 46765 37825 46799 37859
rect 46799 37825 46808 37859
rect 46756 37816 46808 37825
rect 22744 37791 22796 37800
rect 22744 37757 22753 37791
rect 22753 37757 22787 37791
rect 22787 37757 22796 37791
rect 22744 37748 22796 37757
rect 24952 37791 25004 37800
rect 24952 37757 24961 37791
rect 24961 37757 24995 37791
rect 24995 37757 25004 37791
rect 24952 37748 25004 37757
rect 18144 37655 18196 37664
rect 18144 37621 18153 37655
rect 18153 37621 18187 37655
rect 18187 37621 18196 37655
rect 18144 37612 18196 37621
rect 21180 37612 21232 37664
rect 22192 37612 22244 37664
rect 22376 37612 22428 37664
rect 22836 37612 22888 37664
rect 24400 37612 24452 37664
rect 25504 37612 25556 37664
rect 27620 37612 27672 37664
rect 29460 37655 29512 37664
rect 29460 37621 29469 37655
rect 29469 37621 29503 37655
rect 29503 37621 29512 37655
rect 29460 37612 29512 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 18604 37451 18656 37460
rect 18604 37417 18613 37451
rect 18613 37417 18647 37451
rect 18647 37417 18656 37451
rect 18604 37408 18656 37417
rect 19800 37408 19852 37460
rect 22744 37408 22796 37460
rect 24400 37451 24452 37460
rect 24400 37417 24409 37451
rect 24409 37417 24443 37451
rect 24443 37417 24452 37451
rect 24400 37408 24452 37417
rect 20168 37340 20220 37392
rect 21180 37315 21232 37324
rect 21180 37281 21189 37315
rect 21189 37281 21223 37315
rect 21223 37281 21232 37315
rect 21180 37272 21232 37281
rect 21364 37340 21416 37392
rect 23204 37315 23256 37324
rect 23204 37281 23213 37315
rect 23213 37281 23247 37315
rect 23247 37281 23256 37315
rect 23204 37272 23256 37281
rect 29920 37272 29972 37324
rect 1768 37204 1820 37256
rect 18328 37247 18380 37256
rect 18328 37213 18337 37247
rect 18337 37213 18371 37247
rect 18371 37213 18380 37247
rect 18328 37204 18380 37213
rect 18696 37247 18748 37256
rect 18696 37213 18705 37247
rect 18705 37213 18739 37247
rect 18739 37213 18748 37247
rect 18696 37204 18748 37213
rect 20996 37204 21048 37256
rect 18604 37136 18656 37188
rect 21916 37204 21968 37256
rect 23020 37247 23072 37256
rect 23020 37213 23029 37247
rect 23029 37213 23063 37247
rect 23063 37213 23072 37247
rect 23020 37204 23072 37213
rect 24676 37247 24728 37256
rect 22560 37136 22612 37188
rect 24676 37213 24685 37247
rect 24685 37213 24719 37247
rect 24719 37213 24728 37247
rect 24676 37204 24728 37213
rect 24768 37204 24820 37256
rect 18512 37068 18564 37120
rect 19340 37068 19392 37120
rect 24308 37136 24360 37188
rect 24124 37068 24176 37120
rect 24860 37111 24912 37120
rect 24860 37077 24869 37111
rect 24869 37077 24903 37111
rect 24903 37077 24912 37111
rect 24860 37068 24912 37077
rect 26240 37179 26292 37188
rect 26240 37145 26249 37179
rect 26249 37145 26283 37179
rect 26283 37145 26292 37179
rect 26240 37136 26292 37145
rect 27620 37136 27672 37188
rect 28540 37204 28592 37256
rect 28724 37247 28776 37256
rect 28724 37213 28733 37247
rect 28733 37213 28767 37247
rect 28767 37213 28776 37247
rect 28724 37204 28776 37213
rect 29644 37204 29696 37256
rect 27528 37068 27580 37120
rect 27712 37111 27764 37120
rect 27712 37077 27721 37111
rect 27721 37077 27755 37111
rect 27755 37077 27764 37111
rect 27712 37068 27764 37077
rect 28448 37068 28500 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 26240 36907 26292 36916
rect 26240 36873 26249 36907
rect 26249 36873 26283 36907
rect 26283 36873 26292 36907
rect 26240 36864 26292 36873
rect 17960 36796 18012 36848
rect 21732 36796 21784 36848
rect 21916 36796 21968 36848
rect 28724 36864 28776 36916
rect 28448 36839 28500 36848
rect 28448 36805 28457 36839
rect 28457 36805 28491 36839
rect 28491 36805 28500 36839
rect 28448 36796 28500 36805
rect 29460 36796 29512 36848
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 24308 36728 24360 36780
rect 25504 36728 25556 36780
rect 26240 36728 26292 36780
rect 27528 36728 27580 36780
rect 30656 36771 30708 36780
rect 30656 36737 30665 36771
rect 30665 36737 30699 36771
rect 30699 36737 30708 36771
rect 30656 36728 30708 36737
rect 2228 36660 2280 36712
rect 2780 36703 2832 36712
rect 2780 36669 2789 36703
rect 2789 36669 2823 36703
rect 2823 36669 2832 36703
rect 2780 36660 2832 36669
rect 16672 36703 16724 36712
rect 16672 36669 16681 36703
rect 16681 36669 16715 36703
rect 16715 36669 16724 36703
rect 16672 36660 16724 36669
rect 18236 36660 18288 36712
rect 16672 36524 16724 36576
rect 19432 36660 19484 36712
rect 19800 36703 19852 36712
rect 19800 36669 19809 36703
rect 19809 36669 19843 36703
rect 19843 36669 19852 36703
rect 19800 36660 19852 36669
rect 18604 36524 18656 36576
rect 21272 36567 21324 36576
rect 21272 36533 21281 36567
rect 21281 36533 21315 36567
rect 21315 36533 21324 36567
rect 21272 36524 21324 36533
rect 25596 36524 25648 36576
rect 29920 36567 29972 36576
rect 29920 36533 29929 36567
rect 29929 36533 29963 36567
rect 29963 36533 29972 36567
rect 29920 36524 29972 36533
rect 30748 36567 30800 36576
rect 30748 36533 30757 36567
rect 30757 36533 30791 36567
rect 30791 36533 30800 36567
rect 30748 36524 30800 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2228 36363 2280 36372
rect 2228 36329 2237 36363
rect 2237 36329 2271 36363
rect 2271 36329 2280 36363
rect 2228 36320 2280 36329
rect 19800 36320 19852 36372
rect 21732 36363 21784 36372
rect 21732 36329 21741 36363
rect 21741 36329 21775 36363
rect 21775 36329 21784 36363
rect 21732 36320 21784 36329
rect 23020 36320 23072 36372
rect 24952 36320 25004 36372
rect 28540 36320 28592 36372
rect 2412 36116 2464 36168
rect 40684 36252 40736 36304
rect 17500 36227 17552 36236
rect 17500 36193 17509 36227
rect 17509 36193 17543 36227
rect 17543 36193 17552 36227
rect 17500 36184 17552 36193
rect 18236 36227 18288 36236
rect 18236 36193 18245 36227
rect 18245 36193 18279 36227
rect 18279 36193 18288 36227
rect 18236 36184 18288 36193
rect 18604 36184 18656 36236
rect 18512 36116 18564 36168
rect 19432 36116 19484 36168
rect 22652 36184 22704 36236
rect 24400 36184 24452 36236
rect 21088 36159 21140 36168
rect 21088 36125 21097 36159
rect 21097 36125 21131 36159
rect 21131 36125 21140 36159
rect 21088 36116 21140 36125
rect 11980 36048 12032 36100
rect 21456 36116 21508 36168
rect 23480 36116 23532 36168
rect 24584 36116 24636 36168
rect 27344 36184 27396 36236
rect 27436 36184 27488 36236
rect 25320 36116 25372 36168
rect 25504 36116 25556 36168
rect 25964 36116 26016 36168
rect 26700 36116 26752 36168
rect 27896 36116 27948 36168
rect 29000 36159 29052 36168
rect 29000 36125 29009 36159
rect 29009 36125 29043 36159
rect 29043 36125 29052 36159
rect 29000 36116 29052 36125
rect 29920 36116 29972 36168
rect 18328 35980 18380 36032
rect 29092 36048 29144 36100
rect 29644 36048 29696 36100
rect 22560 36023 22612 36032
rect 22560 35989 22569 36023
rect 22569 35989 22603 36023
rect 22603 35989 22612 36023
rect 22560 35980 22612 35989
rect 26608 35980 26660 36032
rect 27712 35980 27764 36032
rect 29460 35980 29512 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 17960 35776 18012 35828
rect 18696 35776 18748 35828
rect 22652 35819 22704 35828
rect 21272 35708 21324 35760
rect 22652 35785 22661 35819
rect 22661 35785 22695 35819
rect 22695 35785 22704 35819
rect 22652 35776 22704 35785
rect 24124 35776 24176 35828
rect 24492 35776 24544 35828
rect 31024 35776 31076 35828
rect 23204 35708 23256 35760
rect 26792 35708 26844 35760
rect 27528 35708 27580 35760
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 15936 35640 15988 35692
rect 19340 35640 19392 35692
rect 21824 35640 21876 35692
rect 22008 35572 22060 35624
rect 23480 35640 23532 35692
rect 24400 35683 24452 35692
rect 24400 35649 24409 35683
rect 24409 35649 24443 35683
rect 24443 35649 24452 35683
rect 24400 35640 24452 35649
rect 24584 35683 24636 35692
rect 24584 35649 24593 35683
rect 24593 35649 24627 35683
rect 24627 35649 24636 35683
rect 24584 35640 24636 35649
rect 26516 35640 26568 35692
rect 27436 35683 27488 35692
rect 27436 35649 27445 35683
rect 27445 35649 27479 35683
rect 27479 35649 27488 35683
rect 27436 35640 27488 35649
rect 28172 35683 28224 35692
rect 28172 35649 28181 35683
rect 28181 35649 28215 35683
rect 28215 35649 28224 35683
rect 28172 35640 28224 35649
rect 20536 35504 20588 35556
rect 24952 35572 25004 35624
rect 25688 35615 25740 35624
rect 25688 35581 25697 35615
rect 25697 35581 25731 35615
rect 25731 35581 25740 35615
rect 25688 35572 25740 35581
rect 26240 35572 26292 35624
rect 2136 35436 2188 35488
rect 25320 35504 25372 35556
rect 26332 35504 26384 35556
rect 27344 35504 27396 35556
rect 29092 35683 29144 35692
rect 29092 35649 29101 35683
rect 29101 35649 29135 35683
rect 29135 35649 29144 35683
rect 29092 35640 29144 35649
rect 30748 35708 30800 35760
rect 48136 35683 48188 35692
rect 48136 35649 48145 35683
rect 48145 35649 48179 35683
rect 48179 35649 48188 35683
rect 48136 35640 48188 35649
rect 28632 35572 28684 35624
rect 30748 35572 30800 35624
rect 24400 35436 24452 35488
rect 26148 35436 26200 35488
rect 28264 35479 28316 35488
rect 28264 35445 28273 35479
rect 28273 35445 28307 35479
rect 28307 35445 28316 35479
rect 28264 35436 28316 35445
rect 28448 35436 28500 35488
rect 30564 35436 30616 35488
rect 47124 35436 47176 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 21824 35275 21876 35284
rect 21824 35241 21833 35275
rect 21833 35241 21867 35275
rect 21867 35241 21876 35275
rect 21824 35232 21876 35241
rect 26332 35275 26384 35284
rect 26332 35241 26341 35275
rect 26341 35241 26375 35275
rect 26375 35241 26384 35275
rect 26332 35232 26384 35241
rect 28448 35232 28500 35284
rect 29000 35232 29052 35284
rect 30748 35232 30800 35284
rect 24768 35164 24820 35216
rect 19432 35096 19484 35148
rect 20168 35096 20220 35148
rect 22100 35096 22152 35148
rect 26608 35164 26660 35216
rect 28264 35164 28316 35216
rect 28908 35164 28960 35216
rect 25596 35139 25648 35148
rect 25596 35105 25605 35139
rect 25605 35105 25639 35139
rect 25639 35105 25648 35139
rect 25596 35096 25648 35105
rect 27252 35096 27304 35148
rect 28632 35139 28684 35148
rect 28632 35105 28641 35139
rect 28641 35105 28675 35139
rect 28675 35105 28684 35139
rect 28632 35096 28684 35105
rect 30564 35139 30616 35148
rect 16856 35071 16908 35080
rect 16856 35037 16865 35071
rect 16865 35037 16899 35071
rect 16899 35037 16908 35071
rect 16856 35028 16908 35037
rect 17040 35071 17092 35080
rect 17040 35037 17049 35071
rect 17049 35037 17083 35071
rect 17083 35037 17092 35071
rect 17040 35028 17092 35037
rect 19340 35071 19392 35080
rect 19340 35037 19349 35071
rect 19349 35037 19383 35071
rect 19383 35037 19392 35071
rect 19340 35028 19392 35037
rect 20352 35028 20404 35080
rect 21272 35028 21324 35080
rect 24860 35028 24912 35080
rect 25136 35028 25188 35080
rect 26332 35028 26384 35080
rect 26516 35071 26568 35080
rect 26516 35037 26525 35071
rect 26525 35037 26559 35071
rect 26559 35037 26568 35071
rect 26516 35028 26568 35037
rect 26608 35071 26660 35080
rect 26608 35037 26617 35071
rect 26617 35037 26651 35071
rect 26651 35037 26660 35071
rect 26884 35071 26936 35080
rect 26608 35028 26660 35037
rect 26884 35037 26893 35071
rect 26893 35037 26927 35071
rect 26927 35037 26936 35071
rect 26884 35028 26936 35037
rect 27712 35071 27764 35080
rect 27712 35037 27721 35071
rect 27721 35037 27755 35071
rect 27755 35037 27764 35071
rect 27712 35028 27764 35037
rect 30564 35105 30573 35139
rect 30573 35105 30607 35139
rect 30607 35105 30616 35139
rect 30564 35096 30616 35105
rect 30932 35096 30984 35148
rect 20812 34960 20864 35012
rect 21456 34960 21508 35012
rect 24032 34960 24084 35012
rect 16764 34892 16816 34944
rect 19432 34935 19484 34944
rect 19432 34901 19441 34935
rect 19441 34901 19475 34935
rect 19475 34901 19484 34935
rect 19432 34892 19484 34901
rect 20536 34892 20588 34944
rect 22376 34892 22428 34944
rect 25872 34935 25924 34944
rect 25872 34901 25881 34935
rect 25881 34901 25915 34935
rect 25915 34901 25924 34935
rect 25872 34892 25924 34901
rect 27436 34892 27488 34944
rect 28172 34960 28224 35012
rect 28540 35003 28592 35012
rect 28540 34969 28549 35003
rect 28549 34969 28583 35003
rect 28583 34969 28592 35003
rect 28540 34960 28592 34969
rect 29000 35028 29052 35080
rect 30288 35071 30340 35080
rect 30288 35037 30297 35071
rect 30297 35037 30331 35071
rect 30331 35037 30340 35071
rect 30288 35028 30340 35037
rect 29828 34960 29880 35012
rect 31024 35028 31076 35080
rect 48228 35028 48280 35080
rect 28724 34892 28776 34944
rect 47860 34892 47912 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 16856 34688 16908 34740
rect 15936 34595 15988 34604
rect 15936 34561 15945 34595
rect 15945 34561 15979 34595
rect 15979 34561 15988 34595
rect 15936 34552 15988 34561
rect 18328 34688 18380 34740
rect 21088 34688 21140 34740
rect 24400 34688 24452 34740
rect 24584 34688 24636 34740
rect 25228 34688 25280 34740
rect 25596 34688 25648 34740
rect 27712 34731 27764 34740
rect 27712 34697 27721 34731
rect 27721 34697 27755 34731
rect 27755 34697 27764 34731
rect 27712 34688 27764 34697
rect 18696 34620 18748 34672
rect 19432 34620 19484 34672
rect 22100 34620 22152 34672
rect 23388 34620 23440 34672
rect 24032 34663 24084 34672
rect 24032 34629 24041 34663
rect 24041 34629 24075 34663
rect 24075 34629 24084 34663
rect 24032 34620 24084 34629
rect 25136 34620 25188 34672
rect 20904 34595 20956 34604
rect 16580 34484 16632 34536
rect 17316 34484 17368 34536
rect 17592 34484 17644 34536
rect 18420 34527 18472 34536
rect 18420 34493 18429 34527
rect 18429 34493 18463 34527
rect 18463 34493 18472 34527
rect 18420 34484 18472 34493
rect 20904 34561 20913 34595
rect 20913 34561 20947 34595
rect 20947 34561 20956 34595
rect 20904 34552 20956 34561
rect 22192 34595 22244 34604
rect 22192 34561 22201 34595
rect 22201 34561 22235 34595
rect 22235 34561 22244 34595
rect 22192 34552 22244 34561
rect 22376 34595 22428 34604
rect 22376 34561 22385 34595
rect 22385 34561 22419 34595
rect 22419 34561 22428 34595
rect 22376 34552 22428 34561
rect 22928 34595 22980 34604
rect 22928 34561 22937 34595
rect 22937 34561 22971 34595
rect 22971 34561 22980 34595
rect 22928 34552 22980 34561
rect 21272 34484 21324 34536
rect 23664 34552 23716 34604
rect 24768 34552 24820 34604
rect 26332 34620 26384 34672
rect 26700 34620 26752 34672
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 25504 34595 25556 34604
rect 25504 34561 25539 34595
rect 25539 34561 25556 34595
rect 25504 34552 25556 34561
rect 25964 34552 26016 34604
rect 23572 34484 23624 34536
rect 23480 34416 23532 34468
rect 26056 34484 26108 34536
rect 26884 34552 26936 34604
rect 27344 34552 27396 34604
rect 28632 34620 28684 34672
rect 30288 34688 30340 34740
rect 26332 34484 26384 34536
rect 26792 34484 26844 34536
rect 28724 34595 28776 34604
rect 28724 34561 28733 34595
rect 28733 34561 28767 34595
rect 28767 34561 28776 34595
rect 28724 34552 28776 34561
rect 28908 34595 28960 34604
rect 28908 34561 28917 34595
rect 28917 34561 28951 34595
rect 28951 34561 28960 34595
rect 28908 34552 28960 34561
rect 28816 34484 28868 34536
rect 29460 34552 29512 34604
rect 30564 34620 30616 34672
rect 29920 34595 29972 34604
rect 29920 34561 29929 34595
rect 29929 34561 29963 34595
rect 29963 34561 29972 34595
rect 47768 34595 47820 34604
rect 29920 34552 29972 34561
rect 47768 34561 47777 34595
rect 47777 34561 47811 34595
rect 47811 34561 47820 34595
rect 47768 34552 47820 34561
rect 19984 34348 20036 34400
rect 20720 34391 20772 34400
rect 20720 34357 20729 34391
rect 20729 34357 20763 34391
rect 20763 34357 20772 34391
rect 20720 34348 20772 34357
rect 21456 34348 21508 34400
rect 24308 34391 24360 34400
rect 24308 34357 24317 34391
rect 24317 34357 24351 34391
rect 24351 34357 24360 34391
rect 24308 34348 24360 34357
rect 25964 34416 26016 34468
rect 30380 34348 30432 34400
rect 47216 34348 47268 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19984 34187 20036 34196
rect 1952 34008 2004 34060
rect 16672 34008 16724 34060
rect 18420 34008 18472 34060
rect 19340 34008 19392 34060
rect 19984 34153 19993 34187
rect 19993 34153 20027 34187
rect 20027 34153 20036 34187
rect 19984 34144 20036 34153
rect 21456 34187 21508 34196
rect 21456 34153 21465 34187
rect 21465 34153 21499 34187
rect 21499 34153 21508 34187
rect 21456 34144 21508 34153
rect 23388 34144 23440 34196
rect 23664 34187 23716 34196
rect 23664 34153 23673 34187
rect 23673 34153 23707 34187
rect 23707 34153 23716 34187
rect 23664 34144 23716 34153
rect 24584 34144 24636 34196
rect 25688 34144 25740 34196
rect 28632 34144 28684 34196
rect 20996 34076 21048 34128
rect 1584 33983 1636 33992
rect 1584 33949 1593 33983
rect 1593 33949 1627 33983
rect 1627 33949 1636 33983
rect 1584 33940 1636 33949
rect 19248 33983 19300 33992
rect 19248 33949 19257 33983
rect 19257 33949 19291 33983
rect 19291 33949 19300 33983
rect 19248 33940 19300 33949
rect 20904 34008 20956 34060
rect 1952 33804 2004 33856
rect 16580 33872 16632 33924
rect 20536 33940 20588 33992
rect 21088 33983 21140 33992
rect 21088 33949 21097 33983
rect 21097 33949 21131 33983
rect 21131 33949 21140 33983
rect 21088 33940 21140 33949
rect 21364 33983 21416 33992
rect 21364 33949 21373 33983
rect 21373 33949 21407 33983
rect 21407 33949 21416 33983
rect 21364 33940 21416 33949
rect 22376 34076 22428 34128
rect 22192 34008 22244 34060
rect 22928 34008 22980 34060
rect 27528 34008 27580 34060
rect 47124 34051 47176 34060
rect 47124 34017 47133 34051
rect 47133 34017 47167 34051
rect 47167 34017 47176 34051
rect 47124 34008 47176 34017
rect 47676 34051 47728 34060
rect 47676 34017 47685 34051
rect 47685 34017 47719 34051
rect 47719 34017 47728 34051
rect 47676 34008 47728 34017
rect 22376 33983 22428 33992
rect 22376 33949 22385 33983
rect 22385 33949 22419 33983
rect 22419 33949 22428 33983
rect 22376 33940 22428 33949
rect 23572 33983 23624 33992
rect 23572 33949 23581 33983
rect 23581 33949 23615 33983
rect 23615 33949 23624 33983
rect 23572 33940 23624 33949
rect 20076 33872 20128 33924
rect 25504 33940 25556 33992
rect 30472 33983 30524 33992
rect 30472 33949 30481 33983
rect 30481 33949 30515 33983
rect 30515 33949 30524 33983
rect 30472 33940 30524 33949
rect 30840 33983 30892 33992
rect 30840 33949 30849 33983
rect 30849 33949 30883 33983
rect 30883 33949 30892 33983
rect 30840 33940 30892 33949
rect 25872 33872 25924 33924
rect 27436 33872 27488 33924
rect 29644 33872 29696 33924
rect 30380 33872 30432 33924
rect 16764 33804 16816 33856
rect 17316 33804 17368 33856
rect 22284 33804 22336 33856
rect 25964 33847 26016 33856
rect 25964 33813 25973 33847
rect 25973 33813 26007 33847
rect 26007 33813 26016 33847
rect 25964 33804 26016 33813
rect 27896 33804 27948 33856
rect 29736 33804 29788 33856
rect 47216 33915 47268 33924
rect 47216 33881 47225 33915
rect 47225 33881 47259 33915
rect 47259 33881 47268 33915
rect 47216 33872 47268 33881
rect 31300 33804 31352 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 17040 33600 17092 33652
rect 19248 33600 19300 33652
rect 16672 33507 16724 33516
rect 16672 33473 16681 33507
rect 16681 33473 16715 33507
rect 16715 33473 16724 33507
rect 16672 33464 16724 33473
rect 17224 33532 17276 33584
rect 17500 33464 17552 33516
rect 20904 33532 20956 33584
rect 24676 33532 24728 33584
rect 28448 33600 28500 33652
rect 29092 33600 29144 33652
rect 47768 33600 47820 33652
rect 19524 33507 19576 33516
rect 19524 33473 19533 33507
rect 19533 33473 19567 33507
rect 19567 33473 19576 33507
rect 19524 33464 19576 33473
rect 20720 33464 20772 33516
rect 21272 33464 21324 33516
rect 22744 33507 22796 33516
rect 22744 33473 22753 33507
rect 22753 33473 22787 33507
rect 22787 33473 22796 33507
rect 22744 33464 22796 33473
rect 24860 33464 24912 33516
rect 28908 33532 28960 33584
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 1860 33396 1912 33448
rect 17040 33396 17092 33448
rect 17316 33396 17368 33448
rect 28632 33507 28684 33516
rect 28632 33473 28641 33507
rect 28641 33473 28675 33507
rect 28675 33473 28684 33507
rect 28632 33464 28684 33473
rect 30472 33464 30524 33516
rect 31024 33464 31076 33516
rect 46848 33507 46900 33516
rect 46848 33473 46857 33507
rect 46857 33473 46891 33507
rect 46891 33473 46900 33507
rect 46848 33464 46900 33473
rect 47768 33464 47820 33516
rect 30840 33439 30892 33448
rect 30840 33405 30849 33439
rect 30849 33405 30883 33439
rect 30883 33405 30892 33439
rect 30840 33396 30892 33405
rect 19340 33328 19392 33380
rect 23572 33328 23624 33380
rect 23664 33328 23716 33380
rect 27620 33328 27672 33380
rect 31576 33328 31628 33380
rect 17224 33260 17276 33312
rect 20720 33260 20772 33312
rect 21364 33260 21416 33312
rect 22376 33260 22428 33312
rect 23112 33260 23164 33312
rect 23848 33260 23900 33312
rect 24952 33260 25004 33312
rect 27344 33260 27396 33312
rect 28540 33260 28592 33312
rect 28724 33260 28776 33312
rect 41420 33260 41472 33312
rect 47860 33303 47912 33312
rect 47860 33269 47869 33303
rect 47869 33269 47903 33303
rect 47903 33269 47912 33303
rect 47860 33260 47912 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1952 33099 2004 33108
rect 1952 33065 1961 33099
rect 1961 33065 1995 33099
rect 1995 33065 2004 33099
rect 1952 33056 2004 33065
rect 16672 33056 16724 33108
rect 17500 33056 17552 33108
rect 17776 33056 17828 33108
rect 22192 33056 22244 33108
rect 24860 33056 24912 33108
rect 25688 33056 25740 33108
rect 26148 33056 26200 33108
rect 27528 33056 27580 33108
rect 29644 33099 29696 33108
rect 1860 32895 1912 32904
rect 1860 32861 1869 32895
rect 1869 32861 1903 32895
rect 1903 32861 1912 32895
rect 1860 32852 1912 32861
rect 17040 32920 17092 32972
rect 18420 32920 18472 32972
rect 17224 32895 17276 32904
rect 17224 32861 17233 32895
rect 17233 32861 17267 32895
rect 17267 32861 17276 32895
rect 17224 32852 17276 32861
rect 19248 32852 19300 32904
rect 18604 32784 18656 32836
rect 19984 32852 20036 32904
rect 22376 32920 22428 32972
rect 24492 32852 24544 32904
rect 26332 32920 26384 32972
rect 27620 32920 27672 32972
rect 21272 32784 21324 32836
rect 27344 32852 27396 32904
rect 28540 32920 28592 32972
rect 29644 33065 29653 33099
rect 29653 33065 29687 33099
rect 29687 33065 29696 33099
rect 29644 33056 29696 33065
rect 28816 32988 28868 33040
rect 31116 32963 31168 32972
rect 31116 32929 31125 32963
rect 31125 32929 31159 32963
rect 31159 32929 31168 32963
rect 31116 32920 31168 32929
rect 47032 32920 47084 32972
rect 29552 32895 29604 32904
rect 26240 32784 26292 32836
rect 28264 32784 28316 32836
rect 29552 32861 29561 32895
rect 29561 32861 29595 32895
rect 29595 32861 29604 32895
rect 29552 32852 29604 32861
rect 46296 32895 46348 32904
rect 46296 32861 46305 32895
rect 46305 32861 46339 32895
rect 46339 32861 46348 32895
rect 46296 32852 46348 32861
rect 30564 32784 30616 32836
rect 31392 32827 31444 32836
rect 31392 32793 31401 32827
rect 31401 32793 31435 32827
rect 31435 32793 31444 32827
rect 31392 32784 31444 32793
rect 33692 32784 33744 32836
rect 46940 32784 46992 32836
rect 48136 32827 48188 32836
rect 48136 32793 48145 32827
rect 48145 32793 48179 32827
rect 48179 32793 48188 32827
rect 48136 32784 48188 32793
rect 2320 32716 2372 32768
rect 18236 32716 18288 32768
rect 19340 32716 19392 32768
rect 20812 32716 20864 32768
rect 25412 32759 25464 32768
rect 25412 32725 25421 32759
rect 25421 32725 25455 32759
rect 25455 32725 25464 32759
rect 25412 32716 25464 32725
rect 28448 32716 28500 32768
rect 29552 32716 29604 32768
rect 30656 32716 30708 32768
rect 31024 32716 31076 32768
rect 31668 32716 31720 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 21272 32555 21324 32564
rect 21272 32521 21281 32555
rect 21281 32521 21315 32555
rect 21315 32521 21324 32555
rect 21272 32512 21324 32521
rect 22744 32512 22796 32564
rect 23112 32512 23164 32564
rect 2320 32487 2372 32496
rect 2320 32453 2329 32487
rect 2329 32453 2363 32487
rect 2363 32453 2372 32487
rect 2320 32444 2372 32453
rect 23848 32487 23900 32496
rect 2136 32419 2188 32428
rect 2136 32385 2145 32419
rect 2145 32385 2179 32419
rect 2179 32385 2188 32419
rect 2136 32376 2188 32385
rect 16672 32376 16724 32428
rect 17776 32419 17828 32428
rect 4620 32308 4672 32360
rect 17224 32308 17276 32360
rect 17776 32385 17785 32419
rect 17785 32385 17819 32419
rect 17819 32385 17828 32419
rect 17776 32376 17828 32385
rect 18972 32376 19024 32428
rect 19340 32419 19392 32428
rect 19340 32385 19349 32419
rect 19349 32385 19383 32419
rect 19383 32385 19392 32419
rect 19340 32376 19392 32385
rect 19984 32376 20036 32428
rect 23848 32453 23857 32487
rect 23857 32453 23891 32487
rect 23891 32453 23900 32487
rect 23848 32444 23900 32453
rect 18052 32351 18104 32360
rect 18052 32317 18061 32351
rect 18061 32317 18095 32351
rect 18095 32317 18104 32351
rect 18052 32308 18104 32317
rect 19248 32308 19300 32360
rect 21180 32308 21232 32360
rect 22560 32376 22612 32428
rect 22928 32419 22980 32428
rect 22928 32385 22937 32419
rect 22937 32385 22971 32419
rect 22971 32385 22980 32419
rect 22928 32376 22980 32385
rect 23572 32419 23624 32428
rect 23572 32385 23581 32419
rect 23581 32385 23615 32419
rect 23615 32385 23624 32419
rect 23572 32376 23624 32385
rect 24952 32376 25004 32428
rect 25596 32444 25648 32496
rect 28632 32512 28684 32564
rect 31392 32512 31444 32564
rect 33692 32555 33744 32564
rect 33692 32521 33701 32555
rect 33701 32521 33735 32555
rect 33735 32521 33744 32555
rect 33692 32512 33744 32521
rect 46940 32555 46992 32564
rect 46940 32521 46949 32555
rect 46949 32521 46983 32555
rect 46983 32521 46992 32555
rect 46940 32512 46992 32521
rect 47032 32512 47084 32564
rect 25872 32444 25924 32496
rect 26240 32444 26292 32496
rect 41420 32444 41472 32496
rect 17684 32240 17736 32292
rect 1400 32172 1452 32224
rect 17224 32215 17276 32224
rect 17224 32181 17233 32215
rect 17233 32181 17267 32215
rect 17267 32181 17276 32215
rect 17224 32172 17276 32181
rect 17316 32172 17368 32224
rect 18696 32172 18748 32224
rect 20720 32240 20772 32292
rect 19340 32172 19392 32224
rect 21364 32172 21416 32224
rect 24584 32308 24636 32360
rect 25964 32308 26016 32360
rect 28172 32419 28224 32428
rect 28172 32385 28181 32419
rect 28181 32385 28215 32419
rect 28215 32385 28224 32419
rect 28172 32376 28224 32385
rect 28448 32376 28500 32428
rect 28540 32376 28592 32428
rect 29000 32419 29052 32428
rect 29000 32385 29009 32419
rect 29009 32385 29043 32419
rect 29043 32385 29052 32419
rect 29000 32376 29052 32385
rect 31300 32419 31352 32428
rect 24860 32240 24912 32292
rect 22376 32215 22428 32224
rect 22376 32181 22385 32215
rect 22385 32181 22419 32215
rect 22419 32181 22428 32215
rect 22376 32172 22428 32181
rect 22468 32172 22520 32224
rect 23940 32172 23992 32224
rect 25136 32172 25188 32224
rect 25320 32172 25372 32224
rect 30840 32308 30892 32360
rect 31300 32385 31309 32419
rect 31309 32385 31343 32419
rect 31343 32385 31352 32419
rect 31300 32376 31352 32385
rect 31484 32419 31536 32428
rect 31484 32385 31493 32419
rect 31493 32385 31527 32419
rect 31527 32385 31536 32419
rect 31484 32376 31536 32385
rect 31576 32419 31628 32428
rect 31576 32385 31585 32419
rect 31585 32385 31619 32419
rect 31619 32385 31628 32419
rect 31576 32376 31628 32385
rect 31760 32376 31812 32428
rect 31024 32308 31076 32360
rect 32680 32308 32732 32360
rect 33692 32376 33744 32428
rect 46204 32376 46256 32428
rect 47952 32419 48004 32428
rect 47952 32385 47961 32419
rect 47961 32385 47995 32419
rect 47995 32385 48004 32419
rect 47952 32376 48004 32385
rect 34152 32308 34204 32360
rect 26884 32240 26936 32292
rect 30472 32240 30524 32292
rect 31300 32240 31352 32292
rect 28080 32172 28132 32224
rect 28264 32172 28316 32224
rect 30196 32215 30248 32224
rect 30196 32181 30205 32215
rect 30205 32181 30239 32215
rect 30239 32181 30248 32215
rect 30196 32172 30248 32181
rect 30564 32172 30616 32224
rect 47400 32308 47452 32360
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 3240 31807 3292 31816
rect 3240 31773 3249 31807
rect 3249 31773 3283 31807
rect 3283 31773 3292 31807
rect 3240 31764 3292 31773
rect 3792 31807 3844 31816
rect 3792 31773 3801 31807
rect 3801 31773 3835 31807
rect 3835 31773 3844 31807
rect 3792 31764 3844 31773
rect 3976 31764 4028 31816
rect 17316 31968 17368 32020
rect 17776 31900 17828 31952
rect 18052 31900 18104 31952
rect 18696 31968 18748 32020
rect 21180 31943 21232 31952
rect 21180 31909 21189 31943
rect 21189 31909 21223 31943
rect 21223 31909 21232 31943
rect 21180 31900 21232 31909
rect 22928 31968 22980 32020
rect 28172 31968 28224 32020
rect 28908 31968 28960 32020
rect 29368 31968 29420 32020
rect 30196 31968 30248 32020
rect 30472 31968 30524 32020
rect 39856 31968 39908 32020
rect 46296 31968 46348 32020
rect 26884 31900 26936 31952
rect 16856 31832 16908 31884
rect 17684 31832 17736 31884
rect 7564 31671 7616 31680
rect 7564 31637 7573 31671
rect 7573 31637 7607 31671
rect 7607 31637 7616 31671
rect 7564 31628 7616 31637
rect 17868 31696 17920 31748
rect 17132 31628 17184 31680
rect 18328 31875 18380 31884
rect 18328 31841 18337 31875
rect 18337 31841 18371 31875
rect 18371 31841 18380 31875
rect 18328 31832 18380 31841
rect 18696 31832 18748 31884
rect 22468 31875 22520 31884
rect 22468 31841 22477 31875
rect 22477 31841 22511 31875
rect 22511 31841 22520 31875
rect 22468 31832 22520 31841
rect 22560 31832 22612 31884
rect 18604 31764 18656 31816
rect 18604 31628 18656 31680
rect 18972 31764 19024 31816
rect 20812 31764 20864 31816
rect 22008 31764 22060 31816
rect 22100 31764 22152 31816
rect 19432 31696 19484 31748
rect 22376 31807 22428 31816
rect 22376 31773 22385 31807
rect 22385 31773 22419 31807
rect 22419 31773 22428 31807
rect 22376 31764 22428 31773
rect 22744 31764 22796 31816
rect 23940 31832 23992 31884
rect 25872 31832 25924 31884
rect 27436 31832 27488 31884
rect 28080 31832 28132 31884
rect 30012 31900 30064 31952
rect 30748 31943 30800 31952
rect 30748 31909 30757 31943
rect 30757 31909 30791 31943
rect 30791 31909 30800 31943
rect 30748 31900 30800 31909
rect 34152 31943 34204 31952
rect 28724 31832 28776 31884
rect 23848 31807 23900 31816
rect 23848 31773 23857 31807
rect 23857 31773 23891 31807
rect 23891 31773 23900 31807
rect 23848 31764 23900 31773
rect 25044 31764 25096 31816
rect 29368 31764 29420 31816
rect 29552 31807 29604 31816
rect 29552 31773 29561 31807
rect 29561 31773 29595 31807
rect 29595 31773 29604 31807
rect 29552 31764 29604 31773
rect 31024 31832 31076 31884
rect 31116 31832 31168 31884
rect 34152 31909 34161 31943
rect 34161 31909 34195 31943
rect 34195 31909 34204 31943
rect 34152 31900 34204 31909
rect 33140 31832 33192 31884
rect 27712 31696 27764 31748
rect 30472 31807 30524 31816
rect 30472 31773 30481 31807
rect 30481 31773 30515 31807
rect 30515 31773 30524 31807
rect 31300 31807 31352 31816
rect 30472 31764 30524 31773
rect 31300 31773 31309 31807
rect 31309 31773 31343 31807
rect 31343 31773 31352 31807
rect 31300 31764 31352 31773
rect 31576 31764 31628 31816
rect 21272 31628 21324 31680
rect 22100 31628 22152 31680
rect 25228 31628 25280 31680
rect 29736 31628 29788 31680
rect 30748 31628 30800 31680
rect 33784 31764 33836 31816
rect 32404 31628 32456 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 17132 31424 17184 31476
rect 17868 31467 17920 31476
rect 17868 31433 17877 31467
rect 17877 31433 17911 31467
rect 17911 31433 17920 31467
rect 17868 31424 17920 31433
rect 19432 31424 19484 31476
rect 21456 31424 21508 31476
rect 23848 31424 23900 31476
rect 24400 31424 24452 31476
rect 27160 31424 27212 31476
rect 1860 31356 1912 31408
rect 18880 31356 18932 31408
rect 2596 31263 2648 31272
rect 2596 31229 2605 31263
rect 2605 31229 2639 31263
rect 2639 31229 2648 31263
rect 2596 31220 2648 31229
rect 4620 31220 4672 31272
rect 6552 31084 6604 31136
rect 16580 31288 16632 31340
rect 16764 31331 16816 31340
rect 16764 31297 16801 31331
rect 16801 31297 16816 31331
rect 16764 31288 16816 31297
rect 17132 31331 17184 31340
rect 19340 31356 19392 31408
rect 22376 31356 22428 31408
rect 22560 31356 22612 31408
rect 27344 31356 27396 31408
rect 27712 31424 27764 31476
rect 28908 31467 28960 31476
rect 28908 31433 28917 31467
rect 28917 31433 28951 31467
rect 28951 31433 28960 31467
rect 28908 31424 28960 31433
rect 33140 31467 33192 31476
rect 33140 31433 33149 31467
rect 33149 31433 33183 31467
rect 33183 31433 33192 31467
rect 33140 31424 33192 31433
rect 33784 31467 33836 31476
rect 33784 31433 33793 31467
rect 33793 31433 33827 31467
rect 33827 31433 33836 31467
rect 33784 31424 33836 31433
rect 46480 31424 46532 31476
rect 46848 31424 46900 31476
rect 17132 31297 17146 31331
rect 17146 31297 17180 31331
rect 17180 31297 17184 31331
rect 17132 31288 17184 31297
rect 17224 31084 17276 31136
rect 19432 31288 19484 31340
rect 20536 31288 20588 31340
rect 24584 31288 24636 31340
rect 25504 31331 25556 31340
rect 25504 31297 25513 31331
rect 25513 31297 25547 31331
rect 25547 31297 25556 31331
rect 25504 31288 25556 31297
rect 31208 31356 31260 31408
rect 19248 31263 19300 31272
rect 19248 31229 19257 31263
rect 19257 31229 19291 31263
rect 19291 31229 19300 31263
rect 19248 31220 19300 31229
rect 19984 31220 20036 31272
rect 20904 31152 20956 31204
rect 20996 31084 21048 31136
rect 22192 31220 22244 31272
rect 24860 31220 24912 31272
rect 25412 31220 25464 31272
rect 27620 31288 27672 31340
rect 28632 31288 28684 31340
rect 28816 31331 28868 31340
rect 28816 31297 28825 31331
rect 28825 31297 28859 31331
rect 28859 31297 28868 31331
rect 28816 31288 28868 31297
rect 29000 31331 29052 31340
rect 29000 31297 29009 31331
rect 29009 31297 29043 31331
rect 29043 31297 29052 31331
rect 29000 31288 29052 31297
rect 30840 31288 30892 31340
rect 32404 31331 32456 31340
rect 32404 31297 32413 31331
rect 32413 31297 32447 31331
rect 32447 31297 32456 31331
rect 32404 31288 32456 31297
rect 32588 31331 32640 31340
rect 32588 31297 32597 31331
rect 32597 31297 32631 31331
rect 32631 31297 32640 31331
rect 32588 31288 32640 31297
rect 32680 31331 32732 31340
rect 32680 31297 32689 31331
rect 32689 31297 32723 31331
rect 32723 31297 32732 31331
rect 32956 31331 33008 31340
rect 32680 31288 32732 31297
rect 32956 31297 32965 31331
rect 32965 31297 32999 31331
rect 32999 31297 33008 31331
rect 32956 31288 33008 31297
rect 33692 31331 33744 31340
rect 33692 31297 33701 31331
rect 33701 31297 33735 31331
rect 33735 31297 33744 31331
rect 33692 31288 33744 31297
rect 28264 31220 28316 31272
rect 30472 31220 30524 31272
rect 31116 31220 31168 31272
rect 32496 31220 32548 31272
rect 22100 31084 22152 31136
rect 25872 31084 25924 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 16580 30880 16632 30932
rect 20904 30880 20956 30932
rect 22192 30880 22244 30932
rect 22560 30880 22612 30932
rect 21640 30812 21692 30864
rect 22008 30812 22060 30864
rect 6552 30787 6604 30796
rect 6552 30753 6561 30787
rect 6561 30753 6595 30787
rect 6595 30753 6604 30787
rect 6552 30744 6604 30753
rect 7564 30744 7616 30796
rect 8208 30787 8260 30796
rect 8208 30753 8217 30787
rect 8217 30753 8251 30787
rect 8251 30753 8260 30787
rect 8208 30744 8260 30753
rect 20996 30744 21048 30796
rect 24676 30880 24728 30932
rect 25504 30923 25556 30932
rect 25504 30889 25513 30923
rect 25513 30889 25547 30923
rect 25547 30889 25556 30923
rect 25504 30880 25556 30889
rect 30196 30923 30248 30932
rect 30196 30889 30205 30923
rect 30205 30889 30239 30923
rect 30239 30889 30248 30923
rect 30196 30880 30248 30889
rect 30840 30880 30892 30932
rect 26332 30812 26384 30864
rect 26976 30855 27028 30864
rect 26976 30821 26985 30855
rect 26985 30821 27019 30855
rect 27019 30821 27028 30855
rect 26976 30812 27028 30821
rect 21272 30719 21324 30728
rect 21272 30685 21281 30719
rect 21281 30685 21315 30719
rect 21315 30685 21324 30719
rect 21272 30676 21324 30685
rect 21456 30719 21508 30728
rect 21456 30685 21463 30719
rect 21463 30685 21508 30719
rect 21456 30676 21508 30685
rect 21732 30719 21784 30728
rect 21732 30685 21746 30719
rect 21746 30685 21780 30719
rect 21780 30685 21784 30719
rect 21732 30676 21784 30685
rect 22560 30676 22612 30728
rect 18880 30608 18932 30660
rect 25228 30676 25280 30728
rect 30288 30744 30340 30796
rect 25320 30651 25372 30660
rect 25320 30617 25345 30651
rect 25345 30617 25372 30651
rect 28540 30676 28592 30728
rect 29000 30676 29052 30728
rect 30656 30719 30708 30728
rect 30656 30685 30665 30719
rect 30665 30685 30699 30719
rect 30699 30685 30708 30719
rect 30656 30676 30708 30685
rect 32404 30719 32456 30728
rect 32404 30685 32413 30719
rect 32413 30685 32447 30719
rect 32447 30685 32456 30719
rect 32404 30676 32456 30685
rect 32588 30812 32640 30864
rect 40408 30744 40460 30796
rect 47032 30744 47084 30796
rect 47676 30744 47728 30796
rect 32680 30719 32732 30728
rect 32680 30685 32689 30719
rect 32689 30685 32723 30719
rect 32723 30685 32732 30719
rect 32956 30719 33008 30728
rect 32680 30676 32732 30685
rect 32956 30685 32965 30719
rect 32965 30685 32999 30719
rect 32999 30685 33008 30719
rect 32956 30676 33008 30685
rect 25320 30608 25372 30617
rect 26516 30608 26568 30660
rect 26792 30651 26844 30660
rect 26792 30617 26801 30651
rect 26801 30617 26835 30651
rect 26835 30617 26844 30651
rect 26792 30608 26844 30617
rect 30288 30608 30340 30660
rect 46020 30608 46072 30660
rect 47768 30608 47820 30660
rect 25596 30540 25648 30592
rect 25964 30540 26016 30592
rect 28264 30540 28316 30592
rect 30380 30540 30432 30592
rect 33140 30583 33192 30592
rect 33140 30549 33149 30583
rect 33149 30549 33183 30583
rect 33183 30549 33192 30583
rect 33140 30540 33192 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 19432 30336 19484 30388
rect 20168 30336 20220 30388
rect 17960 30268 18012 30320
rect 16856 30200 16908 30252
rect 19064 30200 19116 30252
rect 19432 30243 19484 30252
rect 19432 30209 19441 30243
rect 19441 30209 19475 30243
rect 19475 30209 19484 30243
rect 19432 30200 19484 30209
rect 19524 30175 19576 30184
rect 19524 30141 19533 30175
rect 19533 30141 19567 30175
rect 19567 30141 19576 30175
rect 19524 30132 19576 30141
rect 19800 30243 19852 30252
rect 19800 30209 19809 30243
rect 19809 30209 19843 30243
rect 19843 30209 19852 30243
rect 19800 30200 19852 30209
rect 20076 30132 20128 30184
rect 28448 30336 28500 30388
rect 28816 30336 28868 30388
rect 24860 30243 24912 30252
rect 24860 30209 24869 30243
rect 24869 30209 24903 30243
rect 24903 30209 24912 30243
rect 24860 30200 24912 30209
rect 25320 30200 25372 30252
rect 25504 30200 25556 30252
rect 25964 30243 26016 30252
rect 25964 30209 25973 30243
rect 25973 30209 26007 30243
rect 26007 30209 26016 30243
rect 25964 30200 26016 30209
rect 27804 30200 27856 30252
rect 28908 30268 28960 30320
rect 29736 30336 29788 30388
rect 47768 30336 47820 30388
rect 48228 30336 48280 30388
rect 33140 30311 33192 30320
rect 33140 30277 33149 30311
rect 33149 30277 33183 30311
rect 33183 30277 33192 30311
rect 33140 30268 33192 30277
rect 33784 30268 33836 30320
rect 29000 30200 29052 30252
rect 29460 30243 29512 30252
rect 29460 30209 29469 30243
rect 29469 30209 29503 30243
rect 29503 30209 29512 30243
rect 29460 30200 29512 30209
rect 29644 30200 29696 30252
rect 29920 30200 29972 30252
rect 30840 30200 30892 30252
rect 25412 30132 25464 30184
rect 26792 30132 26844 30184
rect 30012 30132 30064 30184
rect 30288 30175 30340 30184
rect 30288 30141 30297 30175
rect 30297 30141 30331 30175
rect 30331 30141 30340 30175
rect 30288 30132 30340 30141
rect 31300 30175 31352 30184
rect 31300 30141 31309 30175
rect 31309 30141 31343 30175
rect 31343 30141 31352 30175
rect 31300 30132 31352 30141
rect 32864 30175 32916 30184
rect 32864 30141 32873 30175
rect 32873 30141 32907 30175
rect 32907 30141 32916 30175
rect 32864 30132 32916 30141
rect 29092 30064 29144 30116
rect 32404 30064 32456 30116
rect 19800 29996 19852 30048
rect 25320 29996 25372 30048
rect 25780 29996 25832 30048
rect 27436 29996 27488 30048
rect 27712 29996 27764 30048
rect 30656 29996 30708 30048
rect 31392 30039 31444 30048
rect 31392 30005 31401 30039
rect 31401 30005 31435 30039
rect 31435 30005 31444 30039
rect 31392 29996 31444 30005
rect 31760 29996 31812 30048
rect 32680 29996 32732 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 17960 29792 18012 29844
rect 19524 29792 19576 29844
rect 19984 29792 20036 29844
rect 22652 29792 22704 29844
rect 29000 29792 29052 29844
rect 29920 29835 29972 29844
rect 29920 29801 29929 29835
rect 29929 29801 29963 29835
rect 29963 29801 29972 29835
rect 29920 29792 29972 29801
rect 30196 29792 30248 29844
rect 31300 29792 31352 29844
rect 33784 29835 33836 29844
rect 33784 29801 33793 29835
rect 33793 29801 33827 29835
rect 33827 29801 33836 29835
rect 33784 29792 33836 29801
rect 19524 29699 19576 29708
rect 19524 29665 19533 29699
rect 19533 29665 19567 29699
rect 19567 29665 19576 29699
rect 19524 29656 19576 29665
rect 20352 29656 20404 29708
rect 18144 29588 18196 29640
rect 19800 29588 19852 29640
rect 20076 29588 20128 29640
rect 20720 29631 20772 29640
rect 20720 29597 20729 29631
rect 20729 29597 20763 29631
rect 20763 29597 20772 29631
rect 20720 29588 20772 29597
rect 24584 29588 24636 29640
rect 24860 29656 24912 29708
rect 27436 29656 27488 29708
rect 32864 29656 32916 29708
rect 25596 29588 25648 29640
rect 27068 29631 27120 29640
rect 27068 29597 27077 29631
rect 27077 29597 27111 29631
rect 27111 29597 27120 29631
rect 27068 29588 27120 29597
rect 29736 29631 29788 29640
rect 29736 29597 29745 29631
rect 29745 29597 29779 29631
rect 29779 29597 29788 29631
rect 29736 29588 29788 29597
rect 30012 29631 30064 29640
rect 30012 29597 30021 29631
rect 30021 29597 30055 29631
rect 30055 29597 30064 29631
rect 33692 29631 33744 29640
rect 30012 29588 30064 29597
rect 33692 29597 33701 29631
rect 33701 29597 33735 29631
rect 33735 29597 33744 29631
rect 33692 29588 33744 29597
rect 48136 29631 48188 29640
rect 48136 29597 48145 29631
rect 48145 29597 48179 29631
rect 48179 29597 48188 29631
rect 48136 29588 48188 29597
rect 20812 29520 20864 29572
rect 27436 29520 27488 29572
rect 28356 29520 28408 29572
rect 32128 29520 32180 29572
rect 20536 29452 20588 29504
rect 23112 29452 23164 29504
rect 27988 29452 28040 29504
rect 30012 29452 30064 29504
rect 47952 29495 48004 29504
rect 47952 29461 47961 29495
rect 47961 29461 47995 29495
rect 47995 29461 48004 29495
rect 47952 29452 48004 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 19984 29248 20036 29300
rect 20904 29248 20956 29300
rect 21732 29248 21784 29300
rect 25412 29291 25464 29300
rect 16856 29180 16908 29232
rect 16672 29155 16724 29164
rect 16672 29121 16681 29155
rect 16681 29121 16715 29155
rect 16715 29121 16724 29155
rect 16672 29112 16724 29121
rect 18236 29112 18288 29164
rect 19892 29112 19944 29164
rect 20076 29112 20128 29164
rect 20536 29155 20588 29164
rect 20536 29121 20545 29155
rect 20545 29121 20579 29155
rect 20579 29121 20588 29155
rect 20536 29112 20588 29121
rect 21916 29180 21968 29232
rect 23020 29180 23072 29232
rect 19432 28976 19484 29028
rect 21824 29112 21876 29164
rect 21180 29044 21232 29096
rect 22100 29112 22152 29164
rect 24032 29112 24084 29164
rect 24584 29112 24636 29164
rect 22928 29087 22980 29096
rect 22928 29053 22937 29087
rect 22937 29053 22971 29087
rect 22971 29053 22980 29087
rect 22928 29044 22980 29053
rect 22652 28976 22704 29028
rect 25412 29257 25421 29291
rect 25421 29257 25455 29291
rect 25455 29257 25464 29291
rect 25412 29248 25464 29257
rect 27436 29291 27488 29300
rect 27436 29257 27445 29291
rect 27445 29257 27479 29291
rect 27479 29257 27488 29291
rect 27436 29248 27488 29257
rect 29736 29248 29788 29300
rect 32128 29248 32180 29300
rect 27712 29155 27764 29164
rect 27712 29121 27721 29155
rect 27721 29121 27755 29155
rect 27755 29121 27764 29155
rect 27988 29155 28040 29164
rect 27712 29112 27764 29121
rect 27988 29121 27997 29155
rect 27997 29121 28031 29155
rect 28031 29121 28040 29155
rect 27988 29112 28040 29121
rect 28816 29155 28868 29164
rect 28816 29121 28825 29155
rect 28825 29121 28859 29155
rect 28859 29121 28868 29155
rect 28816 29112 28868 29121
rect 30288 29112 30340 29164
rect 43352 29180 43404 29232
rect 25136 29087 25188 29096
rect 25136 29053 25145 29087
rect 25145 29053 25179 29087
rect 25179 29053 25188 29087
rect 25136 29044 25188 29053
rect 25688 29044 25740 29096
rect 27804 28976 27856 29028
rect 27988 28976 28040 29028
rect 29000 29044 29052 29096
rect 30564 29112 30616 29164
rect 30748 29155 30800 29164
rect 30748 29121 30757 29155
rect 30757 29121 30791 29155
rect 30791 29121 30800 29155
rect 30748 29112 30800 29121
rect 29644 28976 29696 29028
rect 30012 28976 30064 29028
rect 30656 28976 30708 29028
rect 24400 28951 24452 28960
rect 24400 28917 24409 28951
rect 24409 28917 24443 28951
rect 24443 28917 24452 28951
rect 24400 28908 24452 28917
rect 25504 28908 25556 28960
rect 28264 28908 28316 28960
rect 33692 29112 33744 29164
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 20076 28704 20128 28756
rect 22928 28704 22980 28756
rect 26976 28704 27028 28756
rect 27160 28704 27212 28756
rect 28356 28747 28408 28756
rect 28356 28713 28365 28747
rect 28365 28713 28399 28747
rect 28399 28713 28408 28747
rect 28356 28704 28408 28713
rect 30748 28704 30800 28756
rect 20720 28636 20772 28688
rect 30196 28636 30248 28688
rect 7472 28568 7524 28620
rect 19892 28611 19944 28620
rect 18144 28500 18196 28552
rect 18328 28475 18380 28484
rect 18328 28441 18337 28475
rect 18337 28441 18371 28475
rect 18371 28441 18380 28475
rect 18328 28432 18380 28441
rect 18512 28475 18564 28484
rect 18512 28441 18521 28475
rect 18521 28441 18555 28475
rect 18555 28441 18564 28475
rect 18512 28432 18564 28441
rect 19892 28577 19901 28611
rect 19901 28577 19935 28611
rect 19935 28577 19944 28611
rect 19892 28568 19944 28577
rect 22284 28568 22336 28620
rect 23480 28568 23532 28620
rect 25504 28568 25556 28620
rect 28540 28568 28592 28620
rect 19340 28500 19392 28552
rect 21088 28500 21140 28552
rect 22192 28500 22244 28552
rect 22652 28500 22704 28552
rect 23112 28543 23164 28552
rect 23112 28509 23121 28543
rect 23121 28509 23155 28543
rect 23155 28509 23164 28543
rect 23112 28500 23164 28509
rect 25412 28500 25464 28552
rect 28264 28543 28316 28552
rect 24492 28432 24544 28484
rect 28264 28509 28273 28543
rect 28273 28509 28307 28543
rect 28307 28509 28316 28543
rect 28264 28500 28316 28509
rect 30380 28543 30432 28552
rect 30380 28509 30389 28543
rect 30389 28509 30423 28543
rect 30423 28509 30432 28543
rect 30380 28500 30432 28509
rect 17776 28407 17828 28416
rect 17776 28373 17785 28407
rect 17785 28373 17819 28407
rect 17819 28373 17828 28407
rect 17776 28364 17828 28373
rect 19432 28364 19484 28416
rect 19984 28364 20036 28416
rect 20720 28364 20772 28416
rect 21456 28364 21508 28416
rect 24584 28364 24636 28416
rect 29460 28432 29512 28484
rect 30288 28475 30340 28484
rect 30288 28441 30297 28475
rect 30297 28441 30331 28475
rect 30331 28441 30340 28475
rect 30288 28432 30340 28441
rect 29552 28364 29604 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 18512 28160 18564 28212
rect 19340 28160 19392 28212
rect 22192 28203 22244 28212
rect 17776 28092 17828 28144
rect 19432 28092 19484 28144
rect 16672 28024 16724 28076
rect 19524 28067 19576 28076
rect 19524 28033 19533 28067
rect 19533 28033 19567 28067
rect 19567 28033 19576 28067
rect 19524 28024 19576 28033
rect 22192 28169 22201 28203
rect 22201 28169 22235 28203
rect 22235 28169 22244 28203
rect 22192 28160 22244 28169
rect 25596 28160 25648 28212
rect 20720 28092 20772 28144
rect 21088 28092 21140 28144
rect 21272 28092 21324 28144
rect 22100 28092 22152 28144
rect 21732 28024 21784 28076
rect 23480 28092 23532 28144
rect 24400 28092 24452 28144
rect 29460 28092 29512 28144
rect 29552 28135 29604 28144
rect 29552 28101 29561 28135
rect 29561 28101 29595 28135
rect 29595 28101 29604 28135
rect 29552 28092 29604 28101
rect 30656 28092 30708 28144
rect 24676 28067 24728 28076
rect 20996 27956 21048 28008
rect 22928 27956 22980 28008
rect 24676 28033 24685 28067
rect 24685 28033 24719 28067
rect 24719 28033 24728 28067
rect 24676 28024 24728 28033
rect 26332 28024 26384 28076
rect 30012 28067 30064 28076
rect 30012 28033 30021 28067
rect 30021 28033 30055 28067
rect 30055 28033 30064 28067
rect 30012 28024 30064 28033
rect 30196 28067 30248 28076
rect 30196 28033 30205 28067
rect 30205 28033 30239 28067
rect 30239 28033 30248 28067
rect 30196 28024 30248 28033
rect 31484 28024 31536 28076
rect 24768 27999 24820 28008
rect 18328 27820 18380 27872
rect 19248 27820 19300 27872
rect 21272 27888 21324 27940
rect 22192 27888 22244 27940
rect 24768 27965 24777 27999
rect 24777 27965 24811 27999
rect 24811 27965 24820 27999
rect 24768 27956 24820 27965
rect 20812 27820 20864 27872
rect 21088 27820 21140 27872
rect 23020 27863 23072 27872
rect 23020 27829 23029 27863
rect 23029 27829 23063 27863
rect 23063 27829 23072 27863
rect 23020 27820 23072 27829
rect 23940 27863 23992 27872
rect 23940 27829 23949 27863
rect 23949 27829 23983 27863
rect 23983 27829 23992 27863
rect 23940 27820 23992 27829
rect 24952 27888 25004 27940
rect 25136 27888 25188 27940
rect 24860 27820 24912 27872
rect 30012 27863 30064 27872
rect 30012 27829 30021 27863
rect 30021 27829 30055 27863
rect 30055 27829 30064 27863
rect 30012 27820 30064 27829
rect 38752 27820 38804 27872
rect 46296 28024 46348 28076
rect 46940 27863 46992 27872
rect 46940 27829 46949 27863
rect 46949 27829 46983 27863
rect 46983 27829 46992 27863
rect 46940 27820 46992 27829
rect 47768 27863 47820 27872
rect 47768 27829 47777 27863
rect 47777 27829 47811 27863
rect 47811 27829 47820 27863
rect 47768 27820 47820 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3332 27616 3384 27668
rect 15108 27616 15160 27668
rect 19524 27616 19576 27668
rect 20352 27616 20404 27668
rect 20720 27616 20772 27668
rect 21456 27659 21508 27668
rect 21456 27625 21465 27659
rect 21465 27625 21499 27659
rect 21499 27625 21508 27659
rect 21456 27616 21508 27625
rect 24676 27616 24728 27668
rect 26516 27616 26568 27668
rect 30380 27616 30432 27668
rect 2228 27548 2280 27600
rect 15016 27480 15068 27532
rect 16120 27523 16172 27532
rect 12992 27412 13044 27464
rect 16120 27489 16129 27523
rect 16129 27489 16163 27523
rect 16163 27489 16172 27523
rect 16120 27480 16172 27489
rect 16856 27480 16908 27532
rect 17040 27523 17092 27532
rect 17040 27489 17049 27523
rect 17049 27489 17083 27523
rect 17083 27489 17092 27523
rect 17040 27480 17092 27489
rect 20720 27480 20772 27532
rect 19248 27455 19300 27464
rect 14464 27387 14516 27396
rect 14464 27353 14473 27387
rect 14473 27353 14507 27387
rect 14507 27353 14516 27387
rect 14464 27344 14516 27353
rect 13268 27276 13320 27328
rect 19248 27421 19257 27455
rect 19257 27421 19291 27455
rect 19291 27421 19300 27455
rect 19248 27412 19300 27421
rect 19340 27412 19392 27464
rect 20260 27455 20312 27464
rect 20260 27421 20269 27455
rect 20269 27421 20303 27455
rect 20303 27421 20312 27455
rect 20260 27412 20312 27421
rect 16764 27387 16816 27396
rect 16764 27353 16773 27387
rect 16773 27353 16807 27387
rect 16807 27353 16816 27387
rect 16764 27344 16816 27353
rect 16856 27344 16908 27396
rect 22284 27412 22336 27464
rect 20996 27387 21048 27396
rect 20996 27353 21005 27387
rect 21005 27353 21039 27387
rect 21039 27353 21048 27387
rect 20996 27344 21048 27353
rect 21088 27344 21140 27396
rect 23020 27412 23072 27464
rect 23940 27344 23992 27396
rect 24952 27412 25004 27464
rect 25596 27548 25648 27600
rect 25780 27548 25832 27600
rect 31116 27591 31168 27600
rect 31116 27557 31125 27591
rect 31125 27557 31159 27591
rect 31159 27557 31168 27591
rect 31116 27548 31168 27557
rect 31392 27548 31444 27600
rect 25596 27412 25648 27464
rect 26332 27412 26384 27464
rect 28908 27480 28960 27532
rect 26148 27344 26200 27396
rect 27896 27412 27948 27464
rect 31208 27480 31260 27532
rect 42432 27616 42484 27668
rect 45560 27616 45612 27668
rect 47768 27548 47820 27600
rect 30196 27455 30248 27464
rect 19340 27319 19392 27328
rect 19340 27285 19349 27319
rect 19349 27285 19383 27319
rect 19383 27285 19392 27319
rect 19340 27276 19392 27285
rect 21364 27276 21416 27328
rect 22928 27276 22980 27328
rect 24952 27276 25004 27328
rect 25504 27276 25556 27328
rect 25964 27276 26016 27328
rect 26884 27319 26936 27328
rect 26884 27285 26893 27319
rect 26893 27285 26927 27319
rect 26927 27285 26936 27319
rect 26884 27276 26936 27285
rect 26976 27276 27028 27328
rect 28264 27319 28316 27328
rect 28264 27285 28273 27319
rect 28273 27285 28307 27319
rect 28307 27285 28316 27319
rect 28264 27276 28316 27285
rect 30196 27421 30205 27455
rect 30205 27421 30239 27455
rect 30239 27421 30248 27455
rect 30196 27412 30248 27421
rect 31760 27455 31812 27464
rect 31760 27421 31769 27455
rect 31769 27421 31803 27455
rect 31803 27421 31812 27455
rect 31944 27455 31996 27464
rect 31760 27412 31812 27421
rect 31944 27421 31953 27455
rect 31953 27421 31987 27455
rect 31987 27421 31996 27455
rect 31944 27412 31996 27421
rect 46940 27480 46992 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 32312 27412 32364 27464
rect 31392 27276 31444 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 13268 27115 13320 27124
rect 13268 27081 13277 27115
rect 13277 27081 13311 27115
rect 13311 27081 13320 27115
rect 13268 27072 13320 27081
rect 14464 27072 14516 27124
rect 16764 27072 16816 27124
rect 19432 27115 19484 27124
rect 19432 27081 19441 27115
rect 19441 27081 19475 27115
rect 19475 27081 19484 27115
rect 19432 27072 19484 27081
rect 20260 27072 20312 27124
rect 12440 27004 12492 27056
rect 11244 26868 11296 26920
rect 11520 26911 11572 26920
rect 11520 26877 11529 26911
rect 11529 26877 11563 26911
rect 11563 26877 11572 26911
rect 11520 26868 11572 26877
rect 12348 26868 12400 26920
rect 17408 27004 17460 27056
rect 21456 27004 21508 27056
rect 22192 27047 22244 27056
rect 22192 27013 22201 27047
rect 22201 27013 22235 27047
rect 22235 27013 22244 27047
rect 22928 27072 22980 27124
rect 22192 27004 22244 27013
rect 24492 27004 24544 27056
rect 14280 26979 14332 26988
rect 14280 26945 14289 26979
rect 14289 26945 14323 26979
rect 14323 26945 14332 26979
rect 14280 26936 14332 26945
rect 17224 26936 17276 26988
rect 19340 26979 19392 26988
rect 19340 26945 19349 26979
rect 19349 26945 19383 26979
rect 19383 26945 19392 26979
rect 19340 26936 19392 26945
rect 19984 26936 20036 26988
rect 17960 26868 18012 26920
rect 20720 26936 20772 26988
rect 21272 26936 21324 26988
rect 21364 26936 21416 26988
rect 21916 26979 21968 26988
rect 21916 26945 21926 26979
rect 21926 26945 21960 26979
rect 21960 26945 21968 26979
rect 22100 26979 22152 26988
rect 21916 26936 21968 26945
rect 22100 26945 22109 26979
rect 22109 26945 22143 26979
rect 22143 26945 22152 26979
rect 22100 26936 22152 26945
rect 22560 26936 22612 26988
rect 24768 26936 24820 26988
rect 25136 27047 25188 27056
rect 25136 27013 25170 27047
rect 25170 27013 25188 27047
rect 25136 27004 25188 27013
rect 25780 27004 25832 27056
rect 26976 27072 27028 27124
rect 27620 27072 27672 27124
rect 30472 27072 30524 27124
rect 31484 27115 31536 27124
rect 31484 27081 31493 27115
rect 31493 27081 31527 27115
rect 31527 27081 31536 27115
rect 31484 27072 31536 27081
rect 24952 26911 25004 26920
rect 24952 26877 24961 26911
rect 24961 26877 24995 26911
rect 24995 26877 25004 26911
rect 24952 26868 25004 26877
rect 20996 26800 21048 26852
rect 25688 26868 25740 26920
rect 15200 26732 15252 26784
rect 19984 26732 20036 26784
rect 20812 26732 20864 26784
rect 22100 26732 22152 26784
rect 26516 26936 26568 26988
rect 27528 26979 27580 26988
rect 27528 26945 27537 26979
rect 27537 26945 27571 26979
rect 27571 26945 27580 26979
rect 27528 26936 27580 26945
rect 28264 26936 28316 26988
rect 30656 27047 30708 27056
rect 30656 27013 30665 27047
rect 30665 27013 30699 27047
rect 30699 27013 30708 27047
rect 30656 27004 30708 27013
rect 31208 27004 31260 27056
rect 30380 26979 30432 26988
rect 29736 26868 29788 26920
rect 26240 26800 26292 26852
rect 26332 26800 26384 26852
rect 30380 26945 30389 26979
rect 30389 26945 30423 26979
rect 30423 26945 30432 26979
rect 30380 26936 30432 26945
rect 30564 26979 30616 26988
rect 30564 26945 30573 26979
rect 30573 26945 30607 26979
rect 30607 26945 30616 26979
rect 30564 26936 30616 26945
rect 31392 26979 31444 26988
rect 30472 26868 30524 26920
rect 31392 26945 31401 26979
rect 31401 26945 31435 26979
rect 31435 26945 31444 26979
rect 31392 26936 31444 26945
rect 31576 26979 31628 26988
rect 31576 26945 31585 26979
rect 31585 26945 31619 26979
rect 31619 26945 31628 26979
rect 31576 26936 31628 26945
rect 32312 26979 32364 26988
rect 32312 26945 32321 26979
rect 32321 26945 32355 26979
rect 32355 26945 32364 26979
rect 32312 26936 32364 26945
rect 31944 26868 31996 26920
rect 46572 26868 46624 26920
rect 46756 26868 46808 26920
rect 25688 26732 25740 26784
rect 25780 26775 25832 26784
rect 25780 26741 25789 26775
rect 25789 26741 25823 26775
rect 25823 26741 25832 26775
rect 25780 26732 25832 26741
rect 25964 26732 26016 26784
rect 31300 26732 31352 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 11244 26571 11296 26580
rect 11244 26537 11253 26571
rect 11253 26537 11287 26571
rect 11287 26537 11296 26571
rect 11244 26528 11296 26537
rect 20352 26571 20404 26580
rect 20352 26537 20361 26571
rect 20361 26537 20395 26571
rect 20395 26537 20404 26571
rect 20352 26528 20404 26537
rect 21916 26528 21968 26580
rect 15108 26460 15160 26512
rect 12624 26392 12676 26444
rect 15200 26435 15252 26444
rect 15200 26401 15209 26435
rect 15209 26401 15243 26435
rect 15243 26401 15252 26435
rect 15200 26392 15252 26401
rect 21088 26460 21140 26512
rect 20260 26392 20312 26444
rect 12716 26324 12768 26376
rect 12992 26324 13044 26376
rect 14740 26324 14792 26376
rect 12532 26256 12584 26308
rect 20352 26324 20404 26376
rect 22192 26324 22244 26376
rect 25136 26528 25188 26580
rect 26884 26528 26936 26580
rect 28908 26571 28960 26580
rect 28908 26537 28917 26571
rect 28917 26537 28951 26571
rect 28951 26537 28960 26571
rect 28908 26528 28960 26537
rect 32312 26528 32364 26580
rect 24676 26460 24728 26512
rect 25688 26460 25740 26512
rect 29460 26460 29512 26512
rect 24952 26392 25004 26444
rect 24860 26367 24912 26376
rect 24860 26333 24869 26367
rect 24869 26333 24903 26367
rect 24903 26333 24912 26367
rect 24860 26324 24912 26333
rect 16488 26256 16540 26308
rect 24768 26256 24820 26308
rect 26976 26324 27028 26376
rect 27160 26367 27212 26376
rect 27160 26333 27169 26367
rect 27169 26333 27203 26367
rect 27203 26333 27212 26367
rect 27160 26324 27212 26333
rect 29736 26367 29788 26376
rect 25688 26299 25740 26308
rect 25688 26265 25697 26299
rect 25697 26265 25731 26299
rect 25731 26265 25740 26299
rect 25688 26256 25740 26265
rect 26148 26256 26200 26308
rect 29092 26256 29144 26308
rect 29736 26333 29745 26367
rect 29745 26333 29779 26367
rect 29779 26333 29788 26367
rect 29736 26324 29788 26333
rect 29920 26460 29972 26512
rect 30380 26392 30432 26444
rect 31300 26435 31352 26444
rect 31300 26401 31309 26435
rect 31309 26401 31343 26435
rect 31343 26401 31352 26435
rect 31300 26392 31352 26401
rect 45192 26324 45244 26376
rect 31576 26256 31628 26308
rect 31760 26256 31812 26308
rect 30104 26231 30156 26240
rect 30104 26197 30113 26231
rect 30113 26197 30147 26231
rect 30147 26197 30156 26231
rect 30104 26188 30156 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 11520 25984 11572 26036
rect 12440 25984 12492 26036
rect 16856 25984 16908 26036
rect 22192 25984 22244 26036
rect 24032 25984 24084 26036
rect 27528 26027 27580 26036
rect 27528 25993 27537 26027
rect 27537 25993 27571 26027
rect 27571 25993 27580 26027
rect 27528 25984 27580 25993
rect 29092 26027 29144 26036
rect 29092 25993 29101 26027
rect 29101 25993 29135 26027
rect 29135 25993 29144 26027
rect 29092 25984 29144 25993
rect 31760 25984 31812 26036
rect 10692 25891 10744 25900
rect 10692 25857 10701 25891
rect 10701 25857 10735 25891
rect 10735 25857 10744 25891
rect 10692 25848 10744 25857
rect 12440 25848 12492 25900
rect 14004 25848 14056 25900
rect 16764 25848 16816 25900
rect 13176 25780 13228 25832
rect 13452 25780 13504 25832
rect 11796 25712 11848 25764
rect 14740 25712 14792 25764
rect 22100 25959 22152 25968
rect 22100 25925 22109 25959
rect 22109 25925 22143 25959
rect 22143 25925 22152 25959
rect 22100 25916 22152 25925
rect 22836 25916 22888 25968
rect 18236 25848 18288 25900
rect 19984 25848 20036 25900
rect 21824 25891 21876 25900
rect 21824 25857 21833 25891
rect 21833 25857 21867 25891
rect 21867 25857 21876 25891
rect 21824 25848 21876 25857
rect 23388 25848 23440 25900
rect 25504 25848 25556 25900
rect 29460 25916 29512 25968
rect 30012 25959 30064 25968
rect 30012 25925 30021 25959
rect 30021 25925 30055 25959
rect 30055 25925 30064 25959
rect 30012 25916 30064 25925
rect 18144 25780 18196 25832
rect 28540 25780 28592 25832
rect 30104 25848 30156 25900
rect 46296 25891 46348 25900
rect 30288 25780 30340 25832
rect 46296 25857 46305 25891
rect 46305 25857 46339 25891
rect 46339 25857 46348 25891
rect 46296 25848 46348 25857
rect 12808 25644 12860 25696
rect 14464 25644 14516 25696
rect 15108 25687 15160 25696
rect 15108 25653 15117 25687
rect 15117 25653 15151 25687
rect 15151 25653 15160 25687
rect 15108 25644 15160 25653
rect 15936 25644 15988 25696
rect 18052 25644 18104 25696
rect 18420 25687 18472 25696
rect 18420 25653 18429 25687
rect 18429 25653 18463 25687
rect 18463 25653 18472 25687
rect 18420 25644 18472 25653
rect 25136 25644 25188 25696
rect 25412 25644 25464 25696
rect 29920 25644 29972 25696
rect 46480 25644 46532 25696
rect 47768 25687 47820 25696
rect 47768 25653 47777 25687
rect 47777 25653 47811 25687
rect 47811 25653 47820 25687
rect 47768 25644 47820 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 11796 25483 11848 25492
rect 11796 25449 11805 25483
rect 11805 25449 11839 25483
rect 11839 25449 11848 25483
rect 11796 25440 11848 25449
rect 16764 25483 16816 25492
rect 16764 25449 16773 25483
rect 16773 25449 16807 25483
rect 16807 25449 16816 25483
rect 16764 25440 16816 25449
rect 17960 25440 18012 25492
rect 18236 25483 18288 25492
rect 18236 25449 18245 25483
rect 18245 25449 18279 25483
rect 18279 25449 18288 25483
rect 18236 25440 18288 25449
rect 22836 25440 22888 25492
rect 25780 25440 25832 25492
rect 11612 25372 11664 25424
rect 12624 25372 12676 25424
rect 13360 25372 13412 25424
rect 16488 25372 16540 25424
rect 8300 25304 8352 25356
rect 14464 25347 14516 25356
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 2044 25100 2096 25152
rect 9128 25211 9180 25220
rect 9128 25177 9137 25211
rect 9137 25177 9171 25211
rect 9171 25177 9180 25211
rect 9128 25168 9180 25177
rect 11704 25236 11756 25288
rect 12348 25236 12400 25288
rect 12072 25168 12124 25220
rect 14464 25313 14473 25347
rect 14473 25313 14507 25347
rect 14507 25313 14516 25347
rect 14464 25304 14516 25313
rect 25688 25372 25740 25424
rect 14188 25279 14240 25288
rect 14188 25245 14197 25279
rect 14197 25245 14231 25279
rect 14231 25245 14240 25279
rect 14188 25236 14240 25245
rect 16488 25279 16540 25288
rect 16488 25245 16497 25279
rect 16497 25245 16531 25279
rect 16531 25245 16540 25279
rect 16488 25236 16540 25245
rect 13176 25168 13228 25220
rect 15108 25168 15160 25220
rect 11520 25143 11572 25152
rect 11520 25109 11529 25143
rect 11529 25109 11563 25143
rect 11563 25109 11572 25143
rect 11520 25100 11572 25109
rect 11612 25143 11664 25152
rect 11612 25109 11621 25143
rect 11621 25109 11655 25143
rect 11655 25109 11664 25143
rect 18512 25279 18564 25288
rect 11612 25100 11664 25109
rect 12716 25100 12768 25152
rect 13544 25100 13596 25152
rect 14004 25100 14056 25152
rect 16396 25100 16448 25152
rect 16488 25100 16540 25152
rect 17500 25143 17552 25152
rect 17500 25109 17509 25143
rect 17509 25109 17543 25143
rect 17543 25109 17552 25143
rect 18512 25245 18521 25279
rect 18521 25245 18555 25279
rect 18555 25245 18564 25279
rect 18512 25236 18564 25245
rect 27160 25304 27212 25356
rect 30380 25440 30432 25492
rect 31576 25440 31628 25492
rect 29920 25347 29972 25356
rect 29920 25313 29929 25347
rect 29929 25313 29963 25347
rect 29963 25313 29972 25347
rect 29920 25304 29972 25313
rect 46480 25347 46532 25356
rect 46480 25313 46489 25347
rect 46489 25313 46523 25347
rect 46523 25313 46532 25347
rect 46480 25304 46532 25313
rect 48136 25347 48188 25356
rect 48136 25313 48145 25347
rect 48145 25313 48179 25347
rect 48179 25313 48188 25347
rect 48136 25304 48188 25313
rect 23388 25236 23440 25288
rect 45836 25236 45888 25288
rect 19340 25168 19392 25220
rect 25136 25168 25188 25220
rect 30932 25168 30984 25220
rect 17500 25100 17552 25109
rect 17868 25100 17920 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9128 24896 9180 24948
rect 11520 24896 11572 24948
rect 12716 24896 12768 24948
rect 13544 24896 13596 24948
rect 8944 24760 8996 24812
rect 10692 24760 10744 24812
rect 11796 24828 11848 24880
rect 12808 24871 12860 24880
rect 12808 24837 12817 24871
rect 12817 24837 12851 24871
rect 12851 24837 12860 24871
rect 12808 24828 12860 24837
rect 14188 24896 14240 24948
rect 16764 24896 16816 24948
rect 19340 24896 19392 24948
rect 23388 24896 23440 24948
rect 26148 24939 26200 24948
rect 26148 24905 26157 24939
rect 26157 24905 26191 24939
rect 26191 24905 26200 24939
rect 26148 24896 26200 24905
rect 18420 24828 18472 24880
rect 25412 24828 25464 24880
rect 11612 24760 11664 24812
rect 12072 24760 12124 24812
rect 12532 24803 12584 24812
rect 12532 24769 12541 24803
rect 12541 24769 12575 24803
rect 12575 24769 12584 24803
rect 12532 24760 12584 24769
rect 14188 24760 14240 24812
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 15936 24803 15988 24812
rect 15936 24769 15945 24803
rect 15945 24769 15979 24803
rect 15979 24769 15988 24803
rect 15936 24760 15988 24769
rect 16396 24760 16448 24812
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 17040 24760 17092 24812
rect 18052 24803 18104 24812
rect 18052 24769 18061 24803
rect 18061 24769 18095 24803
rect 18095 24769 18104 24803
rect 18052 24760 18104 24769
rect 11704 24735 11756 24744
rect 11704 24701 11713 24735
rect 11713 24701 11747 24735
rect 11747 24701 11756 24735
rect 11704 24692 11756 24701
rect 13176 24692 13228 24744
rect 9680 24599 9732 24608
rect 9680 24565 9689 24599
rect 9689 24565 9723 24599
rect 9723 24565 9732 24599
rect 9680 24556 9732 24565
rect 10324 24599 10376 24608
rect 10324 24565 10333 24599
rect 10333 24565 10367 24599
rect 10367 24565 10376 24599
rect 10324 24556 10376 24565
rect 13360 24556 13412 24608
rect 19524 24624 19576 24676
rect 22928 24803 22980 24812
rect 20536 24692 20588 24744
rect 22928 24769 22937 24803
rect 22937 24769 22971 24803
rect 22971 24769 22980 24803
rect 22928 24760 22980 24769
rect 28264 24803 28316 24812
rect 28264 24769 28273 24803
rect 28273 24769 28307 24803
rect 28307 24769 28316 24803
rect 28264 24760 28316 24769
rect 30288 24760 30340 24812
rect 30932 24760 30984 24812
rect 38752 24803 38804 24812
rect 38752 24769 38761 24803
rect 38761 24769 38795 24803
rect 38795 24769 38804 24803
rect 38752 24760 38804 24769
rect 45192 24803 45244 24812
rect 45192 24769 45201 24803
rect 45201 24769 45235 24803
rect 45235 24769 45244 24803
rect 45192 24760 45244 24769
rect 46756 24760 46808 24812
rect 47584 24803 47636 24812
rect 47584 24769 47593 24803
rect 47593 24769 47627 24803
rect 47627 24769 47636 24803
rect 47584 24760 47636 24769
rect 21824 24692 21876 24744
rect 24676 24735 24728 24744
rect 24676 24701 24685 24735
rect 24685 24701 24719 24735
rect 24719 24701 24728 24735
rect 24676 24692 24728 24701
rect 25044 24692 25096 24744
rect 22100 24624 22152 24676
rect 26424 24624 26476 24676
rect 40592 24692 40644 24744
rect 40960 24735 41012 24744
rect 40960 24701 40969 24735
rect 40969 24701 41003 24735
rect 41003 24701 41012 24735
rect 45376 24735 45428 24744
rect 40960 24692 41012 24701
rect 45376 24701 45385 24735
rect 45385 24701 45419 24735
rect 45419 24701 45428 24735
rect 45376 24692 45428 24701
rect 46848 24735 46900 24744
rect 46848 24701 46857 24735
rect 46857 24701 46891 24735
rect 46891 24701 46900 24735
rect 46848 24692 46900 24701
rect 16028 24599 16080 24608
rect 16028 24565 16037 24599
rect 16037 24565 16071 24599
rect 16071 24565 16080 24599
rect 16028 24556 16080 24565
rect 17132 24556 17184 24608
rect 20444 24556 20496 24608
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 23020 24556 23072 24608
rect 27344 24556 27396 24608
rect 28356 24599 28408 24608
rect 28356 24565 28365 24599
rect 28365 24565 28399 24599
rect 28399 24565 28408 24599
rect 28356 24556 28408 24565
rect 45560 24624 45612 24676
rect 40960 24556 41012 24608
rect 46480 24556 46532 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 10784 24352 10836 24404
rect 13452 24395 13504 24404
rect 13452 24361 13461 24395
rect 13461 24361 13495 24395
rect 13495 24361 13504 24395
rect 13452 24352 13504 24361
rect 14188 24395 14240 24404
rect 14188 24361 14197 24395
rect 14197 24361 14231 24395
rect 14231 24361 14240 24395
rect 14188 24352 14240 24361
rect 9680 24284 9732 24336
rect 10324 24259 10376 24268
rect 10324 24225 10333 24259
rect 10333 24225 10367 24259
rect 10367 24225 10376 24259
rect 10324 24216 10376 24225
rect 11612 24284 11664 24336
rect 16028 24284 16080 24336
rect 12440 24148 12492 24200
rect 13728 24216 13780 24268
rect 13360 24191 13412 24200
rect 13360 24157 13369 24191
rect 13369 24157 13403 24191
rect 13403 24157 13412 24191
rect 13360 24148 13412 24157
rect 13544 24191 13596 24200
rect 13544 24157 13553 24191
rect 13553 24157 13587 24191
rect 13587 24157 13596 24191
rect 13544 24148 13596 24157
rect 16856 24216 16908 24268
rect 16672 24148 16724 24200
rect 17868 24148 17920 24200
rect 18512 24284 18564 24336
rect 20444 24259 20496 24268
rect 20444 24225 20453 24259
rect 20453 24225 20487 24259
rect 20487 24225 20496 24259
rect 20444 24216 20496 24225
rect 45652 24284 45704 24336
rect 27344 24259 27396 24268
rect 27344 24225 27353 24259
rect 27353 24225 27387 24259
rect 27387 24225 27396 24259
rect 27344 24216 27396 24225
rect 37280 24216 37332 24268
rect 47492 24352 47544 24404
rect 47768 24284 47820 24336
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 20260 24191 20312 24200
rect 20260 24157 20269 24191
rect 20269 24157 20303 24191
rect 20303 24157 20312 24191
rect 20260 24148 20312 24157
rect 22928 24148 22980 24200
rect 23388 24148 23440 24200
rect 27160 24191 27212 24200
rect 27160 24157 27169 24191
rect 27169 24157 27203 24191
rect 27203 24157 27212 24191
rect 27160 24148 27212 24157
rect 16396 24080 16448 24132
rect 17040 24080 17092 24132
rect 39212 24080 39264 24132
rect 46480 24259 46532 24268
rect 46480 24225 46489 24259
rect 46489 24225 46523 24259
rect 46523 24225 46532 24259
rect 46480 24216 46532 24225
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 42984 24148 43036 24200
rect 42800 24080 42852 24132
rect 45928 24148 45980 24200
rect 12072 24055 12124 24064
rect 12072 24021 12081 24055
rect 12081 24021 12115 24055
rect 12115 24021 12124 24055
rect 12072 24012 12124 24021
rect 16764 24055 16816 24064
rect 16764 24021 16773 24055
rect 16773 24021 16807 24055
rect 16807 24021 16816 24055
rect 16764 24012 16816 24021
rect 17868 24055 17920 24064
rect 17868 24021 17877 24055
rect 17877 24021 17911 24055
rect 17911 24021 17920 24055
rect 17868 24012 17920 24021
rect 19432 24012 19484 24064
rect 22744 24055 22796 24064
rect 22744 24021 22753 24055
rect 22753 24021 22787 24055
rect 22787 24021 22796 24055
rect 22744 24012 22796 24021
rect 24124 24012 24176 24064
rect 26056 24012 26108 24064
rect 41236 24012 41288 24064
rect 43168 24055 43220 24064
rect 43168 24021 43177 24055
rect 43177 24021 43211 24055
rect 43211 24021 43220 24055
rect 43168 24012 43220 24021
rect 47584 24012 47636 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 3608 23808 3660 23860
rect 25596 23808 25648 23860
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 12072 23740 12124 23792
rect 16672 23783 16724 23792
rect 16672 23749 16681 23783
rect 16681 23749 16715 23783
rect 16715 23749 16724 23783
rect 16672 23740 16724 23749
rect 14188 23672 14240 23724
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 8576 23647 8628 23656
rect 8576 23613 8585 23647
rect 8585 23613 8619 23647
rect 8619 23613 8628 23647
rect 8576 23604 8628 23613
rect 9772 23647 9824 23656
rect 9772 23613 9781 23647
rect 9781 23613 9815 23647
rect 9815 23613 9824 23647
rect 9772 23604 9824 23613
rect 16580 23604 16632 23656
rect 16764 23604 16816 23656
rect 17132 23715 17184 23724
rect 17132 23681 17141 23715
rect 17141 23681 17175 23715
rect 17175 23681 17184 23715
rect 17132 23672 17184 23681
rect 13728 23536 13780 23588
rect 17868 23740 17920 23792
rect 20168 23740 20220 23792
rect 20812 23740 20864 23792
rect 26056 23783 26108 23792
rect 19432 23672 19484 23724
rect 19892 23672 19944 23724
rect 26056 23749 26065 23783
rect 26065 23749 26099 23783
rect 26099 23749 26108 23783
rect 26056 23740 26108 23749
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 20260 23604 20312 23656
rect 22100 23604 22152 23656
rect 28264 23808 28316 23860
rect 40592 23851 40644 23860
rect 40592 23817 40601 23851
rect 40601 23817 40635 23851
rect 40635 23817 40644 23851
rect 40592 23808 40644 23817
rect 28356 23740 28408 23792
rect 37740 23715 37792 23724
rect 37740 23681 37749 23715
rect 37749 23681 37783 23715
rect 37783 23681 37792 23715
rect 37740 23672 37792 23681
rect 39212 23715 39264 23724
rect 39212 23681 39221 23715
rect 39221 23681 39255 23715
rect 39255 23681 39264 23715
rect 39212 23672 39264 23681
rect 41144 23715 41196 23724
rect 22376 23604 22428 23656
rect 20076 23468 20128 23520
rect 23112 23511 23164 23520
rect 23112 23477 23121 23511
rect 23121 23477 23155 23511
rect 23155 23477 23164 23511
rect 23112 23468 23164 23477
rect 25412 23511 25464 23520
rect 25412 23477 25421 23511
rect 25421 23477 25455 23511
rect 25455 23477 25464 23511
rect 25412 23468 25464 23477
rect 27804 23604 27856 23656
rect 25596 23536 25648 23588
rect 38476 23604 38528 23656
rect 41144 23681 41153 23715
rect 41153 23681 41187 23715
rect 41187 23681 41196 23715
rect 41144 23672 41196 23681
rect 41236 23672 41288 23724
rect 45376 23808 45428 23860
rect 47492 23740 47544 23792
rect 43352 23715 43404 23724
rect 43352 23681 43361 23715
rect 43361 23681 43395 23715
rect 43395 23681 43404 23715
rect 43352 23672 43404 23681
rect 44824 23672 44876 23724
rect 42524 23604 42576 23656
rect 45192 23647 45244 23656
rect 45192 23613 45201 23647
rect 45201 23613 45235 23647
rect 45235 23613 45244 23647
rect 45192 23604 45244 23613
rect 45652 23604 45704 23656
rect 46664 23647 46716 23656
rect 46664 23613 46673 23647
rect 46673 23613 46707 23647
rect 46707 23613 46716 23647
rect 46664 23604 46716 23613
rect 47400 23536 47452 23588
rect 38568 23468 38620 23520
rect 42984 23468 43036 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 8576 23264 8628 23316
rect 2136 23196 2188 23248
rect 39488 23264 39540 23316
rect 43168 23264 43220 23316
rect 43628 23264 43680 23316
rect 47032 23264 47084 23316
rect 47768 23264 47820 23316
rect 47952 23307 48004 23316
rect 47952 23273 47961 23307
rect 47961 23273 47995 23307
rect 47995 23273 48004 23307
rect 47952 23264 48004 23273
rect 13728 23128 13780 23180
rect 17132 23196 17184 23248
rect 18052 23196 18104 23248
rect 20076 23239 20128 23248
rect 20076 23205 20085 23239
rect 20085 23205 20119 23239
rect 20119 23205 20128 23239
rect 20076 23196 20128 23205
rect 20536 23196 20588 23248
rect 8944 23103 8996 23112
rect 8944 23069 8953 23103
rect 8953 23069 8987 23103
rect 8987 23069 8996 23103
rect 8944 23060 8996 23069
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 11704 23060 11756 23112
rect 14740 23103 14792 23112
rect 14740 23069 14749 23103
rect 14749 23069 14783 23103
rect 14783 23069 14792 23103
rect 14740 23060 14792 23069
rect 16764 23171 16816 23180
rect 16764 23137 16773 23171
rect 16773 23137 16807 23171
rect 16807 23137 16816 23171
rect 16764 23128 16816 23137
rect 16580 23060 16632 23112
rect 19892 23103 19944 23112
rect 19892 23069 19901 23103
rect 19901 23069 19935 23103
rect 19935 23069 19944 23103
rect 19892 23060 19944 23069
rect 22744 23128 22796 23180
rect 23204 23128 23256 23180
rect 25412 23171 25464 23180
rect 21732 23103 21784 23112
rect 17868 22992 17920 23044
rect 21732 23069 21741 23103
rect 21741 23069 21775 23103
rect 21775 23069 21784 23103
rect 21732 23060 21784 23069
rect 23112 23060 23164 23112
rect 11520 22924 11572 22976
rect 14372 22924 14424 22976
rect 15384 22924 15436 22976
rect 22100 22924 22152 22976
rect 22744 22924 22796 22976
rect 22836 22924 22888 22976
rect 23296 22924 23348 22976
rect 25412 23137 25421 23171
rect 25421 23137 25455 23171
rect 25455 23137 25464 23171
rect 25412 23128 25464 23137
rect 25964 23128 26016 23180
rect 26240 23128 26292 23180
rect 27896 23171 27948 23180
rect 27896 23137 27905 23171
rect 27905 23137 27939 23171
rect 27939 23137 27948 23171
rect 27896 23128 27948 23137
rect 28080 23128 28132 23180
rect 27804 23103 27856 23112
rect 27804 23069 27813 23103
rect 27813 23069 27847 23103
rect 27847 23069 27856 23103
rect 27804 23060 27856 23069
rect 28448 23060 28500 23112
rect 36452 23060 36504 23112
rect 41144 23196 41196 23248
rect 45192 23196 45244 23248
rect 38384 23171 38436 23180
rect 38384 23137 38393 23171
rect 38393 23137 38427 23171
rect 38427 23137 38436 23171
rect 38384 23128 38436 23137
rect 38936 23128 38988 23180
rect 40592 23128 40644 23180
rect 43352 23128 43404 23180
rect 37740 23103 37792 23112
rect 37740 23069 37749 23103
rect 37749 23069 37783 23103
rect 37783 23069 37792 23103
rect 37740 23060 37792 23069
rect 42800 23060 42852 23112
rect 40040 22992 40092 23044
rect 40776 22992 40828 23044
rect 41788 22992 41840 23044
rect 42524 22992 42576 23044
rect 44824 23060 44876 23112
rect 48136 23060 48188 23112
rect 44272 22992 44324 23044
rect 47216 23035 47268 23044
rect 47216 23001 47225 23035
rect 47225 23001 47259 23035
rect 47259 23001 47268 23035
rect 47216 22992 47268 23001
rect 37740 22924 37792 22976
rect 43168 22924 43220 22976
rect 45100 22924 45152 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 12716 22720 12768 22772
rect 3884 22652 3936 22704
rect 12072 22652 12124 22704
rect 12440 22652 12492 22704
rect 16764 22720 16816 22772
rect 15384 22652 15436 22704
rect 22744 22720 22796 22772
rect 26240 22763 26292 22772
rect 26240 22729 26249 22763
rect 26249 22729 26283 22763
rect 26283 22729 26292 22763
rect 26240 22720 26292 22729
rect 27160 22720 27212 22772
rect 28448 22720 28500 22772
rect 22836 22695 22888 22704
rect 22836 22661 22845 22695
rect 22845 22661 22879 22695
rect 22879 22661 22888 22695
rect 22836 22652 22888 22661
rect 11520 22627 11572 22636
rect 11520 22593 11529 22627
rect 11529 22593 11563 22627
rect 11563 22593 11572 22627
rect 11520 22584 11572 22593
rect 14372 22627 14424 22636
rect 14372 22593 14381 22627
rect 14381 22593 14415 22627
rect 14415 22593 14424 22627
rect 14372 22584 14424 22593
rect 21456 22584 21508 22636
rect 8668 22559 8720 22568
rect 8668 22525 8677 22559
rect 8677 22525 8711 22559
rect 8711 22525 8720 22559
rect 8668 22516 8720 22525
rect 11796 22559 11848 22568
rect 11796 22525 11805 22559
rect 11805 22525 11839 22559
rect 11839 22525 11848 22559
rect 11796 22516 11848 22525
rect 16580 22516 16632 22568
rect 17776 22559 17828 22568
rect 17776 22525 17785 22559
rect 17785 22525 17819 22559
rect 17819 22525 17828 22559
rect 17776 22516 17828 22525
rect 19064 22559 19116 22568
rect 19064 22525 19073 22559
rect 19073 22525 19107 22559
rect 19107 22525 19116 22559
rect 19064 22516 19116 22525
rect 22468 22584 22520 22636
rect 25780 22652 25832 22704
rect 28080 22652 28132 22704
rect 28816 22652 28868 22704
rect 23572 22584 23624 22636
rect 34704 22627 34756 22636
rect 22192 22448 22244 22500
rect 22284 22448 22336 22500
rect 22652 22448 22704 22500
rect 34704 22593 34713 22627
rect 34713 22593 34747 22627
rect 34747 22593 34756 22627
rect 34704 22584 34756 22593
rect 37740 22720 37792 22772
rect 39488 22763 39540 22772
rect 39488 22729 39497 22763
rect 39497 22729 39531 22763
rect 39531 22729 39540 22763
rect 39488 22720 39540 22729
rect 40776 22763 40828 22772
rect 40776 22729 40785 22763
rect 40785 22729 40819 22763
rect 40819 22729 40828 22763
rect 40776 22720 40828 22729
rect 42524 22720 42576 22772
rect 44272 22763 44324 22772
rect 44272 22729 44281 22763
rect 44281 22729 44315 22763
rect 44315 22729 44324 22763
rect 44272 22720 44324 22729
rect 45652 22763 45704 22772
rect 45652 22729 45661 22763
rect 45661 22729 45695 22763
rect 45695 22729 45704 22763
rect 45652 22720 45704 22729
rect 45744 22652 45796 22704
rect 36452 22627 36504 22636
rect 36452 22593 36461 22627
rect 36461 22593 36495 22627
rect 36495 22593 36504 22627
rect 36452 22584 36504 22593
rect 39764 22584 39816 22636
rect 24492 22559 24544 22568
rect 24492 22525 24501 22559
rect 24501 22525 24535 22559
rect 24535 22525 24544 22559
rect 24492 22516 24544 22525
rect 24768 22559 24820 22568
rect 24768 22525 24777 22559
rect 24777 22525 24811 22559
rect 24811 22525 24820 22559
rect 24768 22516 24820 22525
rect 27528 22559 27580 22568
rect 27528 22525 27537 22559
rect 27537 22525 27571 22559
rect 27571 22525 27580 22559
rect 27528 22516 27580 22525
rect 42984 22627 43036 22636
rect 42984 22593 42993 22627
rect 42993 22593 43027 22627
rect 43027 22593 43036 22627
rect 42984 22584 43036 22593
rect 43168 22627 43220 22636
rect 43168 22593 43177 22627
rect 43177 22593 43211 22627
rect 43211 22593 43220 22627
rect 43168 22584 43220 22593
rect 45100 22627 45152 22636
rect 42800 22516 42852 22568
rect 28908 22448 28960 22500
rect 45100 22593 45109 22627
rect 45109 22593 45143 22627
rect 45143 22593 45152 22627
rect 45100 22584 45152 22593
rect 45560 22627 45612 22636
rect 45560 22593 45569 22627
rect 45569 22593 45603 22627
rect 45603 22593 45612 22627
rect 45560 22584 45612 22593
rect 47584 22627 47636 22636
rect 47584 22593 47593 22627
rect 47593 22593 47627 22627
rect 47627 22593 47636 22627
rect 47584 22584 47636 22593
rect 46204 22559 46256 22568
rect 46204 22525 46213 22559
rect 46213 22525 46247 22559
rect 46247 22525 46256 22559
rect 46204 22516 46256 22525
rect 46480 22559 46532 22568
rect 46480 22525 46489 22559
rect 46489 22525 46523 22559
rect 46523 22525 46532 22559
rect 46480 22516 46532 22525
rect 47860 22559 47912 22568
rect 47860 22525 47869 22559
rect 47869 22525 47903 22559
rect 47903 22525 47912 22559
rect 47860 22516 47912 22525
rect 23480 22380 23532 22432
rect 34520 22423 34572 22432
rect 34520 22389 34529 22423
rect 34529 22389 34563 22423
rect 34563 22389 34572 22423
rect 34520 22380 34572 22389
rect 36636 22423 36688 22432
rect 36636 22389 36645 22423
rect 36645 22389 36679 22423
rect 36679 22389 36688 22423
rect 36636 22380 36688 22389
rect 39488 22380 39540 22432
rect 40040 22380 40092 22432
rect 45928 22380 45980 22432
rect 46664 22380 46716 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 8668 22176 8720 22228
rect 13176 22176 13228 22228
rect 14280 22176 14332 22228
rect 14464 22176 14516 22228
rect 17776 22219 17828 22228
rect 17776 22185 17785 22219
rect 17785 22185 17819 22219
rect 17819 22185 17828 22219
rect 17776 22176 17828 22185
rect 19984 22176 20036 22228
rect 21732 22176 21784 22228
rect 23940 22176 23992 22228
rect 24492 22219 24544 22228
rect 24492 22185 24501 22219
rect 24501 22185 24535 22219
rect 24535 22185 24544 22219
rect 24492 22176 24544 22185
rect 27528 22176 27580 22228
rect 34704 22219 34756 22228
rect 34704 22185 34713 22219
rect 34713 22185 34747 22219
rect 34747 22185 34756 22219
rect 34704 22176 34756 22185
rect 34796 22176 34848 22228
rect 45192 22176 45244 22228
rect 48136 22176 48188 22228
rect 8944 22015 8996 22024
rect 8944 21981 8953 22015
rect 8953 21981 8987 22015
rect 8987 21981 8996 22015
rect 10784 22040 10836 22092
rect 8944 21972 8996 21981
rect 11796 22040 11848 22092
rect 12440 22040 12492 22092
rect 13728 22040 13780 22092
rect 12256 21972 12308 22024
rect 13176 21972 13228 22024
rect 13268 22015 13320 22024
rect 13268 21981 13277 22015
rect 13277 21981 13311 22015
rect 13311 21981 13320 22015
rect 14004 22040 14056 22092
rect 14372 22108 14424 22160
rect 17868 22108 17920 22160
rect 43076 22151 43128 22160
rect 19248 22040 19300 22092
rect 19984 22040 20036 22092
rect 43076 22117 43085 22151
rect 43085 22117 43119 22151
rect 43119 22117 43128 22151
rect 43076 22108 43128 22117
rect 45928 22108 45980 22160
rect 16396 22015 16448 22024
rect 13268 21972 13320 21981
rect 16396 21981 16405 22015
rect 16405 21981 16439 22015
rect 16439 21981 16448 22015
rect 16396 21972 16448 21981
rect 17684 22015 17736 22024
rect 17684 21981 17693 22015
rect 17693 21981 17727 22015
rect 17727 21981 17736 22015
rect 17684 21972 17736 21981
rect 19340 21972 19392 22024
rect 20444 22015 20496 22024
rect 20444 21981 20453 22015
rect 20453 21981 20487 22015
rect 20487 21981 20496 22015
rect 20444 21972 20496 21981
rect 12532 21904 12584 21956
rect 15936 21947 15988 21956
rect 15936 21913 15945 21947
rect 15945 21913 15979 21947
rect 15979 21913 15988 21947
rect 15936 21904 15988 21913
rect 20076 21904 20128 21956
rect 22008 21972 22060 22024
rect 22652 22015 22704 22024
rect 22100 21904 22152 21956
rect 22284 21904 22336 21956
rect 22652 21981 22661 22015
rect 22661 21981 22695 22015
rect 22695 21981 22704 22015
rect 22652 21972 22704 21981
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 23480 22015 23532 22024
rect 23480 21981 23489 22015
rect 23489 21981 23523 22015
rect 23523 21981 23532 22015
rect 23480 21972 23532 21981
rect 25780 22040 25832 22092
rect 25872 22040 25924 22092
rect 24676 21972 24728 22024
rect 25504 22015 25556 22024
rect 25504 21981 25513 22015
rect 25513 21981 25547 22015
rect 25547 21981 25556 22015
rect 25504 21972 25556 21981
rect 11520 21836 11572 21888
rect 13268 21836 13320 21888
rect 14648 21836 14700 21888
rect 16580 21879 16632 21888
rect 16580 21845 16589 21879
rect 16589 21845 16623 21879
rect 16623 21845 16632 21879
rect 16580 21836 16632 21845
rect 17040 21836 17092 21888
rect 19432 21836 19484 21888
rect 21088 21879 21140 21888
rect 21088 21845 21097 21879
rect 21097 21845 21131 21879
rect 21131 21845 21140 21879
rect 21088 21836 21140 21845
rect 22468 21836 22520 21888
rect 24308 21904 24360 21956
rect 26976 21972 27028 22024
rect 27804 21972 27856 22024
rect 29368 21972 29420 22024
rect 25872 21904 25924 21956
rect 29736 21972 29788 22024
rect 31208 21972 31260 22024
rect 32404 21947 32456 21956
rect 32404 21913 32413 21947
rect 32413 21913 32447 21947
rect 32447 21913 32456 21947
rect 32404 21904 32456 21913
rect 23112 21836 23164 21888
rect 23388 21879 23440 21888
rect 23388 21845 23397 21879
rect 23397 21845 23431 21879
rect 23431 21845 23440 21879
rect 23388 21836 23440 21845
rect 23572 21836 23624 21888
rect 28816 21879 28868 21888
rect 28816 21845 28825 21879
rect 28825 21845 28859 21879
rect 28859 21845 28868 21879
rect 28816 21836 28868 21845
rect 29460 21836 29512 21888
rect 30380 21879 30432 21888
rect 30380 21845 30389 21879
rect 30389 21845 30423 21879
rect 30423 21845 30432 21879
rect 30380 21836 30432 21845
rect 35348 21972 35400 22024
rect 36360 21972 36412 22024
rect 36636 21972 36688 22024
rect 37740 21972 37792 22024
rect 37004 21904 37056 21956
rect 38844 21972 38896 22024
rect 39764 21972 39816 22024
rect 40040 22015 40092 22024
rect 40040 21981 40049 22015
rect 40049 21981 40083 22015
rect 40083 21981 40092 22015
rect 40040 21972 40092 21981
rect 42432 21972 42484 22024
rect 45192 22015 45244 22024
rect 45192 21981 45201 22015
rect 45201 21981 45235 22015
rect 45235 21981 45244 22015
rect 45192 21972 45244 21981
rect 45376 22015 45428 22024
rect 45376 21981 45385 22015
rect 45385 21981 45419 22015
rect 45419 21981 45428 22015
rect 45376 21972 45428 21981
rect 45836 22015 45888 22024
rect 45836 21981 45845 22015
rect 45845 21981 45879 22015
rect 45879 21981 45888 22015
rect 45836 21972 45888 21981
rect 40316 21904 40368 21956
rect 42708 21947 42760 21956
rect 42708 21913 42717 21947
rect 42717 21913 42751 21947
rect 42751 21913 42760 21947
rect 42708 21904 42760 21913
rect 38292 21836 38344 21888
rect 38568 21836 38620 21888
rect 45560 21904 45612 21956
rect 45744 21904 45796 21956
rect 46572 21904 46624 21956
rect 47216 21904 47268 21956
rect 43168 21879 43220 21888
rect 43168 21845 43177 21879
rect 43177 21845 43211 21879
rect 43211 21845 43220 21879
rect 43168 21836 43220 21845
rect 46664 21836 46716 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 11704 21675 11756 21684
rect 11704 21641 11713 21675
rect 11713 21641 11747 21675
rect 11747 21641 11756 21675
rect 11704 21632 11756 21641
rect 20444 21632 20496 21684
rect 3792 21428 3844 21480
rect 10876 21496 10928 21548
rect 11520 21539 11572 21548
rect 11520 21505 11529 21539
rect 11529 21505 11563 21539
rect 11563 21505 11572 21539
rect 11520 21496 11572 21505
rect 12256 21539 12308 21548
rect 12256 21505 12265 21539
rect 12265 21505 12299 21539
rect 12299 21505 12308 21539
rect 12256 21496 12308 21505
rect 13728 21564 13780 21616
rect 17684 21564 17736 21616
rect 19984 21564 20036 21616
rect 21088 21564 21140 21616
rect 12624 21428 12676 21480
rect 10416 21360 10468 21412
rect 16396 21496 16448 21548
rect 19432 21539 19484 21548
rect 13544 21471 13596 21480
rect 13544 21437 13553 21471
rect 13553 21437 13587 21471
rect 13587 21437 13596 21471
rect 13728 21471 13780 21480
rect 13544 21428 13596 21437
rect 13728 21437 13737 21471
rect 13737 21437 13771 21471
rect 13771 21437 13780 21471
rect 13728 21428 13780 21437
rect 19432 21505 19441 21539
rect 19441 21505 19475 21539
rect 19475 21505 19484 21539
rect 19432 21496 19484 21505
rect 24308 21632 24360 21684
rect 24768 21632 24820 21684
rect 27896 21632 27948 21684
rect 28448 21632 28500 21684
rect 21916 21496 21968 21548
rect 22284 21496 22336 21548
rect 23112 21496 23164 21548
rect 23296 21496 23348 21548
rect 23572 21539 23624 21548
rect 23572 21505 23581 21539
rect 23581 21505 23615 21539
rect 23615 21505 23624 21539
rect 23572 21496 23624 21505
rect 23664 21539 23716 21548
rect 23664 21505 23673 21539
rect 23673 21505 23707 21539
rect 23707 21505 23716 21539
rect 23664 21496 23716 21505
rect 23940 21496 23992 21548
rect 30380 21564 30432 21616
rect 25228 21496 25280 21548
rect 25504 21496 25556 21548
rect 27804 21496 27856 21548
rect 27896 21496 27948 21548
rect 21732 21428 21784 21480
rect 28356 21496 28408 21548
rect 28816 21539 28868 21548
rect 28816 21505 28825 21539
rect 28825 21505 28859 21539
rect 28859 21505 28868 21539
rect 28816 21496 28868 21505
rect 29000 21539 29052 21548
rect 29000 21505 29009 21539
rect 29009 21505 29043 21539
rect 29043 21505 29052 21539
rect 29000 21496 29052 21505
rect 29460 21539 29512 21548
rect 29460 21505 29469 21539
rect 29469 21505 29503 21539
rect 29503 21505 29512 21539
rect 29460 21496 29512 21505
rect 34520 21632 34572 21684
rect 33416 21564 33468 21616
rect 34612 21607 34664 21616
rect 34612 21573 34621 21607
rect 34621 21573 34655 21607
rect 34655 21573 34664 21607
rect 34612 21564 34664 21573
rect 42800 21632 42852 21684
rect 42892 21632 42944 21684
rect 34796 21564 34848 21616
rect 38200 21564 38252 21616
rect 36360 21539 36412 21548
rect 28172 21428 28224 21480
rect 30104 21428 30156 21480
rect 31208 21471 31260 21480
rect 31208 21437 31217 21471
rect 31217 21437 31251 21471
rect 31251 21437 31260 21471
rect 31208 21428 31260 21437
rect 10692 21292 10744 21344
rect 12348 21335 12400 21344
rect 12348 21301 12357 21335
rect 12357 21301 12391 21335
rect 12391 21301 12400 21335
rect 12348 21292 12400 21301
rect 14464 21360 14516 21412
rect 18144 21360 18196 21412
rect 27344 21360 27396 21412
rect 16856 21292 16908 21344
rect 19340 21292 19392 21344
rect 21456 21292 21508 21344
rect 21548 21292 21600 21344
rect 22560 21292 22612 21344
rect 25504 21335 25556 21344
rect 25504 21301 25513 21335
rect 25513 21301 25547 21335
rect 25547 21301 25556 21335
rect 25504 21292 25556 21301
rect 26976 21292 27028 21344
rect 27988 21292 28040 21344
rect 36360 21505 36369 21539
rect 36369 21505 36403 21539
rect 36403 21505 36412 21539
rect 36360 21496 36412 21505
rect 37740 21539 37792 21548
rect 37740 21505 37749 21539
rect 37749 21505 37783 21539
rect 37783 21505 37792 21539
rect 37740 21496 37792 21505
rect 41696 21539 41748 21548
rect 41696 21505 41705 21539
rect 41705 21505 41739 21539
rect 41739 21505 41748 21539
rect 41696 21496 41748 21505
rect 41880 21539 41932 21548
rect 41880 21505 41889 21539
rect 41889 21505 41923 21539
rect 41923 21505 41932 21539
rect 41880 21496 41932 21505
rect 43076 21496 43128 21548
rect 43628 21539 43680 21548
rect 43628 21505 43637 21539
rect 43637 21505 43671 21539
rect 43671 21505 43680 21539
rect 43628 21496 43680 21505
rect 43812 21539 43864 21548
rect 43812 21505 43821 21539
rect 43821 21505 43855 21539
rect 43855 21505 43864 21539
rect 43812 21496 43864 21505
rect 44272 21496 44324 21548
rect 45836 21632 45888 21684
rect 47584 21632 47636 21684
rect 45376 21564 45428 21616
rect 46664 21607 46716 21616
rect 45744 21496 45796 21548
rect 46664 21573 46673 21607
rect 46673 21573 46707 21607
rect 46707 21573 46716 21607
rect 46664 21564 46716 21573
rect 32864 21428 32916 21480
rect 35532 21428 35584 21480
rect 36268 21428 36320 21480
rect 32312 21360 32364 21412
rect 38292 21471 38344 21480
rect 38292 21437 38301 21471
rect 38301 21437 38335 21471
rect 38335 21437 38344 21471
rect 38292 21428 38344 21437
rect 42708 21428 42760 21480
rect 45008 21471 45060 21480
rect 45008 21437 45017 21471
rect 45017 21437 45051 21471
rect 45051 21437 45060 21471
rect 45008 21428 45060 21437
rect 47676 21496 47728 21548
rect 47860 21539 47912 21548
rect 47860 21505 47869 21539
rect 47869 21505 47903 21539
rect 47903 21505 47912 21539
rect 47860 21496 47912 21505
rect 47768 21428 47820 21480
rect 48136 21632 48188 21684
rect 41880 21360 41932 21412
rect 43812 21360 43864 21412
rect 48136 21403 48188 21412
rect 48136 21369 48145 21403
rect 48145 21369 48179 21403
rect 48179 21369 48188 21403
rect 48136 21360 48188 21369
rect 36636 21335 36688 21344
rect 36636 21301 36645 21335
rect 36645 21301 36679 21335
rect 36679 21301 36688 21335
rect 36636 21292 36688 21301
rect 37004 21292 37056 21344
rect 42892 21292 42944 21344
rect 43076 21335 43128 21344
rect 43076 21301 43085 21335
rect 43085 21301 43119 21335
rect 43119 21301 43128 21335
rect 43076 21292 43128 21301
rect 46020 21335 46072 21344
rect 46020 21301 46029 21335
rect 46029 21301 46063 21335
rect 46063 21301 46072 21335
rect 46020 21292 46072 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2596 21088 2648 21140
rect 10416 21088 10468 21140
rect 12072 21088 12124 21140
rect 12624 21131 12676 21140
rect 12624 21097 12633 21131
rect 12633 21097 12667 21131
rect 12667 21097 12676 21131
rect 12624 21088 12676 21097
rect 13728 21088 13780 21140
rect 16212 21131 16264 21140
rect 16212 21097 16221 21131
rect 16221 21097 16255 21131
rect 16255 21097 16264 21131
rect 16212 21088 16264 21097
rect 16488 21088 16540 21140
rect 16856 21088 16908 21140
rect 23296 21131 23348 21140
rect 3976 21020 4028 21072
rect 10324 21020 10376 21072
rect 14372 21020 14424 21072
rect 23296 21097 23305 21131
rect 23305 21097 23339 21131
rect 23339 21097 23348 21131
rect 23296 21088 23348 21097
rect 24676 21131 24728 21140
rect 24676 21097 24685 21131
rect 24685 21097 24719 21131
rect 24719 21097 24728 21131
rect 24676 21088 24728 21097
rect 27804 21088 27856 21140
rect 28172 21088 28224 21140
rect 28448 21088 28500 21140
rect 30104 21131 30156 21140
rect 30104 21097 30113 21131
rect 30113 21097 30147 21131
rect 30147 21097 30156 21131
rect 30104 21088 30156 21097
rect 32680 21131 32732 21140
rect 32680 21097 32689 21131
rect 32689 21097 32723 21131
rect 32723 21097 32732 21131
rect 32680 21088 32732 21097
rect 33416 21131 33468 21140
rect 33416 21097 33425 21131
rect 33425 21097 33459 21131
rect 33459 21097 33468 21131
rect 33416 21088 33468 21097
rect 36268 21088 36320 21140
rect 42708 21088 42760 21140
rect 3424 20952 3476 21004
rect 14004 20952 14056 21004
rect 20444 20952 20496 21004
rect 21548 20995 21600 21004
rect 21548 20961 21557 20995
rect 21557 20961 21591 20995
rect 21591 20961 21600 20995
rect 21548 20952 21600 20961
rect 25504 20995 25556 21004
rect 25504 20961 25513 20995
rect 25513 20961 25547 20995
rect 25547 20961 25556 20995
rect 25504 20952 25556 20961
rect 10416 20927 10468 20936
rect 10416 20893 10425 20927
rect 10425 20893 10459 20927
rect 10459 20893 10468 20927
rect 10416 20884 10468 20893
rect 12072 20884 12124 20936
rect 12900 20927 12952 20936
rect 10692 20859 10744 20868
rect 10692 20825 10701 20859
rect 10701 20825 10735 20859
rect 10735 20825 10744 20859
rect 10692 20816 10744 20825
rect 12348 20816 12400 20868
rect 12900 20893 12909 20927
rect 12909 20893 12943 20927
rect 12943 20893 12952 20927
rect 12900 20884 12952 20893
rect 14188 20884 14240 20936
rect 12808 20791 12860 20800
rect 12808 20757 12817 20791
rect 12817 20757 12851 20791
rect 12851 20757 12860 20791
rect 12808 20748 12860 20757
rect 14188 20748 14240 20800
rect 14556 20884 14608 20936
rect 16580 20884 16632 20936
rect 17408 20927 17460 20936
rect 17408 20893 17417 20927
rect 17417 20893 17451 20927
rect 17451 20893 17460 20927
rect 17408 20884 17460 20893
rect 18144 20927 18196 20936
rect 18144 20893 18153 20927
rect 18153 20893 18187 20927
rect 18187 20893 18196 20927
rect 18144 20884 18196 20893
rect 19248 20884 19300 20936
rect 21456 20884 21508 20936
rect 23204 20884 23256 20936
rect 25320 20927 25372 20936
rect 25320 20893 25329 20927
rect 25329 20893 25363 20927
rect 25363 20893 25372 20927
rect 25320 20884 25372 20893
rect 14372 20748 14424 20800
rect 22100 20816 22152 20868
rect 22560 20816 22612 20868
rect 28172 20952 28224 21004
rect 28356 20952 28408 21004
rect 31116 20952 31168 21004
rect 31576 20952 31628 21004
rect 32220 21020 32272 21072
rect 35532 21020 35584 21072
rect 42892 21020 42944 21072
rect 27804 20884 27856 20936
rect 17040 20748 17092 20800
rect 17960 20748 18012 20800
rect 18144 20748 18196 20800
rect 18328 20748 18380 20800
rect 18420 20748 18472 20800
rect 27896 20816 27948 20868
rect 28172 20816 28224 20868
rect 28448 20884 28500 20936
rect 31208 20884 31260 20936
rect 32312 20884 32364 20936
rect 31116 20816 31168 20868
rect 27160 20748 27212 20800
rect 29000 20748 29052 20800
rect 30196 20748 30248 20800
rect 31576 20816 31628 20868
rect 32220 20816 32272 20868
rect 43628 21088 43680 21140
rect 46480 21088 46532 21140
rect 45928 21020 45980 21072
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 38568 20884 38620 20936
rect 42984 20884 43036 20936
rect 43076 20884 43128 20936
rect 43720 20884 43772 20936
rect 32864 20816 32916 20868
rect 34796 20816 34848 20868
rect 35348 20859 35400 20868
rect 35348 20825 35357 20859
rect 35357 20825 35391 20859
rect 35391 20825 35400 20859
rect 36268 20859 36320 20868
rect 35348 20816 35400 20825
rect 36268 20825 36277 20859
rect 36277 20825 36311 20859
rect 36311 20825 36320 20859
rect 36268 20816 36320 20825
rect 36820 20791 36872 20800
rect 36820 20757 36829 20791
rect 36829 20757 36863 20791
rect 36863 20757 36872 20791
rect 36820 20748 36872 20757
rect 38844 20748 38896 20800
rect 42892 20748 42944 20800
rect 43628 20748 43680 20800
rect 43812 20748 43864 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 3516 20544 3568 20596
rect 10416 20544 10468 20596
rect 12900 20544 12952 20596
rect 13912 20544 13964 20596
rect 32220 20544 32272 20596
rect 32404 20587 32456 20596
rect 32404 20553 32413 20587
rect 32413 20553 32447 20587
rect 32447 20553 32456 20587
rect 32404 20544 32456 20553
rect 11704 20451 11756 20460
rect 11704 20417 11713 20451
rect 11713 20417 11747 20451
rect 11747 20417 11756 20451
rect 11704 20408 11756 20417
rect 12808 20451 12860 20460
rect 12808 20417 12814 20451
rect 12814 20417 12848 20451
rect 12848 20417 12860 20451
rect 12808 20408 12860 20417
rect 13544 20408 13596 20460
rect 14832 20476 14884 20528
rect 14464 20408 14516 20460
rect 3516 20272 3568 20324
rect 11060 20204 11112 20256
rect 11612 20204 11664 20256
rect 12900 20272 12952 20324
rect 14372 20340 14424 20392
rect 16580 20408 16632 20460
rect 17316 20476 17368 20528
rect 17500 20476 17552 20528
rect 18328 20519 18380 20528
rect 18328 20485 18337 20519
rect 18337 20485 18371 20519
rect 18371 20485 18380 20519
rect 18328 20476 18380 20485
rect 19984 20519 20036 20528
rect 19984 20485 19993 20519
rect 19993 20485 20027 20519
rect 20027 20485 20036 20519
rect 19984 20476 20036 20485
rect 25320 20476 25372 20528
rect 17408 20408 17460 20460
rect 22008 20451 22060 20460
rect 22008 20417 22017 20451
rect 22017 20417 22051 20451
rect 22051 20417 22060 20451
rect 22008 20408 22060 20417
rect 25136 20451 25188 20460
rect 25136 20417 25145 20451
rect 25145 20417 25179 20451
rect 25179 20417 25188 20451
rect 25136 20408 25188 20417
rect 27344 20476 27396 20528
rect 27988 20519 28040 20528
rect 27988 20485 27997 20519
rect 27997 20485 28031 20519
rect 28031 20485 28040 20519
rect 27988 20476 28040 20485
rect 26884 20408 26936 20460
rect 29368 20408 29420 20460
rect 36636 20544 36688 20596
rect 36820 20476 36872 20528
rect 43720 20519 43772 20528
rect 43720 20485 43729 20519
rect 43729 20485 43763 20519
rect 43763 20485 43772 20519
rect 43720 20476 43772 20485
rect 46020 20476 46072 20528
rect 47952 20519 48004 20528
rect 47952 20485 47961 20519
rect 47961 20485 47995 20519
rect 47995 20485 48004 20519
rect 47952 20476 48004 20485
rect 22652 20340 22704 20392
rect 27160 20340 27212 20392
rect 42708 20408 42760 20460
rect 43260 20451 43312 20460
rect 43260 20417 43269 20451
rect 43269 20417 43303 20451
rect 43303 20417 43312 20451
rect 43260 20408 43312 20417
rect 43904 20451 43956 20460
rect 43904 20417 43913 20451
rect 43913 20417 43947 20451
rect 43947 20417 43956 20451
rect 43904 20408 43956 20417
rect 44272 20408 44324 20460
rect 47216 20408 47268 20460
rect 18236 20272 18288 20324
rect 25228 20272 25280 20324
rect 14188 20204 14240 20256
rect 14280 20247 14332 20256
rect 14280 20213 14289 20247
rect 14289 20213 14323 20247
rect 14323 20213 14332 20247
rect 14280 20204 14332 20213
rect 15568 20204 15620 20256
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 15752 20204 15804 20213
rect 17040 20247 17092 20256
rect 17040 20213 17049 20247
rect 17049 20213 17083 20247
rect 17083 20213 17092 20247
rect 17040 20204 17092 20213
rect 22100 20204 22152 20256
rect 25596 20204 25648 20256
rect 25872 20204 25924 20256
rect 29460 20247 29512 20256
rect 29460 20213 29469 20247
rect 29469 20213 29503 20247
rect 29503 20213 29512 20247
rect 29460 20204 29512 20213
rect 33508 20204 33560 20256
rect 34704 20340 34756 20392
rect 35256 20340 35308 20392
rect 43812 20340 43864 20392
rect 45560 20340 45612 20392
rect 36544 20272 36596 20324
rect 38752 20204 38804 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4988 20000 5040 20052
rect 13544 20000 13596 20052
rect 14372 20000 14424 20052
rect 14464 20043 14516 20052
rect 14464 20009 14473 20043
rect 14473 20009 14507 20043
rect 14507 20009 14516 20043
rect 14464 20000 14516 20009
rect 16212 20000 16264 20052
rect 27344 20043 27396 20052
rect 22744 19932 22796 19984
rect 27344 20009 27353 20043
rect 27353 20009 27387 20043
rect 27387 20009 27396 20043
rect 27344 20000 27396 20009
rect 28816 20000 28868 20052
rect 30012 20000 30064 20052
rect 36544 20000 36596 20052
rect 45008 20043 45060 20052
rect 45008 20009 45017 20043
rect 45017 20009 45051 20043
rect 45051 20009 45060 20043
rect 45008 20000 45060 20009
rect 47768 20000 47820 20052
rect 20 19864 72 19916
rect 15752 19907 15804 19916
rect 1768 19796 1820 19848
rect 11060 19839 11112 19848
rect 11060 19805 11069 19839
rect 11069 19805 11103 19839
rect 11103 19805 11112 19839
rect 11060 19796 11112 19805
rect 12624 19796 12676 19848
rect 13820 19796 13872 19848
rect 14556 19796 14608 19848
rect 11612 19728 11664 19780
rect 13544 19728 13596 19780
rect 14188 19728 14240 19780
rect 15752 19873 15761 19907
rect 15761 19873 15795 19907
rect 15795 19873 15804 19907
rect 15752 19864 15804 19873
rect 15384 19796 15436 19848
rect 14280 19703 14332 19712
rect 14280 19669 14305 19703
rect 14305 19669 14332 19703
rect 25596 19907 25648 19916
rect 25596 19873 25605 19907
rect 25605 19873 25639 19907
rect 25639 19873 25648 19907
rect 25596 19864 25648 19873
rect 31300 19932 31352 19984
rect 32220 19932 32272 19984
rect 34704 19975 34756 19984
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 19340 19796 19392 19848
rect 21456 19796 21508 19848
rect 24492 19796 24544 19848
rect 26976 19796 27028 19848
rect 20444 19728 20496 19780
rect 22652 19728 22704 19780
rect 25228 19728 25280 19780
rect 25872 19771 25924 19780
rect 25872 19737 25881 19771
rect 25881 19737 25915 19771
rect 25915 19737 25924 19771
rect 25872 19728 25924 19737
rect 27896 19796 27948 19848
rect 29460 19864 29512 19916
rect 28356 19796 28408 19848
rect 14280 19660 14332 19669
rect 19156 19660 19208 19712
rect 25136 19660 25188 19712
rect 25780 19660 25832 19712
rect 26884 19660 26936 19712
rect 28448 19660 28500 19712
rect 28908 19728 28960 19780
rect 31392 19771 31444 19780
rect 31392 19737 31401 19771
rect 31401 19737 31435 19771
rect 31435 19737 31444 19771
rect 31392 19728 31444 19737
rect 34704 19941 34713 19975
rect 34713 19941 34747 19975
rect 34747 19941 34756 19975
rect 34704 19932 34756 19941
rect 43904 19932 43956 19984
rect 47032 19932 47084 19984
rect 35900 19907 35952 19916
rect 32312 19796 32364 19848
rect 33048 19796 33100 19848
rect 35900 19873 35909 19907
rect 35909 19873 35943 19907
rect 35943 19873 35952 19907
rect 35900 19864 35952 19873
rect 32220 19771 32272 19780
rect 32220 19737 32229 19771
rect 32229 19737 32263 19771
rect 32263 19737 32272 19771
rect 32220 19728 32272 19737
rect 32956 19728 33008 19780
rect 34704 19728 34756 19780
rect 43260 19796 43312 19848
rect 43996 19839 44048 19848
rect 43996 19805 44005 19839
rect 44005 19805 44039 19839
rect 44039 19805 44048 19839
rect 43996 19796 44048 19805
rect 42708 19728 42760 19780
rect 37372 19660 37424 19712
rect 46940 19864 46992 19916
rect 47952 19864 48004 19916
rect 45836 19839 45888 19848
rect 45836 19805 45845 19839
rect 45845 19805 45879 19839
rect 45879 19805 45888 19839
rect 45836 19796 45888 19805
rect 46112 19796 46164 19848
rect 47400 19839 47452 19848
rect 47400 19805 47409 19839
rect 47409 19805 47443 19839
rect 47443 19805 47452 19839
rect 47400 19796 47452 19805
rect 45744 19728 45796 19780
rect 45928 19660 45980 19712
rect 48044 19728 48096 19780
rect 46572 19660 46624 19712
rect 46940 19660 46992 19712
rect 47492 19703 47544 19712
rect 47492 19669 47501 19703
rect 47501 19669 47535 19703
rect 47535 19669 47544 19703
rect 47492 19660 47544 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 14924 19456 14976 19508
rect 20444 19499 20496 19508
rect 20444 19465 20453 19499
rect 20453 19465 20487 19499
rect 20487 19465 20496 19499
rect 20444 19456 20496 19465
rect 22836 19456 22888 19508
rect 24492 19499 24544 19508
rect 12900 19431 12952 19440
rect 12900 19397 12909 19431
rect 12909 19397 12943 19431
rect 12943 19397 12952 19431
rect 12900 19388 12952 19397
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 11520 19320 11572 19372
rect 14372 19388 14424 19440
rect 15016 19388 15068 19440
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 14740 19320 14792 19372
rect 14832 19320 14884 19372
rect 19156 19320 19208 19372
rect 22652 19320 22704 19372
rect 24124 19320 24176 19372
rect 24492 19465 24501 19499
rect 24501 19465 24535 19499
rect 24535 19465 24544 19499
rect 24492 19456 24544 19465
rect 28908 19499 28960 19508
rect 28908 19465 28917 19499
rect 28917 19465 28951 19499
rect 28951 19465 28960 19499
rect 28908 19456 28960 19465
rect 43904 19456 43956 19508
rect 46020 19456 46072 19508
rect 29000 19388 29052 19440
rect 30288 19388 30340 19440
rect 33508 19431 33560 19440
rect 33508 19397 33517 19431
rect 33517 19397 33551 19431
rect 33551 19397 33560 19431
rect 33508 19388 33560 19397
rect 36636 19388 36688 19440
rect 28264 19320 28316 19372
rect 28908 19320 28960 19372
rect 33048 19320 33100 19372
rect 33324 19363 33376 19372
rect 33324 19329 33333 19363
rect 33333 19329 33367 19363
rect 33367 19329 33376 19363
rect 33324 19320 33376 19329
rect 37096 19320 37148 19372
rect 42708 19320 42760 19372
rect 43996 19320 44048 19372
rect 45928 19363 45980 19372
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 3424 19116 3476 19168
rect 17224 19252 17276 19304
rect 17776 19295 17828 19304
rect 17776 19261 17785 19295
rect 17785 19261 17819 19295
rect 17819 19261 17828 19295
rect 17776 19252 17828 19261
rect 18236 19252 18288 19304
rect 22744 19295 22796 19304
rect 22744 19261 22753 19295
rect 22753 19261 22787 19295
rect 22787 19261 22796 19295
rect 22744 19252 22796 19261
rect 23664 19252 23716 19304
rect 32588 19295 32640 19304
rect 32588 19261 32597 19295
rect 32597 19261 32631 19295
rect 32631 19261 32640 19295
rect 32588 19252 32640 19261
rect 45928 19329 45937 19363
rect 45937 19329 45971 19363
rect 45971 19329 45980 19363
rect 45928 19320 45980 19329
rect 46112 19320 46164 19372
rect 46572 19363 46624 19372
rect 46572 19329 46581 19363
rect 46581 19329 46615 19363
rect 46615 19329 46624 19363
rect 46572 19320 46624 19329
rect 46664 19320 46716 19372
rect 12808 19116 12860 19168
rect 13912 19116 13964 19168
rect 14832 19116 14884 19168
rect 20720 19116 20772 19168
rect 45744 19184 45796 19236
rect 35624 19159 35676 19168
rect 35624 19125 35633 19159
rect 35633 19125 35667 19159
rect 35667 19125 35676 19159
rect 35624 19116 35676 19125
rect 45468 19159 45520 19168
rect 45468 19125 45477 19159
rect 45477 19125 45511 19159
rect 45511 19125 45520 19159
rect 45468 19116 45520 19125
rect 46204 19159 46256 19168
rect 46204 19125 46213 19159
rect 46213 19125 46247 19159
rect 46247 19125 46256 19159
rect 46204 19116 46256 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 17776 18912 17828 18964
rect 23664 18955 23716 18964
rect 23664 18921 23673 18955
rect 23673 18921 23707 18955
rect 23707 18921 23716 18955
rect 23664 18912 23716 18921
rect 30932 18912 30984 18964
rect 31484 18912 31536 18964
rect 32588 18912 32640 18964
rect 1584 18776 1636 18828
rect 15568 18776 15620 18828
rect 2320 18708 2372 18760
rect 6552 18708 6604 18760
rect 12808 18708 12860 18760
rect 13820 18708 13872 18760
rect 14924 18751 14976 18760
rect 14924 18717 14933 18751
rect 14933 18717 14967 18751
rect 14967 18717 14976 18751
rect 14924 18708 14976 18717
rect 15016 18708 15068 18760
rect 17592 18776 17644 18828
rect 18052 18776 18104 18828
rect 20720 18819 20772 18828
rect 20720 18785 20729 18819
rect 20729 18785 20763 18819
rect 20763 18785 20772 18819
rect 20720 18776 20772 18785
rect 31116 18844 31168 18896
rect 31668 18844 31720 18896
rect 33048 18844 33100 18896
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 22836 18751 22888 18760
rect 1584 18572 1636 18624
rect 17500 18640 17552 18692
rect 22836 18717 22845 18751
rect 22845 18717 22879 18751
rect 22879 18717 22888 18751
rect 22836 18708 22888 18717
rect 23572 18751 23624 18760
rect 23572 18717 23581 18751
rect 23581 18717 23615 18751
rect 23615 18717 23624 18751
rect 23572 18708 23624 18717
rect 27252 18751 27304 18760
rect 27252 18717 27261 18751
rect 27261 18717 27295 18751
rect 27295 18717 27304 18751
rect 27252 18708 27304 18717
rect 30932 18708 30984 18760
rect 31116 18751 31168 18760
rect 31116 18717 31125 18751
rect 31125 18717 31159 18751
rect 31159 18717 31168 18751
rect 31300 18751 31352 18760
rect 31116 18708 31168 18717
rect 31300 18717 31309 18751
rect 31309 18717 31343 18751
rect 31343 18717 31352 18751
rect 31300 18708 31352 18717
rect 22008 18640 22060 18692
rect 22928 18640 22980 18692
rect 27712 18640 27764 18692
rect 31484 18708 31536 18760
rect 13084 18572 13136 18624
rect 14096 18572 14148 18624
rect 14740 18615 14792 18624
rect 14740 18581 14749 18615
rect 14749 18581 14783 18615
rect 14783 18581 14792 18615
rect 14740 18572 14792 18581
rect 23020 18615 23072 18624
rect 23020 18581 23029 18615
rect 23029 18581 23063 18615
rect 23063 18581 23072 18615
rect 23020 18572 23072 18581
rect 31208 18572 31260 18624
rect 31668 18640 31720 18692
rect 32404 18708 32456 18760
rect 32956 18751 33008 18760
rect 32956 18717 32965 18751
rect 32965 18717 32999 18751
rect 32999 18717 33008 18751
rect 32956 18708 33008 18717
rect 33600 18751 33652 18760
rect 33600 18717 33609 18751
rect 33609 18717 33643 18751
rect 33643 18717 33652 18751
rect 33600 18708 33652 18717
rect 46112 18844 46164 18896
rect 43812 18776 43864 18828
rect 45468 18776 45520 18828
rect 47492 18776 47544 18828
rect 48136 18819 48188 18828
rect 48136 18785 48145 18819
rect 48145 18785 48179 18819
rect 48179 18785 48188 18819
rect 48136 18776 48188 18785
rect 36912 18640 36964 18692
rect 37372 18708 37424 18760
rect 45100 18751 45152 18760
rect 42800 18683 42852 18692
rect 32312 18572 32364 18624
rect 37464 18615 37516 18624
rect 37464 18581 37473 18615
rect 37473 18581 37507 18615
rect 37507 18581 37516 18615
rect 37464 18572 37516 18581
rect 42800 18649 42809 18683
rect 42809 18649 42843 18683
rect 42843 18649 42852 18683
rect 42800 18640 42852 18649
rect 44456 18683 44508 18692
rect 44456 18649 44465 18683
rect 44465 18649 44499 18683
rect 44499 18649 44508 18683
rect 44456 18640 44508 18649
rect 45100 18717 45109 18751
rect 45109 18717 45143 18751
rect 45143 18717 45152 18751
rect 45100 18708 45152 18717
rect 45376 18708 45428 18760
rect 45744 18640 45796 18692
rect 44364 18572 44416 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 4620 18368 4672 18420
rect 31300 18411 31352 18420
rect 14096 18300 14148 18352
rect 17224 18343 17276 18352
rect 17224 18309 17233 18343
rect 17233 18309 17267 18343
rect 17267 18309 17276 18343
rect 17224 18300 17276 18309
rect 22560 18300 22612 18352
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 17132 18275 17184 18284
rect 17132 18241 17141 18275
rect 17141 18241 17175 18275
rect 17175 18241 17184 18275
rect 17132 18232 17184 18241
rect 17960 18232 18012 18284
rect 18052 18275 18104 18284
rect 18052 18241 18061 18275
rect 18061 18241 18095 18275
rect 18095 18241 18104 18275
rect 18052 18232 18104 18241
rect 14740 18164 14792 18216
rect 15016 18164 15068 18216
rect 17868 18071 17920 18080
rect 17868 18037 17877 18071
rect 17877 18037 17911 18071
rect 17911 18037 17920 18071
rect 17868 18028 17920 18037
rect 24768 18232 24820 18284
rect 28816 18300 28868 18352
rect 31300 18377 31309 18411
rect 31309 18377 31343 18411
rect 31343 18377 31352 18411
rect 31300 18368 31352 18377
rect 31484 18368 31536 18420
rect 37096 18411 37148 18420
rect 25780 18232 25832 18284
rect 27160 18275 27212 18284
rect 27160 18241 27169 18275
rect 27169 18241 27203 18275
rect 27203 18241 27212 18275
rect 27160 18232 27212 18241
rect 22100 18207 22152 18216
rect 22100 18173 22109 18207
rect 22109 18173 22143 18207
rect 22143 18173 22152 18207
rect 22100 18164 22152 18173
rect 22468 18164 22520 18216
rect 23572 18164 23624 18216
rect 26976 18207 27028 18216
rect 26976 18173 26985 18207
rect 26985 18173 27019 18207
rect 27019 18173 27028 18207
rect 26976 18164 27028 18173
rect 27252 18164 27304 18216
rect 29000 18232 29052 18284
rect 30380 18300 30432 18352
rect 31208 18343 31260 18352
rect 31208 18309 31217 18343
rect 31217 18309 31251 18343
rect 31251 18309 31260 18343
rect 31208 18300 31260 18309
rect 30656 18232 30708 18284
rect 31576 18275 31628 18284
rect 31576 18241 31585 18275
rect 31585 18241 31619 18275
rect 31619 18241 31628 18275
rect 37096 18377 37105 18411
rect 37105 18377 37139 18411
rect 37139 18377 37148 18411
rect 37096 18368 37148 18377
rect 35624 18300 35676 18352
rect 31576 18232 31628 18241
rect 33324 18232 33376 18284
rect 37372 18368 37424 18420
rect 42800 18411 42852 18420
rect 42800 18377 42809 18411
rect 42809 18377 42843 18411
rect 42843 18377 42852 18411
rect 42800 18368 42852 18377
rect 45100 18368 45152 18420
rect 37464 18343 37516 18352
rect 37464 18309 37473 18343
rect 37473 18309 37507 18343
rect 37507 18309 37516 18343
rect 37464 18300 37516 18309
rect 37556 18300 37608 18352
rect 41788 18300 41840 18352
rect 46204 18300 46256 18352
rect 47032 18300 47084 18352
rect 31300 18164 31352 18216
rect 33600 18164 33652 18216
rect 35900 18207 35952 18216
rect 35900 18173 35909 18207
rect 35909 18173 35943 18207
rect 35943 18173 35952 18207
rect 35900 18164 35952 18173
rect 37188 18164 37240 18216
rect 27896 18096 27948 18148
rect 34796 18096 34848 18148
rect 37096 18096 37148 18148
rect 37464 18164 37516 18216
rect 38384 18164 38436 18216
rect 44364 18232 44416 18284
rect 46756 18232 46808 18284
rect 43904 18207 43956 18216
rect 22468 18028 22520 18080
rect 22652 18028 22704 18080
rect 24860 18028 24912 18080
rect 27804 18071 27856 18080
rect 27804 18037 27813 18071
rect 27813 18037 27847 18071
rect 27847 18037 27856 18071
rect 27804 18028 27856 18037
rect 28816 18071 28868 18080
rect 28816 18037 28825 18071
rect 28825 18037 28859 18071
rect 28859 18037 28868 18071
rect 28816 18028 28868 18037
rect 31484 18028 31536 18080
rect 32312 18028 32364 18080
rect 33048 18071 33100 18080
rect 33048 18037 33057 18071
rect 33057 18037 33091 18071
rect 33091 18037 33100 18071
rect 33048 18028 33100 18037
rect 36912 18071 36964 18080
rect 36912 18037 36921 18071
rect 36921 18037 36955 18071
rect 36955 18037 36964 18071
rect 36912 18028 36964 18037
rect 37464 18028 37516 18080
rect 43904 18173 43913 18207
rect 43913 18173 43947 18207
rect 43947 18173 43956 18207
rect 43904 18164 43956 18173
rect 44732 18207 44784 18216
rect 44732 18173 44741 18207
rect 44741 18173 44775 18207
rect 44775 18173 44784 18207
rect 44732 18164 44784 18173
rect 41788 18096 41840 18148
rect 45560 18096 45612 18148
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3056 17824 3108 17876
rect 9772 17824 9824 17876
rect 17040 17824 17092 17876
rect 17592 17824 17644 17876
rect 18328 17824 18380 17876
rect 22100 17824 22152 17876
rect 22560 17867 22612 17876
rect 22560 17833 22569 17867
rect 22569 17833 22603 17867
rect 22603 17833 22612 17867
rect 22560 17824 22612 17833
rect 17776 17756 17828 17808
rect 18236 17756 18288 17808
rect 22284 17756 22336 17808
rect 12808 17663 12860 17672
rect 12808 17629 12817 17663
rect 12817 17629 12851 17663
rect 12851 17629 12860 17663
rect 12808 17620 12860 17629
rect 13820 17620 13872 17672
rect 14832 17620 14884 17672
rect 15384 17552 15436 17604
rect 16764 17620 16816 17672
rect 17592 17552 17644 17604
rect 17776 17552 17828 17604
rect 18328 17620 18380 17672
rect 20536 17620 20588 17672
rect 22652 17688 22704 17740
rect 24860 17688 24912 17740
rect 26148 17824 26200 17876
rect 25596 17688 25648 17740
rect 23020 17620 23072 17672
rect 23388 17620 23440 17672
rect 23572 17663 23624 17672
rect 23572 17629 23581 17663
rect 23581 17629 23615 17663
rect 23615 17629 23624 17663
rect 23572 17620 23624 17629
rect 27160 17824 27212 17876
rect 28724 17824 28776 17876
rect 31300 17824 31352 17876
rect 34796 17824 34848 17876
rect 37464 17824 37516 17876
rect 44272 17824 44324 17876
rect 35440 17756 35492 17808
rect 44180 17756 44232 17808
rect 27804 17688 27856 17740
rect 31576 17688 31628 17740
rect 37096 17688 37148 17740
rect 43904 17688 43956 17740
rect 47492 17688 47544 17740
rect 12624 17484 12676 17536
rect 13452 17527 13504 17536
rect 13452 17493 13461 17527
rect 13461 17493 13495 17527
rect 13495 17493 13504 17527
rect 13452 17484 13504 17493
rect 15292 17527 15344 17536
rect 15292 17493 15301 17527
rect 15301 17493 15335 17527
rect 15335 17493 15344 17527
rect 15292 17484 15344 17493
rect 16856 17484 16908 17536
rect 19248 17552 19300 17604
rect 25872 17552 25924 17604
rect 29000 17620 29052 17672
rect 30380 17663 30432 17672
rect 30380 17629 30389 17663
rect 30389 17629 30423 17663
rect 30423 17629 30432 17663
rect 30380 17620 30432 17629
rect 30656 17620 30708 17672
rect 31116 17663 31168 17672
rect 31116 17629 31125 17663
rect 31125 17629 31159 17663
rect 31159 17629 31168 17663
rect 31116 17620 31168 17629
rect 31300 17663 31352 17672
rect 31300 17629 31309 17663
rect 31309 17629 31343 17663
rect 31343 17629 31352 17663
rect 31300 17620 31352 17629
rect 31484 17620 31536 17672
rect 32312 17663 32364 17672
rect 32312 17629 32321 17663
rect 32321 17629 32355 17663
rect 32355 17629 32364 17663
rect 32312 17620 32364 17629
rect 32864 17620 32916 17672
rect 35440 17663 35492 17672
rect 35440 17629 35449 17663
rect 35449 17629 35483 17663
rect 35483 17629 35492 17663
rect 35440 17620 35492 17629
rect 36176 17663 36228 17672
rect 36176 17629 36185 17663
rect 36185 17629 36219 17663
rect 36219 17629 36228 17663
rect 36176 17620 36228 17629
rect 45100 17620 45152 17672
rect 45376 17663 45428 17672
rect 45376 17629 45385 17663
rect 45385 17629 45419 17663
rect 45419 17629 45428 17663
rect 45376 17620 45428 17629
rect 26792 17552 26844 17604
rect 18236 17527 18288 17536
rect 18236 17493 18245 17527
rect 18245 17493 18279 17527
rect 18279 17493 18288 17527
rect 18236 17484 18288 17493
rect 24124 17484 24176 17536
rect 24952 17527 25004 17536
rect 24952 17493 24961 17527
rect 24961 17493 24995 17527
rect 24995 17493 25004 17527
rect 24952 17484 25004 17493
rect 25412 17484 25464 17536
rect 28816 17552 28868 17604
rect 30932 17552 30984 17604
rect 46296 17552 46348 17604
rect 46940 17552 46992 17604
rect 48136 17595 48188 17604
rect 48136 17561 48145 17595
rect 48145 17561 48179 17595
rect 48179 17561 48188 17595
rect 48136 17552 48188 17561
rect 27620 17484 27672 17536
rect 29644 17527 29696 17536
rect 29644 17493 29653 17527
rect 29653 17493 29687 17527
rect 29687 17493 29696 17527
rect 29644 17484 29696 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 18052 17280 18104 17332
rect 24768 17280 24820 17332
rect 26976 17280 27028 17332
rect 27712 17280 27764 17332
rect 31484 17323 31536 17332
rect 31484 17289 31493 17323
rect 31493 17289 31527 17323
rect 31527 17289 31536 17323
rect 31484 17280 31536 17289
rect 45376 17280 45428 17332
rect 46940 17323 46992 17332
rect 46940 17289 46949 17323
rect 46949 17289 46983 17323
rect 46983 17289 46992 17323
rect 46940 17280 46992 17289
rect 12624 17212 12676 17264
rect 13452 17212 13504 17264
rect 16856 17212 16908 17264
rect 17868 17255 17920 17264
rect 12716 17119 12768 17128
rect 12716 17085 12725 17119
rect 12725 17085 12759 17119
rect 12759 17085 12768 17119
rect 12716 17076 12768 17085
rect 12808 17076 12860 17128
rect 17132 17076 17184 17128
rect 1400 16940 1452 16992
rect 13360 16940 13412 16992
rect 14188 16983 14240 16992
rect 14188 16949 14197 16983
rect 14197 16949 14231 16983
rect 14231 16949 14240 16983
rect 14188 16940 14240 16949
rect 15016 16940 15068 16992
rect 16028 16983 16080 16992
rect 16028 16949 16037 16983
rect 16037 16949 16071 16983
rect 16071 16949 16080 16983
rect 16028 16940 16080 16949
rect 17040 16940 17092 16992
rect 17868 17221 17877 17255
rect 17877 17221 17911 17255
rect 17911 17221 17920 17255
rect 17868 17212 17920 17221
rect 18880 17212 18932 17264
rect 22192 17212 22244 17264
rect 23112 17255 23164 17264
rect 23112 17221 23121 17255
rect 23121 17221 23155 17255
rect 23155 17221 23164 17255
rect 23112 17212 23164 17221
rect 26148 17212 26200 17264
rect 17408 17076 17460 17128
rect 18236 17076 18288 17128
rect 22284 17144 22336 17196
rect 22652 17076 22704 17128
rect 23020 17187 23072 17196
rect 23020 17153 23029 17187
rect 23029 17153 23063 17187
rect 23063 17153 23072 17187
rect 24124 17187 24176 17196
rect 23020 17144 23072 17153
rect 24124 17153 24133 17187
rect 24133 17153 24167 17187
rect 24167 17153 24176 17187
rect 24124 17144 24176 17153
rect 25504 17144 25556 17196
rect 25872 17144 25924 17196
rect 29644 17212 29696 17264
rect 31484 17144 31536 17196
rect 33048 17144 33100 17196
rect 37096 17144 37148 17196
rect 47032 17212 47084 17264
rect 47124 17212 47176 17264
rect 24032 17076 24084 17128
rect 25136 17076 25188 17128
rect 27068 17076 27120 17128
rect 22468 17008 22520 17060
rect 23204 17008 23256 17060
rect 19156 16940 19208 16992
rect 19248 16940 19300 16992
rect 20996 16940 21048 16992
rect 21916 16940 21968 16992
rect 23940 16940 23992 16992
rect 25596 16940 25648 16992
rect 26792 16940 26844 16992
rect 36176 17076 36228 17128
rect 43904 17119 43956 17128
rect 43904 17085 43913 17119
rect 43913 17085 43947 17119
rect 43947 17085 43956 17119
rect 43904 17076 43956 17085
rect 45376 17119 45428 17128
rect 45376 17085 45385 17119
rect 45385 17085 45419 17119
rect 45419 17085 45428 17119
rect 45376 17076 45428 17085
rect 47216 17144 47268 17196
rect 46756 17076 46808 17128
rect 47676 16983 47728 16992
rect 47676 16949 47685 16983
rect 47685 16949 47719 16983
rect 47719 16949 47728 16983
rect 47676 16940 47728 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 12716 16736 12768 16788
rect 16764 16779 16816 16788
rect 16764 16745 16773 16779
rect 16773 16745 16807 16779
rect 16807 16745 16816 16779
rect 16764 16736 16816 16745
rect 17408 16779 17460 16788
rect 17408 16745 17417 16779
rect 17417 16745 17451 16779
rect 17451 16745 17460 16779
rect 17408 16736 17460 16745
rect 18236 16736 18288 16788
rect 22652 16779 22704 16788
rect 22652 16745 22661 16779
rect 22661 16745 22695 16779
rect 22695 16745 22704 16779
rect 22652 16736 22704 16745
rect 23020 16736 23072 16788
rect 17316 16668 17368 16720
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 14832 16600 14884 16652
rect 15016 16643 15068 16652
rect 15016 16609 15025 16643
rect 15025 16609 15059 16643
rect 15059 16609 15068 16643
rect 15016 16600 15068 16609
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 17040 16600 17092 16652
rect 18328 16600 18380 16652
rect 13360 16532 13412 16584
rect 17132 16532 17184 16584
rect 21916 16668 21968 16720
rect 19248 16600 19300 16652
rect 23204 16668 23256 16720
rect 23940 16736 23992 16788
rect 24032 16736 24084 16788
rect 25504 16736 25556 16788
rect 27068 16779 27120 16788
rect 27068 16745 27077 16779
rect 27077 16745 27111 16779
rect 27111 16745 27120 16779
rect 27068 16736 27120 16745
rect 27620 16779 27672 16788
rect 27620 16745 27629 16779
rect 27629 16745 27663 16779
rect 27663 16745 27672 16779
rect 27620 16736 27672 16745
rect 43904 16779 43956 16788
rect 43904 16745 43913 16779
rect 43913 16745 43947 16779
rect 43947 16745 43956 16779
rect 43904 16736 43956 16745
rect 47216 16736 47268 16788
rect 47860 16736 47912 16788
rect 23388 16668 23440 16720
rect 23756 16600 23808 16652
rect 23940 16600 23992 16652
rect 2136 16464 2188 16516
rect 16028 16464 16080 16516
rect 19984 16464 20036 16516
rect 18144 16396 18196 16448
rect 22284 16464 22336 16516
rect 24860 16532 24912 16584
rect 22192 16396 22244 16448
rect 26976 16600 27028 16652
rect 26792 16575 26844 16584
rect 26792 16541 26801 16575
rect 26801 16541 26835 16575
rect 26835 16541 26844 16575
rect 26792 16532 26844 16541
rect 27896 16532 27948 16584
rect 45652 16600 45704 16652
rect 47768 16600 47820 16652
rect 47676 16464 47728 16516
rect 48136 16507 48188 16516
rect 48136 16473 48145 16507
rect 48145 16473 48179 16507
rect 48179 16473 48188 16507
rect 48136 16464 48188 16473
rect 25412 16396 25464 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 18328 16192 18380 16244
rect 18880 16192 18932 16244
rect 19984 16192 20036 16244
rect 19248 16124 19300 16176
rect 39948 16192 40000 16244
rect 1952 16056 2004 16108
rect 14280 15988 14332 16040
rect 18236 16099 18288 16108
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 18236 16056 18288 16065
rect 18420 16056 18472 16108
rect 19156 16056 19208 16108
rect 22560 16124 22612 16176
rect 24032 16124 24084 16176
rect 21640 16056 21692 16108
rect 22100 16031 22152 16040
rect 22100 15997 22109 16031
rect 22109 15997 22143 16031
rect 22143 15997 22152 16031
rect 44732 16099 44784 16108
rect 44732 16065 44741 16099
rect 44741 16065 44775 16099
rect 44775 16065 44784 16099
rect 44732 16056 44784 16065
rect 47768 16099 47820 16108
rect 47768 16065 47777 16099
rect 47777 16065 47811 16099
rect 47811 16065 47820 16099
rect 47768 16056 47820 16065
rect 22100 15988 22152 15997
rect 45100 15988 45152 16040
rect 46112 16031 46164 16040
rect 46112 15997 46121 16031
rect 46121 15997 46155 16031
rect 46155 15997 46164 16031
rect 46112 15988 46164 15997
rect 17960 15963 18012 15972
rect 15384 15895 15436 15904
rect 15384 15861 15393 15895
rect 15393 15861 15427 15895
rect 15427 15861 15436 15895
rect 15384 15852 15436 15861
rect 17960 15929 17969 15963
rect 17969 15929 18003 15963
rect 18003 15929 18012 15963
rect 17960 15920 18012 15929
rect 24952 15920 25004 15972
rect 25136 15920 25188 15972
rect 20812 15852 20864 15904
rect 22192 15852 22244 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 22100 15648 22152 15700
rect 22560 15648 22612 15700
rect 45100 15691 45152 15700
rect 45100 15657 45109 15691
rect 45109 15657 45143 15691
rect 45143 15657 45152 15691
rect 45100 15648 45152 15657
rect 47492 15648 47544 15700
rect 20536 15580 20588 15632
rect 22284 15580 22336 15632
rect 45560 15580 45612 15632
rect 15384 15555 15436 15564
rect 15384 15521 15393 15555
rect 15393 15521 15427 15555
rect 15427 15521 15436 15555
rect 15384 15512 15436 15521
rect 1768 15444 1820 15496
rect 14280 15487 14332 15496
rect 14280 15453 14289 15487
rect 14289 15453 14323 15487
rect 14323 15453 14332 15487
rect 14280 15444 14332 15453
rect 18420 15487 18472 15496
rect 18420 15453 18429 15487
rect 18429 15453 18463 15487
rect 18463 15453 18472 15487
rect 18420 15444 18472 15453
rect 20996 15487 21048 15496
rect 20996 15453 21005 15487
rect 21005 15453 21039 15487
rect 21039 15453 21048 15487
rect 20996 15444 21048 15453
rect 21640 15487 21692 15496
rect 17040 15419 17092 15428
rect 17040 15385 17049 15419
rect 17049 15385 17083 15419
rect 17083 15385 17092 15419
rect 17040 15376 17092 15385
rect 21640 15453 21649 15487
rect 21649 15453 21683 15487
rect 21683 15453 21692 15487
rect 21640 15444 21692 15453
rect 21916 15376 21968 15428
rect 14372 15351 14424 15360
rect 14372 15317 14381 15351
rect 14381 15317 14415 15351
rect 14415 15317 14424 15351
rect 14372 15308 14424 15317
rect 18512 15351 18564 15360
rect 18512 15317 18521 15351
rect 18521 15317 18555 15351
rect 18555 15317 18564 15351
rect 18512 15308 18564 15317
rect 19984 15308 20036 15360
rect 21824 15351 21876 15360
rect 21824 15317 21833 15351
rect 21833 15317 21867 15351
rect 21867 15317 21876 15351
rect 21824 15308 21876 15317
rect 22836 15444 22888 15496
rect 25780 15444 25832 15496
rect 45652 15444 45704 15496
rect 24400 15308 24452 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 14372 15036 14424 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 16580 14968 16632 15020
rect 18236 14968 18288 15020
rect 21548 15036 21600 15088
rect 21916 15036 21968 15088
rect 23756 15036 23808 15088
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 16856 14943 16908 14952
rect 12440 14832 12492 14884
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 18052 14943 18104 14952
rect 18052 14909 18061 14943
rect 18061 14909 18095 14943
rect 18095 14909 18104 14943
rect 18052 14900 18104 14909
rect 22836 15011 22888 15020
rect 22836 14977 22845 15011
rect 22845 14977 22879 15011
rect 22879 14977 22888 15011
rect 22836 14968 22888 14977
rect 23388 14968 23440 15020
rect 45652 14968 45704 15020
rect 20996 14832 21048 14884
rect 15476 14764 15528 14816
rect 19524 14764 19576 14816
rect 22008 14807 22060 14816
rect 22008 14773 22017 14807
rect 22017 14773 22051 14807
rect 22051 14773 22060 14807
rect 22008 14764 22060 14773
rect 22836 14764 22888 14816
rect 46480 14764 46532 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 20996 14603 21048 14612
rect 15476 14467 15528 14476
rect 15476 14433 15485 14467
rect 15485 14433 15519 14467
rect 15519 14433 15528 14467
rect 15476 14424 15528 14433
rect 18236 14492 18288 14544
rect 20996 14569 21005 14603
rect 21005 14569 21039 14603
rect 21039 14569 21048 14603
rect 20996 14560 21048 14569
rect 21548 14560 21600 14612
rect 23112 14560 23164 14612
rect 22192 14492 22244 14544
rect 18144 14467 18196 14476
rect 18144 14433 18153 14467
rect 18153 14433 18187 14467
rect 18187 14433 18196 14467
rect 18144 14424 18196 14433
rect 19524 14467 19576 14476
rect 19524 14433 19533 14467
rect 19533 14433 19567 14467
rect 19567 14433 19576 14467
rect 19524 14424 19576 14433
rect 2688 14356 2740 14408
rect 14280 14356 14332 14408
rect 18236 14356 18288 14408
rect 21916 14424 21968 14476
rect 23756 14424 23808 14476
rect 17132 14331 17184 14340
rect 17132 14297 17141 14331
rect 17141 14297 17175 14331
rect 17175 14297 17184 14331
rect 17132 14288 17184 14297
rect 22008 14356 22060 14408
rect 19432 14288 19484 14340
rect 19984 14288 20036 14340
rect 20996 14288 21048 14340
rect 15200 14220 15252 14272
rect 21640 14263 21692 14272
rect 21640 14229 21649 14263
rect 21649 14229 21683 14263
rect 21683 14229 21692 14263
rect 21640 14220 21692 14229
rect 24308 14356 24360 14408
rect 32864 14356 32916 14408
rect 45008 14399 45060 14408
rect 45008 14365 45017 14399
rect 45017 14365 45051 14399
rect 45051 14365 45060 14399
rect 45008 14356 45060 14365
rect 25136 14288 25188 14340
rect 45192 14331 45244 14340
rect 45192 14297 45201 14331
rect 45201 14297 45235 14331
rect 45235 14297 45244 14331
rect 45192 14288 45244 14297
rect 46848 14331 46900 14340
rect 46848 14297 46857 14331
rect 46857 14297 46891 14331
rect 46891 14297 46900 14331
rect 46848 14288 46900 14297
rect 30380 14220 30432 14272
rect 30564 14220 30616 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 16856 14016 16908 14068
rect 21548 14016 21600 14068
rect 24308 14059 24360 14068
rect 24308 14025 24317 14059
rect 24317 14025 24351 14059
rect 24351 14025 24360 14059
rect 24308 14016 24360 14025
rect 25136 14016 25188 14068
rect 45192 14059 45244 14068
rect 45192 14025 45201 14059
rect 45201 14025 45235 14059
rect 45235 14025 45244 14059
rect 45192 14016 45244 14025
rect 18144 13948 18196 14000
rect 18512 13948 18564 14000
rect 22836 13948 22888 14000
rect 23388 13948 23440 14000
rect 15660 13880 15712 13932
rect 21824 13923 21876 13932
rect 21824 13889 21833 13923
rect 21833 13889 21867 13923
rect 21867 13889 21876 13923
rect 21824 13880 21876 13889
rect 24400 13880 24452 13932
rect 44180 13880 44232 13932
rect 17960 13812 18012 13864
rect 18236 13812 18288 13864
rect 45008 13812 45060 13864
rect 3424 13744 3476 13796
rect 15936 13744 15988 13796
rect 21824 13676 21876 13728
rect 47768 13719 47820 13728
rect 47768 13685 47777 13719
rect 47777 13685 47811 13719
rect 47811 13685 47820 13719
rect 47768 13676 47820 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 17960 13515 18012 13524
rect 17960 13481 17969 13515
rect 17969 13481 18003 13515
rect 18003 13481 18012 13515
rect 17960 13472 18012 13481
rect 19432 13515 19484 13524
rect 19432 13481 19441 13515
rect 19441 13481 19475 13515
rect 19475 13481 19484 13515
rect 19432 13472 19484 13481
rect 21824 13515 21876 13524
rect 21824 13481 21833 13515
rect 21833 13481 21867 13515
rect 21867 13481 21876 13515
rect 21824 13472 21876 13481
rect 14648 13404 14700 13456
rect 15200 13379 15252 13388
rect 15200 13345 15209 13379
rect 15209 13345 15243 13379
rect 15243 13345 15252 13379
rect 15200 13336 15252 13345
rect 24400 13404 24452 13456
rect 21640 13379 21692 13388
rect 21640 13345 21649 13379
rect 21649 13345 21683 13379
rect 21683 13345 21692 13379
rect 21640 13336 21692 13345
rect 30380 13379 30432 13388
rect 30380 13345 30389 13379
rect 30389 13345 30423 13379
rect 30423 13345 30432 13379
rect 30380 13336 30432 13345
rect 30564 13379 30616 13388
rect 30564 13345 30573 13379
rect 30573 13345 30607 13379
rect 30607 13345 30616 13379
rect 30564 13336 30616 13345
rect 47768 13404 47820 13456
rect 46480 13379 46532 13388
rect 46480 13345 46489 13379
rect 46489 13345 46523 13379
rect 46523 13345 46532 13379
rect 46480 13336 46532 13345
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 32220 13243 32272 13252
rect 32220 13209 32229 13243
rect 32229 13209 32263 13243
rect 32263 13209 32272 13243
rect 32220 13200 32272 13209
rect 48136 13243 48188 13252
rect 48136 13209 48145 13243
rect 48145 13209 48179 13243
rect 48179 13209 48188 13243
rect 48136 13200 48188 13209
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 30472 12588 30524 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 46296 12180 46348 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 22468 11772 22520 11824
rect 22284 11679 22336 11688
rect 22284 11645 22293 11679
rect 22293 11645 22327 11679
rect 22327 11645 22336 11679
rect 22284 11636 22336 11645
rect 23940 11679 23992 11688
rect 23940 11645 23949 11679
rect 23949 11645 23983 11679
rect 23983 11645 23992 11679
rect 23940 11636 23992 11645
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 22284 11339 22336 11348
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 46296 11203 46348 11212
rect 46296 11169 46305 11203
rect 46305 11169 46339 11203
rect 46339 11169 46348 11203
rect 46296 11160 46348 11169
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 38844 11092 38896 11144
rect 46020 11024 46072 11076
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 3148 10956 3200 11008
rect 12440 10956 12492 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 47124 10616 47176 10668
rect 47492 10616 47544 10668
rect 46296 10412 46348 10464
rect 47676 10455 47728 10464
rect 47676 10421 47685 10455
rect 47685 10421 47719 10455
rect 47719 10421 47728 10455
rect 47676 10412 47728 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 47676 10072 47728 10124
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 47860 9571 47912 9580
rect 47860 9537 47869 9571
rect 47869 9537 47903 9571
rect 47903 9537 47912 9571
rect 47860 9528 47912 9537
rect 48228 9392 48280 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 47768 8891 47820 8900
rect 47768 8857 47777 8891
rect 47777 8857 47811 8891
rect 47811 8857 47820 8891
rect 47768 8848 47820 8857
rect 28540 8780 28592 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 46940 8483 46992 8492
rect 46940 8449 46949 8483
rect 46949 8449 46983 8483
rect 46983 8449 46992 8483
rect 46940 8440 46992 8449
rect 47124 8304 47176 8356
rect 3148 8236 3200 8288
rect 18052 8236 18104 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 46756 7896 46808 7948
rect 45468 7803 45520 7812
rect 45468 7769 45477 7803
rect 45477 7769 45511 7803
rect 45511 7769 45520 7803
rect 45468 7760 45520 7769
rect 45560 7803 45612 7812
rect 45560 7769 45569 7803
rect 45569 7769 45603 7803
rect 45603 7769 45612 7803
rect 47032 7803 47084 7812
rect 45560 7760 45612 7769
rect 47032 7769 47041 7803
rect 47041 7769 47075 7803
rect 47075 7769 47084 7803
rect 47032 7760 47084 7769
rect 47124 7803 47176 7812
rect 47124 7769 47133 7803
rect 47133 7769 47167 7803
rect 47167 7769 47176 7803
rect 47124 7760 47176 7769
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 46940 7488 46992 7540
rect 47032 7488 47084 7540
rect 45560 7352 45612 7404
rect 46204 7395 46256 7404
rect 46204 7361 46213 7395
rect 46213 7361 46247 7395
rect 46247 7361 46256 7395
rect 46204 7352 46256 7361
rect 48136 7395 48188 7404
rect 48136 7361 48145 7395
rect 48145 7361 48179 7395
rect 48179 7361 48188 7395
rect 48136 7352 48188 7361
rect 2044 7216 2096 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3424 6808 3476 6860
rect 17132 6808 17184 6860
rect 47308 6851 47360 6860
rect 47308 6817 47317 6851
rect 47317 6817 47351 6851
rect 47351 6817 47360 6851
rect 47308 6808 47360 6817
rect 47216 6740 47268 6792
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 46664 6400 46716 6452
rect 47952 6307 48004 6316
rect 47952 6273 47961 6307
rect 47961 6273 47995 6307
rect 47995 6273 48004 6307
rect 47952 6264 48004 6273
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3976 5720 4028 5772
rect 43168 5763 43220 5772
rect 43168 5729 43177 5763
rect 43177 5729 43211 5763
rect 43211 5729 43220 5763
rect 43168 5720 43220 5729
rect 6644 5652 6696 5704
rect 37280 5627 37332 5636
rect 37280 5593 37289 5627
rect 37289 5593 37323 5627
rect 37323 5593 37332 5627
rect 37280 5584 37332 5593
rect 38476 5584 38528 5636
rect 42248 5627 42300 5636
rect 42248 5593 42257 5627
rect 42257 5593 42291 5627
rect 42291 5593 42300 5627
rect 42248 5584 42300 5593
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 42248 5312 42300 5364
rect 45928 5312 45980 5364
rect 37740 5287 37792 5296
rect 37740 5253 37749 5287
rect 37749 5253 37783 5287
rect 37783 5253 37792 5287
rect 37740 5244 37792 5253
rect 40408 5219 40460 5228
rect 37648 5151 37700 5160
rect 37648 5117 37657 5151
rect 37657 5117 37691 5151
rect 37691 5117 37700 5151
rect 37648 5108 37700 5117
rect 38476 5151 38528 5160
rect 38476 5117 38485 5151
rect 38485 5117 38519 5151
rect 38519 5117 38528 5151
rect 38476 5108 38528 5117
rect 40408 5185 40417 5219
rect 40417 5185 40451 5219
rect 40451 5185 40460 5219
rect 40408 5176 40460 5185
rect 42892 5176 42944 5228
rect 48320 5176 48372 5228
rect 41236 5108 41288 5160
rect 39120 4972 39172 5024
rect 39948 4972 40000 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 37280 4768 37332 4820
rect 40408 4768 40460 4820
rect 41512 4700 41564 4752
rect 39948 4675 40000 4684
rect 39948 4641 39957 4675
rect 39957 4641 39991 4675
rect 39991 4641 40000 4675
rect 39948 4632 40000 4641
rect 41788 4675 41840 4684
rect 41788 4641 41797 4675
rect 41797 4641 41831 4675
rect 41831 4641 41840 4675
rect 41788 4632 41840 4641
rect 45468 4700 45520 4752
rect 46204 4700 46256 4752
rect 43168 4675 43220 4684
rect 43168 4641 43177 4675
rect 43177 4641 43211 4675
rect 43211 4641 43220 4675
rect 43168 4632 43220 4641
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 18052 4564 18104 4616
rect 21916 4564 21968 4616
rect 37280 4607 37332 4616
rect 37280 4573 37289 4607
rect 37289 4573 37323 4607
rect 37323 4573 37332 4607
rect 37280 4564 37332 4573
rect 39120 4607 39172 4616
rect 39120 4573 39129 4607
rect 39129 4573 39163 4607
rect 39163 4573 39172 4607
rect 39120 4564 39172 4573
rect 47400 4632 47452 4684
rect 46848 4564 46900 4616
rect 40132 4539 40184 4548
rect 40132 4505 40141 4539
rect 40141 4505 40175 4539
rect 40175 4505 40184 4539
rect 40132 4496 40184 4505
rect 14188 4428 14240 4480
rect 18236 4428 18288 4480
rect 22376 4428 22428 4480
rect 42524 4428 42576 4480
rect 46480 4428 46532 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 37280 4224 37332 4276
rect 27160 4199 27212 4208
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 2964 3952 3016 4004
rect 11796 4088 11848 4140
rect 12808 4088 12860 4140
rect 12992 4088 13044 4140
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 10416 3952 10468 4004
rect 15016 3952 15068 4004
rect 15568 4088 15620 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 16120 4020 16172 4072
rect 17592 4088 17644 4140
rect 19248 4131 19300 4140
rect 17408 4020 17460 4072
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 20076 4088 20128 4140
rect 20812 4088 20864 4140
rect 18788 4020 18840 4072
rect 27160 4165 27169 4199
rect 27169 4165 27203 4199
rect 27203 4165 27212 4199
rect 27160 4156 27212 4165
rect 22560 4020 22612 4072
rect 22192 3952 22244 4004
rect 25688 4088 25740 4140
rect 24308 4020 24360 4072
rect 31024 4088 31076 4140
rect 28080 4063 28132 4072
rect 28080 4029 28089 4063
rect 28089 4029 28123 4063
rect 28123 4029 28132 4063
rect 28080 4020 28132 4029
rect 31116 4020 31168 4072
rect 31576 4088 31628 4140
rect 37648 4156 37700 4208
rect 40316 4199 40368 4208
rect 37740 4088 37792 4140
rect 38200 4088 38252 4140
rect 40316 4165 40325 4199
rect 40325 4165 40359 4199
rect 40359 4165 40368 4199
rect 40316 4156 40368 4165
rect 46664 4199 46716 4208
rect 46664 4165 46673 4199
rect 46673 4165 46707 4199
rect 46707 4165 46716 4199
rect 46664 4156 46716 4165
rect 47768 4199 47820 4208
rect 47768 4165 47777 4199
rect 47777 4165 47811 4199
rect 47811 4165 47820 4199
rect 47768 4156 47820 4165
rect 39304 4088 39356 4140
rect 40040 4088 40092 4140
rect 36544 4020 36596 4072
rect 41236 4131 41288 4140
rect 41236 4097 41245 4131
rect 41245 4097 41279 4131
rect 41279 4097 41288 4131
rect 41236 4088 41288 4097
rect 42524 4088 42576 4140
rect 42892 4063 42944 4072
rect 42892 4029 42901 4063
rect 42901 4029 42935 4063
rect 42935 4029 42944 4063
rect 42892 4020 42944 4029
rect 28816 3952 28868 4004
rect 1584 3884 1636 3936
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 7380 3884 7432 3936
rect 11244 3884 11296 3936
rect 12072 3884 12124 3936
rect 14556 3884 14608 3936
rect 14740 3884 14792 3936
rect 15292 3927 15344 3936
rect 15292 3893 15301 3927
rect 15301 3893 15335 3927
rect 15335 3893 15344 3927
rect 15292 3884 15344 3893
rect 15384 3884 15436 3936
rect 16028 3884 16080 3936
rect 16856 3884 16908 3936
rect 17500 3884 17552 3936
rect 18696 3927 18748 3936
rect 18696 3893 18705 3927
rect 18705 3893 18739 3927
rect 18739 3893 18748 3927
rect 18696 3884 18748 3893
rect 19340 3927 19392 3936
rect 19340 3893 19349 3927
rect 19349 3893 19383 3927
rect 19383 3893 19392 3927
rect 19340 3884 19392 3893
rect 20536 3884 20588 3936
rect 21824 3884 21876 3936
rect 22836 3927 22888 3936
rect 22836 3893 22845 3927
rect 22845 3893 22879 3927
rect 22879 3893 22888 3927
rect 22836 3884 22888 3893
rect 23388 3884 23440 3936
rect 24860 3927 24912 3936
rect 24860 3893 24869 3927
rect 24869 3893 24903 3927
rect 24903 3893 24912 3927
rect 24860 3884 24912 3893
rect 25596 3927 25648 3936
rect 25596 3893 25605 3927
rect 25605 3893 25639 3927
rect 25639 3893 25648 3927
rect 25596 3884 25648 3893
rect 25964 3884 26016 3936
rect 37372 3927 37424 3936
rect 37372 3893 37381 3927
rect 37381 3893 37415 3927
rect 37415 3893 37424 3927
rect 37372 3884 37424 3893
rect 40224 3884 40276 3936
rect 41420 3884 41472 3936
rect 46296 3884 46348 3936
rect 47860 3927 47912 3936
rect 47860 3893 47869 3927
rect 47869 3893 47903 3927
rect 47903 3893 47912 3927
rect 47860 3884 47912 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3884 3680 3936 3732
rect 44456 3680 44508 3732
rect 6552 3612 6604 3664
rect 1768 3544 1820 3596
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 11520 3587 11572 3596
rect 11520 3553 11529 3587
rect 11529 3553 11563 3587
rect 11563 3553 11572 3587
rect 11520 3544 11572 3553
rect 7196 3476 7248 3528
rect 10416 3519 10468 3528
rect 1308 3408 1360 3460
rect 10416 3485 10425 3519
rect 10425 3485 10459 3519
rect 10459 3485 10468 3519
rect 10416 3476 10468 3485
rect 10968 3476 11020 3528
rect 13636 3476 13688 3528
rect 14280 3612 14332 3664
rect 16672 3612 16724 3664
rect 17408 3655 17460 3664
rect 17408 3621 17417 3655
rect 17417 3621 17451 3655
rect 17451 3621 17460 3655
rect 17408 3612 17460 3621
rect 18052 3655 18104 3664
rect 18052 3621 18061 3655
rect 18061 3621 18095 3655
rect 18095 3621 18104 3655
rect 18052 3612 18104 3621
rect 18144 3612 18196 3664
rect 22652 3612 22704 3664
rect 24308 3612 24360 3664
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 14740 3519 14792 3528
rect 14740 3485 14749 3519
rect 14749 3485 14783 3519
rect 14783 3485 14792 3519
rect 14740 3476 14792 3485
rect 15016 3476 15068 3528
rect 15384 3519 15436 3528
rect 2780 3383 2832 3392
rect 2780 3349 2789 3383
rect 2789 3349 2823 3383
rect 2823 3349 2832 3383
rect 2780 3340 2832 3349
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 8392 3340 8444 3392
rect 10324 3340 10376 3392
rect 10508 3383 10560 3392
rect 10508 3349 10517 3383
rect 10517 3349 10551 3383
rect 10551 3349 10560 3383
rect 10508 3340 10560 3349
rect 10876 3340 10928 3392
rect 11520 3340 11572 3392
rect 13820 3340 13872 3392
rect 14372 3408 14424 3460
rect 15108 3408 15160 3460
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 16028 3519 16080 3528
rect 16028 3485 16037 3519
rect 16037 3485 16071 3519
rect 16071 3485 16080 3519
rect 16028 3476 16080 3485
rect 22284 3544 22336 3596
rect 25596 3612 25648 3664
rect 25688 3612 25740 3664
rect 37004 3612 37056 3664
rect 40132 3612 40184 3664
rect 24860 3587 24912 3596
rect 24860 3553 24869 3587
rect 24869 3553 24903 3587
rect 24903 3553 24912 3587
rect 24860 3544 24912 3553
rect 25136 3587 25188 3596
rect 25136 3553 25145 3587
rect 25145 3553 25179 3587
rect 25179 3553 25188 3587
rect 25136 3544 25188 3553
rect 25228 3544 25280 3596
rect 16856 3476 16908 3528
rect 17500 3476 17552 3528
rect 18696 3476 18748 3528
rect 17592 3408 17644 3460
rect 17776 3408 17828 3460
rect 18788 3408 18840 3460
rect 19524 3519 19576 3528
rect 19524 3485 19533 3519
rect 19533 3485 19567 3519
rect 19567 3485 19576 3519
rect 20260 3519 20312 3528
rect 19524 3476 19576 3485
rect 20260 3485 20269 3519
rect 20269 3485 20303 3519
rect 20303 3485 20312 3519
rect 20260 3476 20312 3485
rect 20536 3476 20588 3528
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 22100 3476 22152 3528
rect 22836 3519 22888 3528
rect 22836 3485 22845 3519
rect 22845 3485 22879 3519
rect 22879 3485 22888 3519
rect 22836 3476 22888 3485
rect 23204 3476 23256 3528
rect 27436 3476 27488 3528
rect 30932 3544 30984 3596
rect 32220 3544 32272 3596
rect 32956 3544 33008 3596
rect 36544 3544 36596 3596
rect 47860 3612 47912 3664
rect 41788 3587 41840 3596
rect 41788 3553 41797 3587
rect 41797 3553 41831 3587
rect 41831 3553 41840 3587
rect 41788 3544 41840 3553
rect 42432 3544 42484 3596
rect 46296 3587 46348 3596
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 31300 3476 31352 3528
rect 26608 3408 26660 3460
rect 26792 3408 26844 3460
rect 38292 3476 38344 3528
rect 40224 3519 40276 3528
rect 40224 3485 40233 3519
rect 40233 3485 40267 3519
rect 40267 3485 40276 3519
rect 40224 3476 40276 3485
rect 41052 3519 41104 3528
rect 41052 3485 41061 3519
rect 41061 3485 41095 3519
rect 41095 3485 41104 3519
rect 41052 3476 41104 3485
rect 45192 3519 45244 3528
rect 25228 3340 25280 3392
rect 26884 3340 26936 3392
rect 31484 3340 31536 3392
rect 33140 3383 33192 3392
rect 33140 3349 33149 3383
rect 33149 3349 33183 3383
rect 33183 3349 33192 3383
rect 33140 3340 33192 3349
rect 39856 3408 39908 3460
rect 41328 3408 41380 3460
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 47492 3408 47544 3460
rect 48964 3408 49016 3460
rect 42340 3340 42392 3392
rect 42616 3340 42668 3392
rect 45376 3340 45428 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2688 3136 2740 3188
rect 12992 3179 13044 3188
rect 2780 3068 2832 3120
rect 7380 3111 7432 3120
rect 7380 3077 7389 3111
rect 7389 3077 7423 3111
rect 7423 3077 7432 3111
rect 7380 3068 7432 3077
rect 12992 3145 13001 3179
rect 13001 3145 13035 3179
rect 13035 3145 13044 3179
rect 12992 3136 13044 3145
rect 13820 3111 13872 3120
rect 13820 3077 13829 3111
rect 13829 3077 13863 3111
rect 13863 3077 13872 3111
rect 13820 3068 13872 3077
rect 14556 3136 14608 3188
rect 17040 3136 17092 3188
rect 18236 3136 18288 3188
rect 19248 3136 19300 3188
rect 17776 3068 17828 3120
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 10968 3000 11020 3009
rect 664 2932 716 2984
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 11980 2975 12032 2984
rect 11980 2941 11989 2975
rect 11989 2941 12023 2975
rect 12023 2941 12032 2975
rect 11980 2932 12032 2941
rect 6460 2864 6512 2916
rect 8208 2864 8260 2916
rect 13636 3043 13688 3052
rect 13636 3009 13645 3043
rect 13645 3009 13679 3043
rect 13679 3009 13688 3043
rect 13636 3000 13688 3009
rect 12808 2932 12860 2984
rect 15108 2975 15160 2984
rect 15108 2941 15117 2975
rect 15117 2941 15151 2975
rect 15151 2941 15160 2975
rect 20536 3136 20588 3188
rect 21916 3179 21968 3188
rect 21916 3145 21925 3179
rect 21925 3145 21959 3179
rect 21959 3145 21968 3179
rect 21916 3136 21968 3145
rect 22560 3179 22612 3188
rect 22560 3145 22569 3179
rect 22569 3145 22603 3179
rect 22603 3145 22612 3179
rect 22560 3136 22612 3145
rect 19524 3111 19576 3120
rect 19524 3077 19533 3111
rect 19533 3077 19567 3111
rect 19567 3077 19576 3111
rect 19524 3068 19576 3077
rect 19708 3068 19760 3120
rect 22928 3068 22980 3120
rect 20720 3000 20772 3052
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 22376 3000 22428 3052
rect 27068 3136 27120 3188
rect 39856 3179 39908 3188
rect 23388 3111 23440 3120
rect 23388 3077 23397 3111
rect 23397 3077 23431 3111
rect 23431 3077 23440 3111
rect 23388 3068 23440 3077
rect 23480 3068 23532 3120
rect 26056 3068 26108 3120
rect 26884 3068 26936 3120
rect 28080 3111 28132 3120
rect 28080 3077 28089 3111
rect 28089 3077 28123 3111
rect 28123 3077 28132 3111
rect 28080 3068 28132 3077
rect 28632 3068 28684 3120
rect 33140 3111 33192 3120
rect 33140 3077 33149 3111
rect 33149 3077 33183 3111
rect 33183 3077 33192 3111
rect 33140 3068 33192 3077
rect 39856 3145 39865 3179
rect 39865 3145 39899 3179
rect 39899 3145 39908 3179
rect 39856 3136 39908 3145
rect 41052 3136 41104 3188
rect 42616 3111 42668 3120
rect 23204 3043 23256 3052
rect 15108 2932 15160 2941
rect 18144 2864 18196 2916
rect 20168 2932 20220 2984
rect 23204 3009 23213 3043
rect 23213 3009 23247 3043
rect 23247 3009 23256 3043
rect 23204 3000 23256 3009
rect 26424 3000 26476 3052
rect 32956 3043 33008 3052
rect 32956 3009 32965 3043
rect 32965 3009 32999 3043
rect 32999 3009 33008 3043
rect 32956 3000 33008 3009
rect 39948 3000 40000 3052
rect 40592 3000 40644 3052
rect 41236 3000 41288 3052
rect 20260 2864 20312 2916
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 10324 2796 10376 2848
rect 22008 2864 22060 2916
rect 22560 2864 22612 2916
rect 23480 2864 23532 2916
rect 27160 2932 27212 2984
rect 32220 2932 32272 2984
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 39304 2932 39356 2984
rect 40684 2975 40736 2984
rect 20536 2796 20588 2848
rect 38384 2864 38436 2916
rect 40040 2864 40092 2916
rect 40684 2941 40693 2975
rect 40693 2941 40727 2975
rect 40727 2941 40736 2975
rect 40684 2932 40736 2941
rect 41512 2864 41564 2916
rect 42616 3077 42625 3111
rect 42625 3077 42659 3111
rect 42659 3077 42668 3111
rect 42616 3068 42668 3077
rect 45376 3111 45428 3120
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 42432 3043 42484 3052
rect 42432 3009 42441 3043
rect 42441 3009 42475 3043
rect 42475 3009 42484 3043
rect 42432 3000 42484 3009
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 46756 3000 46808 3052
rect 43168 2975 43220 2984
rect 43168 2941 43177 2975
rect 43177 2941 43211 2975
rect 43211 2941 43220 2975
rect 43168 2932 43220 2941
rect 47676 2932 47728 2984
rect 30656 2796 30708 2848
rect 38292 2796 38344 2848
rect 41328 2796 41380 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2872 2524 2924 2576
rect 9036 2524 9088 2576
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 6184 2456 6236 2508
rect 6736 2499 6788 2508
rect 6736 2465 6745 2499
rect 6745 2465 6779 2499
rect 6779 2465 6788 2499
rect 6736 2456 6788 2465
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 9772 2456 9824 2508
rect 15200 2592 15252 2644
rect 10048 2524 10100 2576
rect 16764 2456 16816 2508
rect 20076 2592 20128 2644
rect 20444 2592 20496 2644
rect 22100 2592 22152 2644
rect 23480 2592 23532 2644
rect 27436 2635 27488 2644
rect 25044 2567 25096 2576
rect 25044 2533 25053 2567
rect 25053 2533 25087 2567
rect 25087 2533 25096 2567
rect 25044 2524 25096 2533
rect 27436 2601 27445 2635
rect 27445 2601 27479 2635
rect 27479 2601 27488 2635
rect 27436 2592 27488 2601
rect 35348 2592 35400 2644
rect 35900 2592 35952 2644
rect 40316 2635 40368 2644
rect 40316 2601 40325 2635
rect 40325 2601 40359 2635
rect 40359 2601 40368 2635
rect 40316 2592 40368 2601
rect 40592 2635 40644 2644
rect 40592 2601 40601 2635
rect 40601 2601 40635 2635
rect 40635 2601 40644 2635
rect 40592 2592 40644 2601
rect 48044 2635 48096 2644
rect 48044 2601 48053 2635
rect 48053 2601 48087 2635
rect 48087 2601 48096 2635
rect 48044 2592 48096 2601
rect 23940 2456 23992 2508
rect 27988 2456 28040 2508
rect 32680 2456 32732 2508
rect 35900 2456 35952 2508
rect 41880 2524 41932 2576
rect 2596 2320 2648 2372
rect 5172 2388 5224 2440
rect 14188 2431 14240 2440
rect 14188 2397 14197 2431
rect 14197 2397 14231 2431
rect 14231 2397 14240 2431
rect 14188 2388 14240 2397
rect 15292 2388 15344 2440
rect 16120 2388 16172 2440
rect 19340 2388 19392 2440
rect 23204 2388 23256 2440
rect 26976 2431 27028 2440
rect 26976 2397 26985 2431
rect 26985 2397 27019 2431
rect 27019 2397 27028 2431
rect 26976 2388 27028 2397
rect 28356 2388 28408 2440
rect 29644 2388 29696 2440
rect 35440 2388 35492 2440
rect 10508 2320 10560 2372
rect 15476 2320 15528 2372
rect 20628 2320 20680 2372
rect 21916 2320 21968 2372
rect 24492 2320 24544 2372
rect 27068 2320 27120 2372
rect 11980 2252 12032 2304
rect 15568 2252 15620 2304
rect 15752 2295 15804 2304
rect 15752 2261 15761 2295
rect 15761 2261 15795 2295
rect 15795 2261 15804 2295
rect 15752 2252 15804 2261
rect 21732 2252 21784 2304
rect 27344 2252 27396 2304
rect 29736 2295 29788 2304
rect 29736 2261 29745 2295
rect 29745 2261 29779 2295
rect 29779 2261 29788 2295
rect 29736 2252 29788 2261
rect 32496 2252 32548 2304
rect 40684 2456 40736 2508
rect 42524 2456 42576 2508
rect 38016 2388 38068 2440
rect 38200 2388 38252 2440
rect 40040 2431 40092 2440
rect 36084 2320 36136 2372
rect 39304 2320 39356 2372
rect 40040 2397 40049 2431
rect 40049 2397 40083 2431
rect 40083 2397 40092 2431
rect 40040 2388 40092 2397
rect 40592 2388 40644 2440
rect 43812 2388 43864 2440
rect 47032 2388 47084 2440
rect 46388 2320 46440 2372
rect 48044 2320 48096 2372
rect 45468 2295 45520 2304
rect 45468 2261 45477 2295
rect 45477 2261 45511 2295
rect 45511 2261 45520 2295
rect 45468 2252 45520 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 4068 2048 4120 2100
rect 10048 2048 10100 2100
rect 21180 1980 21232 2032
rect 45468 1980 45520 2032
rect 15752 1912 15804 1964
rect 37372 1912 37424 1964
rect 29736 1844 29788 1896
rect 41420 1844 41472 1896
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4752 49314
rect 4498 49200 4610 49286
rect 32 19922 60 49200
rect 1858 47696 1914 47705
rect 1858 47631 1914 47640
rect 1872 46646 1900 47631
rect 1964 47054 1992 49200
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2044 46980 2096 46986
rect 2044 46922 2096 46928
rect 1860 46640 1912 46646
rect 1860 46582 1912 46588
rect 1768 45960 1820 45966
rect 1768 45902 1820 45908
rect 1780 45490 1808 45902
rect 1768 45484 1820 45490
rect 1768 45426 1820 45432
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1676 43240 1728 43246
rect 1676 43182 1728 43188
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1584 41540 1636 41546
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1596 35465 1624 35634
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1584 33992 1636 33998
rect 1584 33934 1636 33940
rect 1400 33448 1452 33454
rect 1398 33416 1400 33425
rect 1452 33416 1454 33425
rect 1398 33351 1454 33360
rect 1596 32745 1624 33934
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 1400 32224 1452 32230
rect 1400 32166 1452 32172
rect 1412 31890 1440 32166
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1688 26234 1716 43182
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 1872 40225 1900 40394
rect 1952 40384 2004 40390
rect 1952 40326 2004 40332
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1780 36786 1808 37198
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1964 34066 1992 40326
rect 1952 34060 2004 34066
rect 1952 34002 2004 34008
rect 1952 33856 2004 33862
rect 1952 33798 2004 33804
rect 1860 33448 1912 33454
rect 1860 33390 1912 33396
rect 1872 32910 1900 33390
rect 1964 33114 1992 33798
rect 1952 33108 2004 33114
rect 1952 33050 2004 33056
rect 1860 32904 1912 32910
rect 1860 32846 1912 32852
rect 1872 31414 1900 32846
rect 1860 31408 1912 31414
rect 1860 31350 1912 31356
rect 1596 26206 1716 26234
rect 2056 26234 2084 46922
rect 2608 46918 2636 49200
rect 3252 47054 3280 49200
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3422 47016 3478 47025
rect 3422 46951 3478 46960
rect 2596 46912 2648 46918
rect 2596 46854 2648 46860
rect 2136 46368 2188 46374
rect 2136 46310 2188 46316
rect 2778 46336 2834 46345
rect 2148 35894 2176 46310
rect 2778 46271 2834 46280
rect 2792 45422 2820 46271
rect 2320 45416 2372 45422
rect 2320 45358 2372 45364
rect 2780 45416 2832 45422
rect 2780 45358 2832 45364
rect 2332 45082 2360 45358
rect 2320 45076 2372 45082
rect 2320 45018 2372 45024
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36718 2820 36751
rect 2228 36712 2280 36718
rect 2228 36654 2280 36660
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 2240 36378 2268 36654
rect 2228 36372 2280 36378
rect 2228 36314 2280 36320
rect 2412 36168 2464 36174
rect 2412 36110 2464 36116
rect 2148 35866 2268 35894
rect 2136 35488 2188 35494
rect 2136 35430 2188 35436
rect 2148 32434 2176 35430
rect 2136 32428 2188 32434
rect 2136 32370 2188 32376
rect 2240 27606 2268 35866
rect 2320 32768 2372 32774
rect 2320 32710 2372 32716
rect 2332 32502 2360 32710
rect 2320 32496 2372 32502
rect 2320 32438 2372 32444
rect 2228 27600 2280 27606
rect 2228 27542 2280 27548
rect 2424 26234 2452 36110
rect 3238 32056 3294 32065
rect 3238 31991 3294 32000
rect 3252 31822 3280 31991
rect 3240 31816 3292 31822
rect 3240 31758 3292 31764
rect 2596 31272 2648 31278
rect 2596 31214 2648 31220
rect 2056 26206 2176 26234
rect 20 19916 72 19922
rect 20 19858 72 19864
rect 1596 18834 1624 26206
rect 1858 25256 1914 25265
rect 1858 25191 1860 25200
rect 1912 25191 1914 25200
rect 1860 25162 1912 25168
rect 2044 25152 2096 25158
rect 2044 25094 2096 25100
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 23225 1900 23666
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 1584 18624 1636 18630
rect 1584 18566 1636 18572
rect 1596 18426 1624 18566
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17785 1440 18226
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1872 16425 1900 16594
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1964 6914 1992 16050
rect 2056 7274 2084 25094
rect 2148 23254 2176 26206
rect 2332 26206 2452 26234
rect 2136 23248 2188 23254
rect 2136 23190 2188 23196
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2332 18766 2360 26206
rect 2608 21146 2636 31214
rect 3330 28656 3386 28665
rect 3330 28591 3386 28600
rect 3344 27674 3372 28591
rect 3332 27668 3384 27674
rect 3332 27610 3384 27616
rect 2596 21140 2648 21146
rect 2596 21082 2648 21088
rect 3436 21010 3464 46951
rect 3896 46646 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4724 47054 4752 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49314 7186 50000
rect 7074 49286 7328 49314
rect 7074 49200 7186 49286
rect 5828 47054 5856 49200
rect 7300 47054 7328 49286
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49314 13626 50000
rect 13514 49286 13768 49314
rect 13514 49200 13626 49286
rect 4712 47048 4764 47054
rect 4712 46990 4764 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7288 47048 7340 47054
rect 7288 46990 7340 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 4988 46980 5040 46986
rect 4988 46922 5040 46928
rect 6644 46980 6696 46986
rect 6644 46922 6696 46928
rect 3884 46640 3936 46646
rect 3884 46582 3936 46588
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 3988 46170 4016 46446
rect 3976 46164 4028 46170
rect 3976 46106 4028 46112
rect 3514 44976 3570 44985
rect 3514 44911 3570 44920
rect 3424 21004 3476 21010
rect 3424 20946 3476 20952
rect 3528 20602 3556 44911
rect 3792 44872 3844 44878
rect 3792 44814 3844 44820
rect 3698 43616 3754 43625
rect 3698 43551 3754 43560
rect 3606 31376 3662 31385
rect 3606 31311 3662 31320
rect 3620 23866 3648 31311
rect 3712 26234 3740 43551
rect 3804 31822 3832 44814
rect 3882 39536 3938 39545
rect 3882 39471 3938 39480
rect 3792 31816 3844 31822
rect 3792 31758 3844 31764
rect 3712 26206 3832 26234
rect 3608 23860 3660 23866
rect 3608 23802 3660 23808
rect 3804 21486 3832 26206
rect 3896 22710 3924 39471
rect 3976 31816 4028 31822
rect 3976 31758 4028 31764
rect 3884 22704 3936 22710
rect 3884 22646 3936 22652
rect 3792 21480 3844 21486
rect 3792 21422 3844 21428
rect 3988 21078 4016 31758
rect 3976 21072 4028 21078
rect 3976 21014 4028 21020
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3516 20324 3568 20330
rect 3516 20266 3568 20272
rect 3528 19825 3556 20266
rect 3514 19816 3570 19825
rect 3514 19751 3570 19760
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 3436 18465 3464 19110
rect 3422 18456 3478 18465
rect 3422 18391 3478 18400
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3068 17105 3096 17818
rect 3054 17096 3110 17105
rect 3054 17031 3110 17040
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 2148 16250 2176 16458
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 1964 6886 2084 6914
rect 2056 4146 2084 6886
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1320 800 1348 3402
rect 1596 2514 1624 3878
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 3058 1808 3538
rect 2700 3534 2728 14350
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3436 13705 3464 13738
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10305 3188 10950
rect 3146 10296 3202 10305
rect 3146 10231 3202 10240
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 7585 3188 8230
rect 3146 7576 3202 7585
rect 3146 7511 3202 7520
rect 4080 6914 4108 46922
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4620 32360 4672 32366
rect 4620 32302 4672 32308
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4632 31278 4660 32302
rect 4620 31272 4672 31278
rect 4620 31214 4672 31220
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4632 18426 4660 31214
rect 5000 20058 5028 46922
rect 5172 46504 5224 46510
rect 5172 46446 5224 46452
rect 5184 46170 5212 46446
rect 5172 46164 5224 46170
rect 5172 46106 5224 46112
rect 6552 31136 6604 31142
rect 6552 31078 6604 31084
rect 6564 30802 6592 31078
rect 6552 30796 6604 30802
rect 6552 30738 6604 30744
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3422 6896 3478 6905
rect 3422 6831 3424 6840
rect 3476 6831 3478 6840
rect 3988 6886 4108 6914
rect 3424 6802 3476 6808
rect 3988 5778 4016 6886
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2700 3194 2728 3470
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2792 3126 2820 3334
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2884 2582 2912 3878
rect 2976 3505 3004 3946
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 2962 3496 3018 3505
rect 2962 3431 3018 3440
rect 2872 2576 2924 2582
rect 2872 2518 2924 2524
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2608 800 2636 2314
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 2792 785 2820 2450
rect 3896 800 3924 3674
rect 6564 3670 6592 18702
rect 6656 5710 6684 46922
rect 7472 46912 7524 46918
rect 7472 46854 7524 46860
rect 7484 28626 7512 46854
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9496 46980 9548 46986
rect 9496 46922 9548 46928
rect 8312 45526 8432 45554
rect 7564 31680 7616 31686
rect 7564 31622 7616 31628
rect 7576 30802 7604 31622
rect 7564 30796 7616 30802
rect 7564 30738 7616 30744
rect 8208 30796 8260 30802
rect 8208 30738 8260 30744
rect 7472 28620 7524 28626
rect 7472 28562 7524 28568
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 6196 2514 6224 3470
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4080 1465 4108 2042
rect 4066 1456 4122 1465
rect 4066 1391 4122 1400
rect 5184 800 5212 2382
rect 6472 800 6500 2858
rect 6748 2514 6776 3334
rect 7208 3058 7236 3470
rect 7392 3126 7420 3878
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7116 800 7144 2450
rect 7760 800 7788 2926
rect 8220 2922 8248 30738
rect 8312 25362 8340 45526
rect 9508 38418 9536 46922
rect 10980 46374 11008 49200
rect 10968 46368 11020 46374
rect 10968 46310 11020 46316
rect 11624 46034 11652 49200
rect 12268 47122 12296 49200
rect 12256 47116 12308 47122
rect 12256 47058 12308 47064
rect 12912 46918 12940 49200
rect 13740 47138 13768 49286
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49314 16202 50000
rect 16090 49286 16528 49314
rect 16090 49200 16202 49286
rect 14200 47954 14228 49200
rect 14200 47926 14320 47954
rect 13740 47110 14228 47138
rect 14200 47054 14228 47110
rect 14188 47048 14240 47054
rect 14188 46990 14240 46996
rect 12900 46912 12952 46918
rect 12900 46854 12952 46860
rect 14292 46510 14320 47926
rect 15016 46980 15068 46986
rect 15016 46922 15068 46928
rect 11888 46504 11940 46510
rect 11888 46446 11940 46452
rect 13544 46504 13596 46510
rect 13544 46446 13596 46452
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 11612 46028 11664 46034
rect 11612 45970 11664 45976
rect 11900 45626 11928 46446
rect 13556 46170 13584 46446
rect 14200 46170 14228 46446
rect 13544 46164 13596 46170
rect 13544 46106 13596 46112
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 11980 45960 12032 45966
rect 11980 45902 12032 45908
rect 14096 45960 14148 45966
rect 14096 45902 14148 45908
rect 11888 45620 11940 45626
rect 11888 45562 11940 45568
rect 9496 38412 9548 38418
rect 9496 38354 9548 38360
rect 11992 36106 12020 45902
rect 14108 41138 14136 45902
rect 14096 41132 14148 41138
rect 14096 41074 14148 41080
rect 11980 36100 12032 36106
rect 11980 36042 12032 36048
rect 15028 27538 15056 46922
rect 15488 45554 15516 49200
rect 16500 47054 16528 49286
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49314 27150 50000
rect 26712 49286 27150 49314
rect 17420 47410 17448 49200
rect 16960 47382 17448 47410
rect 18604 47456 18656 47462
rect 18604 47398 18656 47404
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 15488 45526 16160 45554
rect 15936 35692 15988 35698
rect 15936 35634 15988 35640
rect 15948 34610 15976 35634
rect 15936 34604 15988 34610
rect 15936 34546 15988 34552
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 15016 27532 15068 27538
rect 15016 27474 15068 27480
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 12440 27056 12492 27062
rect 12440 26998 12492 27004
rect 11244 26920 11296 26926
rect 11244 26862 11296 26868
rect 11520 26920 11572 26926
rect 11520 26862 11572 26868
rect 12348 26920 12400 26926
rect 12348 26862 12400 26868
rect 11256 26586 11284 26862
rect 11244 26580 11296 26586
rect 11244 26522 11296 26528
rect 11532 26042 11560 26862
rect 11520 26036 11572 26042
rect 11520 25978 11572 25984
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 8300 25356 8352 25362
rect 8300 25298 8352 25304
rect 9128 25220 9180 25226
rect 9128 25162 9180 25168
rect 9140 24954 9168 25162
rect 9128 24948 9180 24954
rect 9128 24890 9180 24896
rect 10704 24818 10732 25842
rect 11796 25764 11848 25770
rect 11796 25706 11848 25712
rect 11808 25498 11836 25706
rect 11796 25492 11848 25498
rect 11796 25434 11848 25440
rect 11612 25424 11664 25430
rect 11612 25366 11664 25372
rect 11624 25158 11652 25366
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11520 25152 11572 25158
rect 11520 25094 11572 25100
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 11532 24954 11560 25094
rect 11520 24948 11572 24954
rect 11520 24890 11572 24896
rect 8944 24812 8996 24818
rect 8944 24754 8996 24760
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 8588 23322 8616 23598
rect 8576 23316 8628 23322
rect 8576 23258 8628 23264
rect 8956 23118 8984 24754
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 10324 24608 10376 24614
rect 10324 24550 10376 24556
rect 9692 24342 9720 24550
rect 9680 24336 9732 24342
rect 9680 24278 9732 24284
rect 10336 24274 10364 24550
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8680 22234 8708 22510
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8956 22030 8984 23054
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 9784 17882 9812 23598
rect 10704 23118 10732 24754
rect 10784 24404 10836 24410
rect 10784 24346 10836 24352
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10796 22098 10824 24346
rect 11624 24342 11652 24754
rect 11716 24750 11744 25230
rect 11808 24886 11836 25434
rect 12360 25294 12388 26862
rect 12452 26042 12480 26998
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12072 25220 12124 25226
rect 12072 25162 12124 25168
rect 11796 24880 11848 24886
rect 11796 24822 11848 24828
rect 12084 24818 12112 25162
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 11704 24744 11756 24750
rect 11704 24686 11756 24692
rect 11612 24336 11664 24342
rect 11612 24278 11664 24284
rect 12084 24070 12112 24754
rect 12452 24206 12480 25842
rect 12544 24818 12572 26250
rect 12636 25430 12664 26386
rect 13004 26382 13032 27406
rect 14464 27396 14516 27402
rect 14464 27338 14516 27344
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 13280 27130 13308 27270
rect 14476 27130 14504 27338
rect 13268 27124 13320 27130
rect 13268 27066 13320 27072
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 12624 25424 12676 25430
rect 12624 25366 12676 25372
rect 12728 25158 12756 26318
rect 14004 25900 14056 25906
rect 14004 25842 14056 25848
rect 13176 25832 13228 25838
rect 13176 25774 13228 25780
rect 13452 25832 13504 25838
rect 13452 25774 13504 25780
rect 12808 25696 12860 25702
rect 12808 25638 12860 25644
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12728 24954 12756 25094
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 12084 23798 12112 24006
rect 12072 23792 12124 23798
rect 12072 23734 12124 23740
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11520 22976 11572 22982
rect 11520 22918 11572 22924
rect 11532 22642 11560 22918
rect 11520 22636 11572 22642
rect 11520 22578 11572 22584
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10796 21570 10824 22034
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 10796 21554 10916 21570
rect 11532 21554 11560 21830
rect 11716 21690 11744 23054
rect 12728 22778 12756 24890
rect 12820 24886 12848 25638
rect 13188 25226 13216 25774
rect 13360 25424 13412 25430
rect 13360 25366 13412 25372
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 12808 24880 12860 24886
rect 12808 24822 12860 24828
rect 13188 24750 13216 25162
rect 13176 24744 13228 24750
rect 13176 24686 13228 24692
rect 13372 24614 13400 25366
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13372 24206 13400 24550
rect 13464 24410 13492 25774
rect 14016 25158 14044 25842
rect 14188 25288 14240 25294
rect 14188 25230 14240 25236
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 13556 24954 13584 25094
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13556 24206 13584 24890
rect 13728 24268 13780 24274
rect 13728 24210 13780 24216
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13740 23594 13768 24210
rect 13728 23588 13780 23594
rect 13728 23530 13780 23536
rect 13740 23186 13768 23530
rect 13728 23180 13780 23186
rect 13728 23122 13780 23128
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12072 22704 12124 22710
rect 12072 22646 12124 22652
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11808 22098 11836 22510
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 10796 21548 10928 21554
rect 10796 21542 10876 21548
rect 10876 21490 10928 21496
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10428 21146 10456 21354
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10324 21072 10376 21078
rect 10322 21040 10324 21049
rect 10376 21040 10378 21049
rect 10322 20975 10378 20984
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 10428 20602 10456 20878
rect 10704 20874 10732 21286
rect 10692 20868 10744 20874
rect 10692 20810 10744 20816
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 11072 19854 11100 20198
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 11532 19378 11560 21490
rect 11716 20466 11744 21626
rect 12084 21146 12112 22646
rect 12452 22098 12480 22646
rect 12440 22092 12492 22098
rect 12728 22094 12756 22714
rect 13176 22228 13228 22234
rect 13176 22170 13228 22176
rect 12440 22034 12492 22040
rect 12544 22066 12756 22094
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12268 21554 12296 21966
rect 12544 21962 12572 22066
rect 13188 22030 13216 22170
rect 14016 22098 14044 25094
rect 14200 24954 14228 25230
rect 14188 24948 14240 24954
rect 14188 24890 14240 24896
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 14200 24410 14228 24754
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14200 22114 14228 23666
rect 14292 22234 14320 26930
rect 15120 26518 15148 27610
rect 16132 27538 16160 45526
rect 16672 36712 16724 36718
rect 16672 36654 16724 36660
rect 16684 36582 16712 36654
rect 16672 36576 16724 36582
rect 16672 36518 16724 36524
rect 16580 34536 16632 34542
rect 16580 34478 16632 34484
rect 16592 33930 16620 34478
rect 16684 34066 16712 36518
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 16764 34944 16816 34950
rect 16764 34886 16816 34892
rect 16672 34060 16724 34066
rect 16672 34002 16724 34008
rect 16580 33924 16632 33930
rect 16580 33866 16632 33872
rect 16776 33862 16804 34886
rect 16868 34746 16896 35022
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 16764 33856 16816 33862
rect 16764 33798 16816 33804
rect 16672 33516 16724 33522
rect 16672 33458 16724 33464
rect 16684 33114 16712 33458
rect 16672 33108 16724 33114
rect 16672 33050 16724 33056
rect 16684 32434 16712 33050
rect 16672 32428 16724 32434
rect 16672 32370 16724 32376
rect 16580 31340 16632 31346
rect 16684 31328 16712 32370
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16764 31340 16816 31346
rect 16684 31300 16764 31328
rect 16580 31282 16632 31288
rect 16764 31282 16816 31288
rect 16592 30938 16620 31282
rect 16580 30932 16632 30938
rect 16580 30874 16632 30880
rect 16868 30258 16896 31826
rect 16960 31754 16988 47382
rect 17224 47252 17276 47258
rect 17224 47194 17276 47200
rect 17236 37874 17264 47194
rect 18144 38480 18196 38486
rect 18144 38422 18196 38428
rect 17224 37868 17276 37874
rect 17224 37810 17276 37816
rect 18156 37670 18184 38422
rect 18144 37664 18196 37670
rect 18144 37606 18196 37612
rect 17960 36848 18012 36854
rect 17960 36790 18012 36796
rect 17500 36236 17552 36242
rect 17500 36178 17552 36184
rect 17040 35080 17092 35086
rect 17040 35022 17092 35028
rect 17052 33658 17080 35022
rect 17316 34536 17368 34542
rect 17316 34478 17368 34484
rect 17328 33862 17356 34478
rect 17316 33856 17368 33862
rect 17316 33798 17368 33804
rect 17040 33652 17092 33658
rect 17040 33594 17092 33600
rect 17224 33584 17276 33590
rect 17224 33526 17276 33532
rect 17040 33448 17092 33454
rect 17040 33390 17092 33396
rect 17052 32978 17080 33390
rect 17236 33318 17264 33526
rect 17328 33454 17356 33798
rect 17512 33522 17540 36178
rect 17972 35834 18000 36790
rect 17960 35828 18012 35834
rect 17960 35770 18012 35776
rect 17592 34536 17644 34542
rect 17592 34478 17644 34484
rect 17500 33516 17552 33522
rect 17500 33458 17552 33464
rect 17316 33448 17368 33454
rect 17316 33390 17368 33396
rect 17224 33312 17276 33318
rect 17224 33254 17276 33260
rect 17040 32972 17092 32978
rect 17040 32914 17092 32920
rect 17236 32910 17264 33254
rect 17512 33114 17540 33458
rect 17500 33108 17552 33114
rect 17500 33050 17552 33056
rect 17224 32904 17276 32910
rect 17224 32846 17276 32852
rect 17236 32366 17264 32846
rect 17224 32360 17276 32366
rect 17224 32302 17276 32308
rect 17224 32224 17276 32230
rect 17224 32166 17276 32172
rect 17316 32224 17368 32230
rect 17316 32166 17368 32172
rect 16960 31726 17080 31754
rect 16856 30252 16908 30258
rect 16856 30194 16908 30200
rect 16868 29238 16896 30194
rect 16856 29232 16908 29238
rect 16856 29174 16908 29180
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16684 28082 16712 29106
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 17052 27538 17080 31726
rect 17132 31680 17184 31686
rect 17132 31622 17184 31628
rect 17144 31482 17172 31622
rect 17132 31476 17184 31482
rect 17132 31418 17184 31424
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 16120 27532 16172 27538
rect 16120 27474 16172 27480
rect 16856 27532 16908 27538
rect 16856 27474 16908 27480
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 16868 27402 16896 27474
rect 16764 27396 16816 27402
rect 16764 27338 16816 27344
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16776 27130 16804 27338
rect 16764 27124 16816 27130
rect 16764 27066 16816 27072
rect 17144 26874 17172 31282
rect 17236 31142 17264 32166
rect 17328 32026 17356 32166
rect 17316 32020 17368 32026
rect 17316 31962 17368 31968
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 17408 27056 17460 27062
rect 17408 26998 17460 27004
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 16960 26846 17172 26874
rect 15200 26784 15252 26790
rect 15200 26726 15252 26732
rect 15108 26512 15160 26518
rect 15108 26454 15160 26460
rect 15212 26450 15240 26726
rect 15200 26444 15252 26450
rect 15200 26386 15252 26392
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14752 25770 14780 26318
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 14740 25764 14792 25770
rect 14740 25706 14792 25712
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14476 25362 14504 25638
rect 14464 25356 14516 25362
rect 14464 25298 14516 25304
rect 14752 24818 14780 25706
rect 15108 25696 15160 25702
rect 15108 25638 15160 25644
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 15120 25226 15148 25638
rect 15108 25220 15160 25226
rect 15108 25162 15160 25168
rect 15948 24818 15976 25638
rect 16500 25430 16528 26250
rect 16856 26036 16908 26042
rect 16856 25978 16908 25984
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 16776 25498 16804 25842
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16488 25424 16540 25430
rect 16488 25366 16540 25372
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 16500 25158 16528 25230
rect 16396 25152 16448 25158
rect 16396 25094 16448 25100
rect 16488 25152 16540 25158
rect 16488 25094 16540 25100
rect 16408 24818 16436 25094
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 14752 23118 14780 24754
rect 16028 24608 16080 24614
rect 16028 24550 16080 24556
rect 16040 24342 16068 24550
rect 16028 24336 16080 24342
rect 16028 24278 16080 24284
rect 16408 24138 16436 24754
rect 16396 24132 16448 24138
rect 16396 24074 16448 24080
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14384 22642 14412 22918
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14372 22160 14424 22166
rect 14200 22108 14372 22114
rect 14200 22102 14424 22108
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 14200 22086 14412 22102
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 13280 21894 13308 21966
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13740 21622 13768 22034
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 12256 21548 12308 21554
rect 12308 21508 12480 21536
rect 12256 21490 12308 21496
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 12084 20942 12112 21082
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 12360 20874 12388 21286
rect 12348 20868 12400 20874
rect 12348 20810 12400 20816
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11624 19786 11652 20198
rect 12452 19836 12480 21508
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 12636 21146 12664 21422
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12820 20466 12848 20742
rect 12912 20602 12940 20878
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 13556 20466 13584 21422
rect 13740 21146 13768 21422
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 14004 21004 14056 21010
rect 14004 20946 14056 20952
rect 14016 20913 14044 20946
rect 14200 20942 14228 22086
rect 14476 21418 14504 22170
rect 14752 22094 14780 23054
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15396 22710 15424 22918
rect 15384 22704 15436 22710
rect 15384 22646 15436 22652
rect 14660 22066 14780 22094
rect 14660 21894 14688 22066
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 14372 21072 14424 21078
rect 14370 21040 14372 21049
rect 14424 21040 14426 21049
rect 14370 20975 14426 20984
rect 14188 20936 14240 20942
rect 14002 20904 14058 20913
rect 14188 20878 14240 20884
rect 14002 20839 14058 20848
rect 14188 20800 14240 20806
rect 14372 20800 14424 20806
rect 14240 20760 14372 20788
rect 14188 20742 14240 20748
rect 14372 20742 14424 20748
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 12820 20369 12848 20402
rect 12806 20360 12862 20369
rect 12806 20295 12862 20304
rect 12900 20324 12952 20330
rect 12900 20266 12952 20272
rect 12624 19848 12676 19854
rect 12452 19808 12624 19836
rect 12624 19790 12676 19796
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 12912 19446 12940 20266
rect 13556 20058 13584 20402
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13556 19786 13584 19994
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 12900 19440 12952 19446
rect 12900 19382 12952 19388
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12820 18766 12848 19110
rect 13832 18766 13860 19790
rect 13924 19174 13952 20538
rect 14476 20466 14504 21354
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14462 20360 14518 20369
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14200 19786 14228 20198
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14292 19718 14320 20198
rect 14384 20058 14412 20334
rect 14462 20295 14518 20304
rect 14476 20058 14504 20295
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14280 19712 14332 19718
rect 14200 19660 14280 19666
rect 14200 19654 14332 19660
rect 14200 19638 14320 19654
rect 14200 19378 14228 19638
rect 14384 19446 14412 19994
rect 14568 19854 14596 20878
rect 14832 20528 14884 20534
rect 14832 20470 14884 20476
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14844 19378 14872 20470
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 12820 17678 12848 18702
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13096 18290 13124 18566
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13832 17678 13860 18702
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 18358 14136 18566
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12636 17270 12664 17478
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12820 17134 12848 17614
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 17270 13492 17478
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12728 16794 12756 17070
rect 14200 16998 14228 19314
rect 14752 19258 14780 19314
rect 14752 19230 14872 19258
rect 14844 19174 14872 19230
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14752 18222 14780 18566
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14844 17678 14872 19110
rect 14936 18766 14964 19450
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 15028 18766 15056 19382
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15028 18222 15056 18702
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 13372 16590 13400 16934
rect 14844 16658 14872 17614
rect 15396 17610 15424 19790
rect 15580 18834 15608 20198
rect 15764 19922 15792 20198
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 16658 15056 16934
rect 15304 16658 15332 17478
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13372 15026 13400 16526
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14292 15502 14320 15982
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15396 15570 15424 15846
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12452 11014 12480 14826
rect 14292 14414 14320 15438
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14384 15094 14412 15302
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15488 14482 15516 14758
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14660 12434 14688 13398
rect 15212 13394 15240 14214
rect 15672 13938 15700 14962
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15948 13802 15976 21898
rect 16408 21554 16436 21966
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 16500 21146 16528 25094
rect 16776 24954 16804 25434
rect 16764 24948 16816 24954
rect 16764 24890 16816 24896
rect 16868 24818 16896 25978
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 16684 23798 16712 24142
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 16672 23792 16724 23798
rect 16672 23734 16724 23740
rect 16776 23662 16804 24006
rect 16868 23730 16896 24210
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16592 23118 16620 23598
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 16592 22574 16620 23054
rect 16776 22778 16804 23122
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16212 21140 16264 21146
rect 16212 21082 16264 21088
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16224 20058 16252 21082
rect 16592 20942 16620 21830
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16868 21146 16896 21286
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16592 20466 16620 20878
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16040 16522 16068 16934
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 16592 15026 16620 20402
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 16794 16804 17614
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16868 17270 16896 17478
rect 16856 17264 16908 17270
rect 16856 17206 16908 17212
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16868 14074 16896 14894
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 14660 12406 14872 12434
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10428 3534 10456 3946
rect 11244 3936 11296 3942
rect 11808 3924 11836 4082
rect 12072 3936 12124 3942
rect 11808 3896 12072 3924
rect 11244 3878 11296 3884
rect 12072 3878 12124 3884
rect 11256 3602 11284 3878
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 8404 800 8432 3334
rect 10336 2854 10364 3334
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 9048 800 9076 2518
rect 9784 2514 9812 2790
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 10060 2106 10088 2518
rect 10520 2378 10548 3334
rect 10888 2774 10916 3334
rect 10980 3058 11008 3470
rect 11532 3398 11560 3538
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 12820 2990 12848 4082
rect 13004 3194 13032 4082
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13648 3058 13676 3470
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13832 3126 13860 3334
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 10888 2746 11008 2774
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 10048 2100 10100 2106
rect 10048 2042 10100 2048
rect 10980 800 11008 2746
rect 11992 2310 12020 2926
rect 14200 2446 14228 4422
rect 14292 3670 14320 4558
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14280 3664 14332 3670
rect 14280 3606 14332 3612
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14384 2774 14412 3402
rect 14568 3194 14596 3878
rect 14752 3534 14780 3878
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14292 2746 14412 2774
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 14292 1578 14320 2746
rect 14200 1550 14320 1578
rect 14200 800 14228 1550
rect 14844 800 14872 12406
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 15028 3534 15056 3946
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15108 3460 15160 3466
rect 15108 3402 15160 3408
rect 15120 2990 15148 3402
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 15212 2650 15240 4082
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15304 2446 15332 3878
rect 15396 3534 15424 3878
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15488 800 15516 2314
rect 15580 2310 15608 4082
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16040 3534 16068 3878
rect 16132 3602 16160 4014
rect 16684 3670 16712 4082
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16868 3534 16896 3878
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16960 2774 16988 26846
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 17052 24138 17080 24754
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 17040 24132 17092 24138
rect 17040 24074 17092 24080
rect 17144 23730 17172 24550
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17144 23254 17172 23666
rect 17132 23248 17184 23254
rect 17132 23190 17184 23196
rect 17236 22094 17264 26930
rect 17052 22066 17264 22094
rect 17052 21894 17080 22066
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 17420 20942 17448 26998
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 17052 20262 17080 20742
rect 17316 20528 17368 20534
rect 17316 20470 17368 20476
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17052 17882 17080 20198
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17236 18358 17264 19246
rect 17224 18352 17276 18358
rect 17224 18294 17276 18300
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 17144 17134 17172 18226
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17052 16658 17080 16934
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17144 16590 17172 17070
rect 17328 16726 17356 20470
rect 17420 20466 17448 20878
rect 17512 20534 17540 25094
rect 17500 20528 17552 20534
rect 17500 20470 17552 20476
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17604 18834 17632 34478
rect 17776 33108 17828 33114
rect 17776 33050 17828 33056
rect 17788 32434 17816 33050
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17684 32292 17736 32298
rect 17684 32234 17736 32240
rect 17696 31890 17724 32234
rect 17788 31958 17816 32370
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 18064 31958 18092 32302
rect 17776 31952 17828 31958
rect 17776 31894 17828 31900
rect 18052 31952 18104 31958
rect 18052 31894 18104 31900
rect 17684 31884 17736 31890
rect 17684 31826 17736 31832
rect 17868 31748 17920 31754
rect 17868 31690 17920 31696
rect 17880 31482 17908 31690
rect 17868 31476 17920 31482
rect 17868 31418 17920 31424
rect 17960 30320 18012 30326
rect 17960 30262 18012 30268
rect 17972 29850 18000 30262
rect 17960 29844 18012 29850
rect 17960 29786 18012 29792
rect 18156 29646 18184 37606
rect 18616 37466 18644 47398
rect 18708 46918 18736 49200
rect 19248 47116 19300 47122
rect 19248 47058 19300 47064
rect 18696 46912 18748 46918
rect 18696 46854 18748 46860
rect 19064 38752 19116 38758
rect 19064 38694 19116 38700
rect 18604 37460 18656 37466
rect 18604 37402 18656 37408
rect 18328 37256 18380 37262
rect 18328 37198 18380 37204
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18236 36712 18288 36718
rect 18236 36654 18288 36660
rect 18248 36242 18276 36654
rect 18236 36236 18288 36242
rect 18236 36178 18288 36184
rect 18340 36038 18368 37198
rect 18604 37188 18656 37194
rect 18604 37130 18656 37136
rect 18512 37120 18564 37126
rect 18512 37062 18564 37068
rect 18524 36174 18552 37062
rect 18616 36582 18644 37130
rect 18604 36576 18656 36582
rect 18604 36518 18656 36524
rect 18616 36242 18644 36518
rect 18604 36236 18656 36242
rect 18604 36178 18656 36184
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 18328 36032 18380 36038
rect 18328 35974 18380 35980
rect 18340 34746 18368 35974
rect 18328 34740 18380 34746
rect 18328 34682 18380 34688
rect 18420 34536 18472 34542
rect 18420 34478 18472 34484
rect 18432 34066 18460 34478
rect 18420 34060 18472 34066
rect 18420 34002 18472 34008
rect 18420 32972 18472 32978
rect 18420 32914 18472 32920
rect 18236 32768 18288 32774
rect 18236 32710 18288 32716
rect 18248 31872 18276 32710
rect 18432 32008 18460 32914
rect 18616 32842 18644 36178
rect 18708 35834 18736 37198
rect 18696 35828 18748 35834
rect 18696 35770 18748 35776
rect 18708 34678 18736 35770
rect 18696 34672 18748 34678
rect 18696 34614 18748 34620
rect 18604 32836 18656 32842
rect 18604 32778 18656 32784
rect 18972 32428 19024 32434
rect 18972 32370 19024 32376
rect 18696 32224 18748 32230
rect 18696 32166 18748 32172
rect 18708 32026 18736 32166
rect 18696 32020 18748 32026
rect 18432 31980 18644 32008
rect 18328 31884 18380 31890
rect 18248 31844 18328 31872
rect 18328 31826 18380 31832
rect 18616 31822 18644 31980
rect 18696 31962 18748 31968
rect 18696 31884 18748 31890
rect 18696 31826 18748 31832
rect 18604 31816 18656 31822
rect 18604 31758 18656 31764
rect 18604 31680 18656 31686
rect 18708 31668 18736 31826
rect 18984 31822 19012 32370
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 18656 31640 18736 31668
rect 18604 31622 18656 31628
rect 18880 31408 18932 31414
rect 18880 31350 18932 31356
rect 18892 30666 18920 31350
rect 18880 30660 18932 30666
rect 18880 30602 18932 30608
rect 19076 30258 19104 38694
rect 19260 38350 19288 47058
rect 19996 46918 20024 49200
rect 20168 47048 20220 47054
rect 20168 46990 20220 46996
rect 19984 46912 20036 46918
rect 19984 46854 20036 46860
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19892 46504 19944 46510
rect 19892 46446 19944 46452
rect 19904 46170 19932 46446
rect 19892 46164 19944 46170
rect 19892 46106 19944 46112
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19248 38344 19300 38350
rect 19248 38286 19300 38292
rect 19340 38208 19392 38214
rect 19340 38150 19392 38156
rect 19352 37126 19380 38150
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19800 37936 19852 37942
rect 19800 37878 19852 37884
rect 19432 37800 19484 37806
rect 19432 37742 19484 37748
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 19444 36718 19472 37742
rect 19812 37466 19840 37878
rect 19800 37460 19852 37466
rect 19800 37402 19852 37408
rect 20180 37398 20208 46990
rect 20536 46980 20588 46986
rect 20536 46922 20588 46928
rect 20260 45960 20312 45966
rect 20260 45902 20312 45908
rect 20168 37392 20220 37398
rect 20168 37334 20220 37340
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19432 36712 19484 36718
rect 19432 36654 19484 36660
rect 19800 36712 19852 36718
rect 19800 36654 19852 36660
rect 19812 36378 19840 36654
rect 19800 36372 19852 36378
rect 19800 36314 19852 36320
rect 19432 36168 19484 36174
rect 19432 36110 19484 36116
rect 19340 35692 19392 35698
rect 19340 35634 19392 35640
rect 19352 35086 19380 35634
rect 19444 35154 19472 36110
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19432 35148 19484 35154
rect 19432 35090 19484 35096
rect 20168 35148 20220 35154
rect 20168 35090 20220 35096
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 19432 34944 19484 34950
rect 19432 34886 19484 34892
rect 19444 34678 19472 34886
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19432 34672 19484 34678
rect 19432 34614 19484 34620
rect 19984 34400 20036 34406
rect 19984 34342 20036 34348
rect 19996 34202 20024 34342
rect 19984 34196 20036 34202
rect 19984 34138 20036 34144
rect 19340 34060 19392 34066
rect 19340 34002 19392 34008
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19260 33658 19288 33934
rect 19248 33652 19300 33658
rect 19248 33594 19300 33600
rect 19352 33386 19380 34002
rect 20076 33924 20128 33930
rect 20076 33866 20128 33872
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19524 33516 19576 33522
rect 19524 33458 19576 33464
rect 19536 33425 19564 33458
rect 19522 33416 19578 33425
rect 19340 33380 19392 33386
rect 19522 33351 19578 33360
rect 19340 33322 19392 33328
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19984 32904 20036 32910
rect 19984 32846 20036 32852
rect 19260 32366 19288 32846
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19352 32434 19380 32710
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19996 32434 20024 32846
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19248 32360 19300 32366
rect 19248 32302 19300 32308
rect 19260 31278 19288 32302
rect 19340 32224 19392 32230
rect 19340 32166 19392 32172
rect 19352 31414 19380 32166
rect 19432 31748 19484 31754
rect 19432 31690 19484 31696
rect 19444 31482 19472 31690
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 19340 31408 19392 31414
rect 19340 31350 19392 31356
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19248 31272 19300 31278
rect 19444 31249 19472 31282
rect 19984 31272 20036 31278
rect 19248 31214 19300 31220
rect 19430 31240 19486 31249
rect 20088 31249 20116 33866
rect 19984 31214 20036 31220
rect 20074 31240 20130 31249
rect 19430 31175 19486 31184
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19444 30258 19472 30330
rect 19064 30252 19116 30258
rect 19064 30194 19116 30200
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 19800 30252 19852 30258
rect 19800 30194 19852 30200
rect 19524 30184 19576 30190
rect 19524 30126 19576 30132
rect 19536 29850 19564 30126
rect 19812 30054 19840 30194
rect 19800 30048 19852 30054
rect 19800 29990 19852 29996
rect 19996 30002 20024 31214
rect 20074 31175 20130 31184
rect 20088 30190 20116 31175
rect 20180 30394 20208 35090
rect 20168 30388 20220 30394
rect 20168 30330 20220 30336
rect 20076 30184 20128 30190
rect 20076 30126 20128 30132
rect 19524 29844 19576 29850
rect 19524 29786 19576 29792
rect 19524 29708 19576 29714
rect 19524 29650 19576 29656
rect 18144 29640 18196 29646
rect 19536 29594 19564 29650
rect 19812 29646 19840 29990
rect 19996 29974 20208 30002
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 18144 29582 18196 29588
rect 18156 29186 18184 29582
rect 19444 29566 19564 29594
rect 19800 29640 19852 29646
rect 19800 29582 19852 29588
rect 18156 29170 18276 29186
rect 18156 29164 18288 29170
rect 18156 29158 18236 29164
rect 18156 28558 18184 29158
rect 18236 29106 18288 29112
rect 19444 29034 19472 29566
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19996 29306 20024 29786
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 19984 29300 20036 29306
rect 19984 29242 20036 29248
rect 20088 29170 20116 29582
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 19432 29028 19484 29034
rect 19432 28970 19484 28976
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 18328 28484 18380 28490
rect 18328 28426 18380 28432
rect 18512 28484 18564 28490
rect 18512 28426 18564 28432
rect 17776 28416 17828 28422
rect 17776 28358 17828 28364
rect 17788 28150 17816 28358
rect 17776 28144 17828 28150
rect 17776 28086 17828 28092
rect 18340 27878 18368 28426
rect 18524 28218 18552 28426
rect 19352 28218 19380 28494
rect 19444 28422 19472 28970
rect 19904 28626 19932 29106
rect 20088 28762 20116 29106
rect 20076 28756 20128 28762
rect 20076 28698 20128 28704
rect 19892 28620 19944 28626
rect 19892 28562 19944 28568
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 18512 28212 18564 28218
rect 18512 28154 18564 28160
rect 19340 28212 19392 28218
rect 19340 28154 19392 28160
rect 18328 27872 18380 27878
rect 18328 27814 18380 27820
rect 19248 27872 19300 27878
rect 19248 27814 19300 27820
rect 19260 27470 19288 27814
rect 19352 27470 19380 28154
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19248 27464 19300 27470
rect 19248 27406 19300 27412
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19352 26994 19380 27270
rect 19444 27130 19472 28086
rect 19524 28076 19576 28082
rect 19524 28018 19576 28024
rect 19536 27674 19564 28018
rect 19524 27668 19576 27674
rect 19524 27610 19576 27616
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19996 26994 20024 28358
rect 20180 27690 20208 29974
rect 20088 27662 20208 27690
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 17960 26920 18012 26926
rect 17960 26862 18012 26868
rect 17972 25498 18000 26862
rect 19984 26784 20036 26790
rect 19984 26726 20036 26732
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19996 25906 20024 26726
rect 18236 25900 18288 25906
rect 18236 25842 18288 25848
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18052 25696 18104 25702
rect 18052 25638 18104 25644
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17868 25152 17920 25158
rect 17868 25094 17920 25100
rect 17880 24206 17908 25094
rect 18064 24818 18092 25638
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17880 23798 17908 24006
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18064 23254 18092 23598
rect 18052 23248 18104 23254
rect 18052 23190 18104 23196
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17776 22568 17828 22574
rect 17776 22510 17828 22516
rect 17788 22234 17816 22510
rect 17776 22228 17828 22234
rect 17776 22170 17828 22176
rect 17880 22166 17908 22986
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17696 21622 17724 21966
rect 17684 21616 17736 21622
rect 17684 21558 17736 21564
rect 17880 19854 17908 22102
rect 18156 22094 18184 25774
rect 18248 25498 18276 25842
rect 18420 25696 18472 25702
rect 18420 25638 18472 25644
rect 18236 25492 18288 25498
rect 18236 25434 18288 25440
rect 18432 24886 18460 25638
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18420 24880 18472 24886
rect 18420 24822 18472 24828
rect 18524 24342 18552 25230
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 19352 24954 19380 25162
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 19524 24676 19576 24682
rect 19524 24618 19576 24624
rect 18512 24336 18564 24342
rect 18512 24278 18564 24284
rect 19536 24206 19564 24618
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19444 23730 19472 24006
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19904 23118 19932 23666
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19996 22681 20024 25842
rect 20088 23526 20116 27662
rect 20272 27554 20300 45902
rect 20548 45554 20576 46922
rect 20640 46510 20668 49200
rect 20812 47252 20864 47258
rect 20812 47194 20864 47200
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 20548 45526 20668 45554
rect 20352 39500 20404 39506
rect 20352 39442 20404 39448
rect 20364 38962 20392 39442
rect 20352 38956 20404 38962
rect 20352 38898 20404 38904
rect 20364 35086 20392 38898
rect 20536 38888 20588 38894
rect 20536 38830 20588 38836
rect 20548 37806 20576 38830
rect 20536 37800 20588 37806
rect 20536 37742 20588 37748
rect 20536 35556 20588 35562
rect 20536 35498 20588 35504
rect 20352 35080 20404 35086
rect 20352 35022 20404 35028
rect 20364 29714 20392 35022
rect 20548 34950 20576 35498
rect 20536 34944 20588 34950
rect 20536 34886 20588 34892
rect 20548 33998 20576 34886
rect 20536 33992 20588 33998
rect 20536 33934 20588 33940
rect 20548 31346 20576 33934
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 20352 29708 20404 29714
rect 20352 29650 20404 29656
rect 20536 29504 20588 29510
rect 20536 29446 20588 29452
rect 20548 29170 20576 29446
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20352 27668 20404 27674
rect 20352 27610 20404 27616
rect 20180 27526 20300 27554
rect 20180 23798 20208 27526
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20272 27130 20300 27406
rect 20260 27124 20312 27130
rect 20260 27066 20312 27072
rect 20272 26450 20300 27066
rect 20364 26586 20392 27610
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 20260 26444 20312 26450
rect 20260 26386 20312 26392
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20260 24200 20312 24206
rect 20260 24142 20312 24148
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20272 23662 20300 24142
rect 20260 23656 20312 23662
rect 20260 23598 20312 23604
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20076 23248 20128 23254
rect 20076 23190 20128 23196
rect 19982 22672 20038 22681
rect 19982 22607 20038 22616
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 17972 22066 18184 22094
rect 17972 20806 18000 22066
rect 18144 21412 18196 21418
rect 18144 21354 18196 21360
rect 18156 20942 18184 21354
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 18418 20904 18474 20913
rect 18418 20839 18474 20848
rect 18432 20806 18460 20839
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17788 18970 17816 19246
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17420 16794 17448 17070
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17040 15428 17092 15434
rect 17040 15370 17092 15376
rect 17052 3194 17080 15370
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 17144 6866 17172 14282
rect 17512 12434 17540 18634
rect 18064 18290 18092 18770
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17604 17610 17632 17818
rect 17776 17808 17828 17814
rect 17776 17750 17828 17756
rect 17788 17610 17816 17750
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17880 17270 17908 18022
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17972 15978 18000 18226
rect 18064 17338 18092 18226
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18156 16454 18184 20742
rect 18340 20534 18368 20742
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18236 20324 18288 20330
rect 18236 20266 18288 20272
rect 18248 19310 18276 20266
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 18248 18766 18276 19246
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18248 17814 18276 18702
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 18236 17808 18288 17814
rect 18236 17750 18288 17756
rect 18340 17678 18368 17818
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 17134 18276 17478
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18248 16794 18276 17070
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18248 16114 18276 16730
rect 18340 16658 18368 17614
rect 18880 17264 18932 17270
rect 18880 17206 18932 17212
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18340 16250 18368 16594
rect 18892 16250 18920 17206
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 18248 15026 18276 16050
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17972 13530 18000 13806
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17512 12406 17724 12434
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17420 3670 17448 4014
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17512 3534 17540 3878
rect 17500 3528 17552 3534
rect 17406 3496 17462 3505
rect 17500 3470 17552 3476
rect 17604 3466 17632 4082
rect 17406 3431 17462 3440
rect 17592 3460 17644 3466
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16776 2746 16988 2774
rect 16776 2514 16804 2746
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15764 1970 15792 2246
rect 15752 1964 15804 1970
rect 15752 1906 15804 1912
rect 16132 800 16160 2382
rect 17420 800 17448 3431
rect 17592 3402 17644 3408
rect 17696 3097 17724 12406
rect 18064 8294 18092 14894
rect 18248 14550 18276 14962
rect 18236 14544 18288 14550
rect 18236 14486 18288 14492
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18156 14006 18184 14418
rect 18236 14408 18288 14414
rect 18340 14362 18368 16186
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18432 15502 18460 16050
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18288 14356 18368 14362
rect 18236 14350 18368 14356
rect 18248 14334 18368 14350
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18248 13870 18276 14334
rect 18524 14006 18552 15302
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18064 3670 18092 4558
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17788 3126 17816 3402
rect 17776 3120 17828 3126
rect 17682 3088 17738 3097
rect 17776 3062 17828 3068
rect 17682 3023 17738 3032
rect 18156 2922 18184 3606
rect 18248 3194 18276 4422
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18708 3534 18736 3878
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18800 3466 18828 4014
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 18708 870 18920 898
rect 18708 800 18736 870
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 18892 762 18920 870
rect 19076 762 19104 22510
rect 19996 22234 20024 22607
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19984 22092 20036 22098
rect 19984 22034 20036 22040
rect 19260 20942 19288 22034
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19352 21350 19380 21966
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19444 21554 19472 21830
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19996 21622 20024 22034
rect 20088 21962 20116 23190
rect 20076 21956 20128 21962
rect 20076 21898 20128 21904
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19352 19854 19380 21286
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19984 20528 20036 20534
rect 19982 20496 19984 20505
rect 20036 20496 20038 20505
rect 19982 20431 20038 20440
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 19168 19378 19196 19654
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19168 16998 19196 19314
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19260 16998 19288 17546
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19168 16114 19196 16934
rect 19260 16658 19288 16934
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 16182 19288 16594
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19996 16250 20024 16458
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19536 14482 19564 14758
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19996 14346 20024 15302
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19444 13530 19472 14282
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 20364 12434 20392 26318
rect 20536 24744 20588 24750
rect 20536 24686 20588 24692
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20456 24274 20484 24550
rect 20444 24268 20496 24274
rect 20444 24210 20496 24216
rect 20548 23254 20576 24686
rect 20536 23248 20588 23254
rect 20536 23190 20588 23196
rect 20444 22024 20496 22030
rect 20444 21966 20496 21972
rect 20456 21690 20484 21966
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20456 21010 20484 21626
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 20456 19514 20484 19722
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20548 15638 20576 17614
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20364 12406 20484 12434
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19260 3194 19288 4082
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19352 2446 19380 3878
rect 19524 3528 19576 3534
rect 19444 3488 19524 3516
rect 19444 3074 19472 3488
rect 19524 3470 19576 3476
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19524 3120 19576 3126
rect 19444 3068 19524 3074
rect 19444 3062 19576 3068
rect 19708 3120 19760 3126
rect 19708 3062 19760 3068
rect 19444 3046 19564 3062
rect 19720 2774 19748 3062
rect 19982 2952 20038 2961
rect 19982 2887 20038 2896
rect 19628 2746 19748 2774
rect 19340 2440 19392 2446
rect 19628 2428 19656 2746
rect 19340 2382 19392 2388
rect 19444 2400 19656 2428
rect 19444 2258 19472 2400
rect 19352 2230 19472 2258
rect 19352 800 19380 2230
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2887
rect 20088 2650 20116 4082
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20166 3088 20222 3097
rect 20166 3023 20222 3032
rect 20180 2990 20208 3023
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20272 2922 20300 3470
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20456 2650 20484 12406
rect 20640 4049 20668 45526
rect 20824 39030 20852 47194
rect 20996 47048 21048 47054
rect 20996 46990 21048 46996
rect 21008 46034 21036 46990
rect 21284 46034 21312 49200
rect 22560 47456 22612 47462
rect 22560 47398 22612 47404
rect 22572 47258 22600 47398
rect 22560 47252 22612 47258
rect 22560 47194 22612 47200
rect 22008 47048 22060 47054
rect 22008 46990 22060 46996
rect 24860 47048 24912 47054
rect 24860 46990 24912 46996
rect 22020 46646 22048 46990
rect 24872 46646 24900 46990
rect 22008 46640 22060 46646
rect 22008 46582 22060 46588
rect 24860 46640 24912 46646
rect 24860 46582 24912 46588
rect 25148 46510 25176 49200
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 25136 46504 25188 46510
rect 25136 46446 25188 46452
rect 24780 46170 24808 46446
rect 24768 46164 24820 46170
rect 24768 46106 24820 46112
rect 25792 46034 25820 49200
rect 20996 46028 21048 46034
rect 20996 45970 21048 45976
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 25780 46028 25832 46034
rect 25780 45970 25832 45976
rect 25228 45960 25280 45966
rect 25228 45902 25280 45908
rect 20996 45892 21048 45898
rect 20996 45834 21048 45840
rect 21008 45626 21036 45834
rect 24492 45824 24544 45830
rect 24492 45766 24544 45772
rect 20996 45620 21048 45626
rect 20996 45562 21048 45568
rect 20904 45484 20956 45490
rect 20904 45426 20956 45432
rect 20916 41414 20944 45426
rect 20916 41386 21680 41414
rect 20812 39024 20864 39030
rect 20812 38966 20864 38972
rect 21364 38548 21416 38554
rect 21364 38490 21416 38496
rect 20812 38208 20864 38214
rect 20812 38150 20864 38156
rect 20824 37942 20852 38150
rect 20812 37936 20864 37942
rect 20812 37878 20864 37884
rect 21180 37664 21232 37670
rect 21180 37606 21232 37612
rect 21192 37330 21220 37606
rect 21376 37398 21404 38490
rect 21364 37392 21416 37398
rect 21364 37334 21416 37340
rect 21180 37324 21232 37330
rect 21180 37266 21232 37272
rect 20996 37256 21048 37262
rect 20996 37198 21048 37204
rect 20812 35012 20864 35018
rect 20812 34954 20864 34960
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20732 33522 20760 34342
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20824 33402 20852 34954
rect 20904 34604 20956 34610
rect 20904 34546 20956 34552
rect 20916 34066 20944 34546
rect 21008 34134 21036 37198
rect 21272 36576 21324 36582
rect 21272 36518 21324 36524
rect 21088 36168 21140 36174
rect 21088 36110 21140 36116
rect 21100 34746 21128 36110
rect 21284 35766 21312 36518
rect 21456 36168 21508 36174
rect 21456 36110 21508 36116
rect 21272 35760 21324 35766
rect 21272 35702 21324 35708
rect 21284 35086 21312 35702
rect 21272 35080 21324 35086
rect 21272 35022 21324 35028
rect 21088 34740 21140 34746
rect 21088 34682 21140 34688
rect 21284 34542 21312 35022
rect 21468 35018 21496 36110
rect 21456 35012 21508 35018
rect 21456 34954 21508 34960
rect 21272 34536 21324 34542
rect 21272 34478 21324 34484
rect 20996 34128 21048 34134
rect 20996 34070 21048 34076
rect 20904 34060 20956 34066
rect 20904 34002 20956 34008
rect 20916 33590 20944 34002
rect 21088 33992 21140 33998
rect 21088 33934 21140 33940
rect 20904 33584 20956 33590
rect 20904 33526 20956 33532
rect 20824 33374 20944 33402
rect 20720 33312 20772 33318
rect 20720 33254 20772 33260
rect 20732 32298 20760 33254
rect 20812 32768 20864 32774
rect 20812 32710 20864 32716
rect 20720 32292 20772 32298
rect 20720 32234 20772 32240
rect 20732 29646 20760 32234
rect 20824 31822 20852 32710
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 20916 31210 20944 33374
rect 20904 31204 20956 31210
rect 20904 31146 20956 31152
rect 20996 31136 21048 31142
rect 20996 31078 21048 31084
rect 20904 30932 20956 30938
rect 20904 30874 20956 30880
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20732 28694 20760 29582
rect 20812 29572 20864 29578
rect 20812 29514 20864 29520
rect 20720 28688 20772 28694
rect 20720 28630 20772 28636
rect 20720 28416 20772 28422
rect 20720 28358 20772 28364
rect 20732 28150 20760 28358
rect 20720 28144 20772 28150
rect 20720 28086 20772 28092
rect 20732 27690 20760 28086
rect 20824 27878 20852 29514
rect 20916 29306 20944 30874
rect 21008 30802 21036 31078
rect 20996 30796 21048 30802
rect 20996 30738 21048 30744
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 21008 29073 21036 30738
rect 20994 29064 21050 29073
rect 20994 28999 21050 29008
rect 21008 28014 21036 28999
rect 21100 28558 21128 33934
rect 21284 33522 21312 34478
rect 21456 34400 21508 34406
rect 21456 34342 21508 34348
rect 21468 34202 21496 34342
rect 21456 34196 21508 34202
rect 21456 34138 21508 34144
rect 21364 33992 21416 33998
rect 21364 33934 21416 33940
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 21376 33318 21404 33934
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21272 32836 21324 32842
rect 21272 32778 21324 32784
rect 21284 32570 21312 32778
rect 21272 32564 21324 32570
rect 21272 32506 21324 32512
rect 21180 32360 21232 32366
rect 21180 32302 21232 32308
rect 21192 31958 21220 32302
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21180 31952 21232 31958
rect 21180 31894 21232 31900
rect 21376 31754 21404 32166
rect 21376 31726 21496 31754
rect 21272 31680 21324 31686
rect 21272 31622 21324 31628
rect 21284 30734 21312 31622
rect 21468 31482 21496 31726
rect 21456 31476 21508 31482
rect 21456 31418 21508 31424
rect 21468 30734 21496 31418
rect 21652 30870 21680 41386
rect 22100 39296 22152 39302
rect 22100 39238 22152 39244
rect 22112 39030 22140 39238
rect 22100 39024 22152 39030
rect 22100 38966 22152 38972
rect 22560 39024 22612 39030
rect 22560 38966 22612 38972
rect 22572 38554 22600 38966
rect 24124 38888 24176 38894
rect 24124 38830 24176 38836
rect 22560 38548 22612 38554
rect 22560 38490 22612 38496
rect 22836 38344 22888 38350
rect 22836 38286 22888 38292
rect 22376 38004 22428 38010
rect 22376 37946 22428 37952
rect 22388 37670 22416 37946
rect 22744 37800 22796 37806
rect 22744 37742 22796 37748
rect 22192 37664 22244 37670
rect 22192 37606 22244 37612
rect 22376 37664 22428 37670
rect 22376 37606 22428 37612
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 21928 36854 21956 37198
rect 21732 36848 21784 36854
rect 21732 36790 21784 36796
rect 21916 36848 21968 36854
rect 21916 36790 21968 36796
rect 21744 36378 21772 36790
rect 21732 36372 21784 36378
rect 21732 36314 21784 36320
rect 21824 35692 21876 35698
rect 21824 35634 21876 35640
rect 21836 35290 21864 35634
rect 21824 35284 21876 35290
rect 21824 35226 21876 35232
rect 21640 30864 21692 30870
rect 21640 30806 21692 30812
rect 21272 30728 21324 30734
rect 21272 30670 21324 30676
rect 21456 30728 21508 30734
rect 21732 30728 21784 30734
rect 21456 30670 21508 30676
rect 21652 30676 21732 30682
rect 21652 30670 21784 30676
rect 21652 30654 21772 30670
rect 21180 29096 21232 29102
rect 21180 29038 21232 29044
rect 21088 28552 21140 28558
rect 21088 28494 21140 28500
rect 21100 28150 21128 28494
rect 21088 28144 21140 28150
rect 21088 28086 21140 28092
rect 20996 28008 21048 28014
rect 20996 27950 21048 27956
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 21088 27872 21140 27878
rect 21088 27814 21140 27820
rect 20732 27674 20852 27690
rect 20720 27668 20852 27674
rect 20772 27662 20852 27668
rect 20720 27610 20772 27616
rect 20720 27532 20772 27538
rect 20720 27474 20772 27480
rect 20732 26994 20760 27474
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20824 26790 20852 27662
rect 21100 27402 21128 27814
rect 20996 27396 21048 27402
rect 20996 27338 21048 27344
rect 21088 27396 21140 27402
rect 21088 27338 21140 27344
rect 21008 26858 21036 27338
rect 20996 26852 21048 26858
rect 20996 26794 21048 26800
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 21100 26518 21128 27338
rect 21088 26512 21140 26518
rect 21088 26454 21140 26460
rect 20812 23792 20864 23798
rect 20812 23734 20864 23740
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18834 20760 19110
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20824 15910 20852 23734
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 21100 21622 21128 21830
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 21008 15502 21036 16934
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 21008 14618 21036 14826
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 21008 14346 21036 14554
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20626 4040 20682 4049
rect 20626 3975 20682 3984
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20548 3534 20576 3878
rect 20824 3534 20852 4082
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20548 2854 20576 3130
rect 20720 3052 20772 3058
rect 20640 3012 20720 3040
rect 20640 2961 20668 3012
rect 20720 2994 20772 3000
rect 20626 2952 20682 2961
rect 20626 2887 20682 2896
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20640 800 20668 2314
rect 21192 2038 21220 29038
rect 21456 28416 21508 28422
rect 21456 28358 21508 28364
rect 21272 28144 21324 28150
rect 21272 28086 21324 28092
rect 21284 27946 21312 28086
rect 21272 27940 21324 27946
rect 21272 27882 21324 27888
rect 21284 26994 21312 27882
rect 21468 27674 21496 28358
rect 21456 27668 21508 27674
rect 21456 27610 21508 27616
rect 21364 27328 21416 27334
rect 21364 27270 21416 27276
rect 21376 26994 21404 27270
rect 21468 27062 21496 27610
rect 21456 27056 21508 27062
rect 21456 26998 21508 27004
rect 21272 26988 21324 26994
rect 21272 26930 21324 26936
rect 21364 26988 21416 26994
rect 21364 26930 21416 26936
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21468 21350 21496 22578
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21560 21010 21588 21286
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21468 19854 21496 20878
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21652 17252 21680 30654
rect 21732 29300 21784 29306
rect 21732 29242 21784 29248
rect 21744 28082 21772 29242
rect 21928 29238 21956 36790
rect 22008 35624 22060 35630
rect 22008 35566 22060 35572
rect 22020 31822 22048 35566
rect 22100 35148 22152 35154
rect 22100 35090 22152 35096
rect 22112 34678 22140 35090
rect 22100 34672 22152 34678
rect 22100 34614 22152 34620
rect 22204 34610 22232 37606
rect 22756 37466 22784 37742
rect 22848 37670 22876 38286
rect 23204 38276 23256 38282
rect 23204 38218 23256 38224
rect 22836 37664 22888 37670
rect 22836 37606 22888 37612
rect 22744 37460 22796 37466
rect 22744 37402 22796 37408
rect 22560 37188 22612 37194
rect 22560 37130 22612 37136
rect 22572 36038 22600 37130
rect 22652 36236 22704 36242
rect 22652 36178 22704 36184
rect 22560 36032 22612 36038
rect 22560 35974 22612 35980
rect 22572 35034 22600 35974
rect 22664 35834 22692 36178
rect 22652 35828 22704 35834
rect 22652 35770 22704 35776
rect 22572 35006 22692 35034
rect 22376 34944 22428 34950
rect 22376 34886 22428 34892
rect 22388 34610 22416 34886
rect 22192 34604 22244 34610
rect 22192 34546 22244 34552
rect 22376 34604 22428 34610
rect 22376 34546 22428 34552
rect 22204 34218 22232 34546
rect 22204 34190 22324 34218
rect 22192 34060 22244 34066
rect 22192 34002 22244 34008
rect 22204 33114 22232 34002
rect 22296 33946 22324 34190
rect 22388 34134 22416 34546
rect 22376 34128 22428 34134
rect 22376 34070 22428 34076
rect 22376 33992 22428 33998
rect 22296 33940 22376 33946
rect 22296 33934 22428 33940
rect 22296 33918 22416 33934
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22192 33108 22244 33114
rect 22192 33050 22244 33056
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 22112 31686 22140 31758
rect 22100 31680 22152 31686
rect 22100 31622 22152 31628
rect 22112 31142 22140 31622
rect 22192 31272 22244 31278
rect 22192 31214 22244 31220
rect 22100 31136 22152 31142
rect 22100 31078 22152 31084
rect 22008 30864 22060 30870
rect 22008 30806 22060 30812
rect 21916 29232 21968 29238
rect 21916 29174 21968 29180
rect 21824 29164 21876 29170
rect 21824 29106 21876 29112
rect 21732 28076 21784 28082
rect 21732 28018 21784 28024
rect 21836 25906 21864 29106
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 21928 26586 21956 26930
rect 21916 26580 21968 26586
rect 21916 26522 21968 26528
rect 21824 25900 21876 25906
rect 21824 25842 21876 25848
rect 21836 24750 21864 25842
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 21744 22234 21772 23054
rect 21732 22228 21784 22234
rect 21732 22170 21784 22176
rect 22020 22094 22048 30806
rect 22112 29170 22140 31078
rect 22204 30938 22232 31214
rect 22192 30932 22244 30938
rect 22192 30874 22244 30880
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22296 28626 22324 33798
rect 22376 33312 22428 33318
rect 22376 33254 22428 33260
rect 22388 32978 22416 33254
rect 22376 32972 22428 32978
rect 22376 32914 22428 32920
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 22376 32224 22428 32230
rect 22376 32166 22428 32172
rect 22468 32224 22520 32230
rect 22468 32166 22520 32172
rect 22388 31822 22416 32166
rect 22480 31890 22508 32166
rect 22572 31890 22600 32370
rect 22468 31884 22520 31890
rect 22468 31826 22520 31832
rect 22560 31884 22612 31890
rect 22560 31826 22612 31832
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22376 31408 22428 31414
rect 22376 31350 22428 31356
rect 22560 31408 22612 31414
rect 22560 31350 22612 31356
rect 22388 30682 22416 31350
rect 22572 30938 22600 31350
rect 22560 30932 22612 30938
rect 22560 30874 22612 30880
rect 22560 30728 22612 30734
rect 22388 30676 22560 30682
rect 22388 30670 22612 30676
rect 22388 30654 22600 30670
rect 22284 28620 22336 28626
rect 22284 28562 22336 28568
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 22204 28218 22232 28494
rect 22192 28212 22244 28218
rect 22192 28154 22244 28160
rect 22100 28144 22152 28150
rect 22100 28086 22152 28092
rect 22112 26994 22140 28086
rect 22192 27940 22244 27946
rect 22192 27882 22244 27888
rect 22204 27062 22232 27882
rect 22296 27470 22324 28562
rect 22284 27464 22336 27470
rect 22284 27406 22336 27412
rect 22192 27056 22244 27062
rect 22192 26998 22244 27004
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 22112 26897 22140 26930
rect 22098 26888 22154 26897
rect 22098 26823 22154 26832
rect 22100 26784 22152 26790
rect 22100 26726 22152 26732
rect 22112 25974 22140 26726
rect 22204 26382 22232 26998
rect 22192 26376 22244 26382
rect 22192 26318 22244 26324
rect 22204 26042 22232 26318
rect 22192 26036 22244 26042
rect 22192 25978 22244 25984
rect 22100 25968 22152 25974
rect 22100 25910 22152 25916
rect 22100 24676 22152 24682
rect 22100 24618 22152 24624
rect 22112 23662 22140 24618
rect 22388 24614 22416 30654
rect 22664 29850 22692 35006
rect 22744 33516 22796 33522
rect 22744 33458 22796 33464
rect 22756 32570 22784 33458
rect 22744 32564 22796 32570
rect 22744 32506 22796 32512
rect 22756 31822 22784 32506
rect 22744 31816 22796 31822
rect 22744 31758 22796 31764
rect 22652 29844 22704 29850
rect 22652 29786 22704 29792
rect 22558 29064 22614 29073
rect 22664 29034 22692 29786
rect 22558 28999 22614 29008
rect 22652 29028 22704 29034
rect 22572 28937 22600 28999
rect 22652 28970 22704 28976
rect 22558 28928 22614 28937
rect 22558 28863 22614 28872
rect 22572 26994 22600 28863
rect 22664 28558 22692 28970
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 22560 26988 22612 26994
rect 22560 26930 22612 26936
rect 22848 26330 22876 37606
rect 23216 37330 23244 38218
rect 23204 37324 23256 37330
rect 23204 37266 23256 37272
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 23032 36378 23060 37198
rect 23020 36372 23072 36378
rect 23020 36314 23072 36320
rect 23216 35766 23244 37266
rect 24136 37126 24164 38830
rect 24504 38350 24532 45766
rect 25240 45490 25268 45902
rect 25412 45892 25464 45898
rect 25412 45834 25464 45840
rect 25228 45484 25280 45490
rect 25228 45426 25280 45432
rect 25424 45082 25452 45834
rect 26712 45554 26740 49286
rect 27038 49200 27150 49286
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49314 31014 50000
rect 30760 49286 31014 49314
rect 28368 47054 28396 49200
rect 29656 47054 29684 49200
rect 30104 47184 30156 47190
rect 30104 47126 30156 47132
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 26436 45526 26740 45554
rect 25412 45076 25464 45082
rect 25412 45018 25464 45024
rect 25320 44872 25372 44878
rect 25320 44814 25372 44820
rect 25332 43722 25360 44814
rect 25780 43784 25832 43790
rect 25780 43726 25832 43732
rect 25320 43716 25372 43722
rect 25320 43658 25372 43664
rect 24584 39364 24636 39370
rect 24584 39306 24636 39312
rect 24596 39098 24624 39306
rect 24584 39092 24636 39098
rect 24584 39034 24636 39040
rect 24676 38956 24728 38962
rect 24676 38898 24728 38904
rect 24492 38344 24544 38350
rect 24492 38286 24544 38292
rect 24492 38208 24544 38214
rect 24492 38150 24544 38156
rect 24504 37942 24532 38150
rect 24492 37936 24544 37942
rect 24492 37878 24544 37884
rect 24400 37664 24452 37670
rect 24400 37606 24452 37612
rect 24412 37466 24440 37606
rect 24400 37460 24452 37466
rect 24400 37402 24452 37408
rect 24308 37188 24360 37194
rect 24308 37130 24360 37136
rect 24124 37120 24176 37126
rect 24124 37062 24176 37068
rect 23480 36168 23532 36174
rect 23480 36110 23532 36116
rect 23204 35760 23256 35766
rect 23204 35702 23256 35708
rect 23492 35698 23520 36110
rect 24136 35834 24164 37062
rect 24320 36786 24348 37130
rect 24308 36780 24360 36786
rect 24308 36722 24360 36728
rect 24124 35828 24176 35834
rect 24124 35770 24176 35776
rect 23480 35692 23532 35698
rect 23480 35634 23532 35640
rect 23388 34672 23440 34678
rect 23388 34614 23440 34620
rect 22928 34604 22980 34610
rect 22928 34546 22980 34552
rect 22940 34066 22968 34546
rect 23400 34202 23428 34614
rect 23492 34474 23520 35634
rect 24032 35012 24084 35018
rect 24032 34954 24084 34960
rect 24044 34678 24072 34954
rect 24032 34672 24084 34678
rect 24032 34614 24084 34620
rect 23664 34604 23716 34610
rect 23664 34546 23716 34552
rect 23572 34536 23624 34542
rect 23572 34478 23624 34484
rect 23480 34468 23532 34474
rect 23480 34410 23532 34416
rect 23388 34196 23440 34202
rect 23388 34138 23440 34144
rect 22928 34060 22980 34066
rect 22928 34002 22980 34008
rect 23112 33312 23164 33318
rect 23112 33254 23164 33260
rect 23124 32570 23152 33254
rect 23112 32564 23164 32570
rect 23112 32506 23164 32512
rect 22928 32428 22980 32434
rect 22928 32370 22980 32376
rect 22940 32026 22968 32370
rect 22928 32020 22980 32026
rect 22928 31962 22980 31968
rect 23400 31929 23428 34138
rect 23584 33998 23612 34478
rect 23676 34202 23704 34546
rect 24320 34406 24348 36722
rect 24412 36242 24440 37402
rect 24688 37262 24716 38898
rect 24952 37800 25004 37806
rect 24952 37742 25004 37748
rect 24676 37256 24728 37262
rect 24676 37198 24728 37204
rect 24768 37256 24820 37262
rect 24768 37198 24820 37204
rect 24400 36236 24452 36242
rect 24400 36178 24452 36184
rect 24412 35698 24440 36178
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 24492 35828 24544 35834
rect 24492 35770 24544 35776
rect 24400 35692 24452 35698
rect 24400 35634 24452 35640
rect 24504 35578 24532 35770
rect 24596 35698 24624 36110
rect 24584 35692 24636 35698
rect 24584 35634 24636 35640
rect 24412 35550 24532 35578
rect 24412 35494 24440 35550
rect 24400 35488 24452 35494
rect 24400 35430 24452 35436
rect 24596 34746 24624 35634
rect 24780 35222 24808 37198
rect 24860 37120 24912 37126
rect 24860 37062 24912 37068
rect 24768 35216 24820 35222
rect 24768 35158 24820 35164
rect 24400 34740 24452 34746
rect 24400 34682 24452 34688
rect 24584 34740 24636 34746
rect 24584 34682 24636 34688
rect 24308 34400 24360 34406
rect 24308 34342 24360 34348
rect 23664 34196 23716 34202
rect 23664 34138 23716 34144
rect 23572 33992 23624 33998
rect 23572 33934 23624 33940
rect 23676 33386 23704 34138
rect 23572 33380 23624 33386
rect 23572 33322 23624 33328
rect 23664 33380 23716 33386
rect 23664 33322 23716 33328
rect 23584 32434 23612 33322
rect 23848 33312 23900 33318
rect 23848 33254 23900 33260
rect 23860 32502 23888 33254
rect 23848 32496 23900 32502
rect 23848 32438 23900 32444
rect 23572 32428 23624 32434
rect 23572 32370 23624 32376
rect 23940 32224 23992 32230
rect 23940 32166 23992 32172
rect 23386 31920 23442 31929
rect 23952 31890 23980 32166
rect 23386 31855 23442 31864
rect 23940 31884 23992 31890
rect 23940 31826 23992 31832
rect 23848 31816 23900 31822
rect 23848 31758 23900 31764
rect 23860 31482 23888 31758
rect 24412 31482 24440 34682
rect 24596 34202 24624 34682
rect 24780 34610 24808 35158
rect 24872 35086 24900 37062
rect 24964 36378 24992 37742
rect 25504 37664 25556 37670
rect 25504 37606 25556 37612
rect 25516 36786 25544 37606
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 24952 36372 25004 36378
rect 24952 36314 25004 36320
rect 25516 36174 25544 36722
rect 25596 36576 25648 36582
rect 25596 36518 25648 36524
rect 25320 36168 25372 36174
rect 25240 36128 25320 36156
rect 24952 35624 25004 35630
rect 24952 35566 25004 35572
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 24768 34604 24820 34610
rect 24768 34546 24820 34552
rect 24584 34196 24636 34202
rect 24584 34138 24636 34144
rect 24964 33674 24992 35566
rect 25136 35080 25188 35086
rect 25136 35022 25188 35028
rect 25148 34678 25176 35022
rect 25240 34746 25268 36128
rect 25320 36110 25372 36116
rect 25504 36168 25556 36174
rect 25504 36110 25556 36116
rect 25320 35556 25372 35562
rect 25320 35498 25372 35504
rect 25228 34740 25280 34746
rect 25228 34682 25280 34688
rect 25136 34672 25188 34678
rect 25136 34614 25188 34620
rect 25332 34610 25360 35498
rect 25608 35154 25636 36518
rect 25688 35624 25740 35630
rect 25688 35566 25740 35572
rect 25596 35148 25648 35154
rect 25596 35090 25648 35096
rect 25608 34746 25636 35090
rect 25596 34740 25648 34746
rect 25596 34682 25648 34688
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25504 34604 25556 34610
rect 25504 34546 25556 34552
rect 25516 34354 25544 34546
rect 25240 34326 25544 34354
rect 24964 33646 25176 33674
rect 24676 33584 24728 33590
rect 24676 33526 24728 33532
rect 24492 32904 24544 32910
rect 24688 32892 24716 33526
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24872 33114 24900 33458
rect 24952 33312 25004 33318
rect 24952 33254 25004 33260
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24544 32864 24716 32892
rect 24492 32846 24544 32852
rect 24584 32360 24636 32366
rect 24584 32302 24636 32308
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 24400 31476 24452 31482
rect 24400 31418 24452 31424
rect 24596 31346 24624 32302
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 24688 30938 24716 32864
rect 24964 32434 24992 33254
rect 24952 32428 25004 32434
rect 24952 32370 25004 32376
rect 24860 32292 24912 32298
rect 24860 32234 24912 32240
rect 24872 31278 24900 32234
rect 25148 32230 25176 33646
rect 25136 32224 25188 32230
rect 25136 32166 25188 32172
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 24860 31272 24912 31278
rect 24860 31214 24912 31220
rect 24676 30932 24728 30938
rect 24676 30874 24728 30880
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24872 29714 24900 30194
rect 24860 29708 24912 29714
rect 24860 29650 24912 29656
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 23112 29504 23164 29510
rect 23112 29446 23164 29452
rect 23020 29232 23072 29238
rect 23124 29220 23152 29446
rect 23072 29192 23152 29220
rect 23020 29174 23072 29180
rect 22928 29096 22980 29102
rect 22928 29038 22980 29044
rect 22940 28762 22968 29038
rect 22928 28756 22980 28762
rect 22928 28698 22980 28704
rect 23124 28558 23152 29192
rect 24596 29170 24624 29582
rect 24032 29164 24084 29170
rect 24032 29106 24084 29112
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 23480 28620 23532 28626
rect 23480 28562 23532 28568
rect 23112 28552 23164 28558
rect 23112 28494 23164 28500
rect 23492 28150 23520 28562
rect 23480 28144 23532 28150
rect 23480 28086 23532 28092
rect 22928 28008 22980 28014
rect 22928 27950 22980 27956
rect 22940 27334 22968 27950
rect 23020 27872 23072 27878
rect 23020 27814 23072 27820
rect 23940 27872 23992 27878
rect 23940 27814 23992 27820
rect 23032 27470 23060 27814
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 23952 27402 23980 27814
rect 23940 27396 23992 27402
rect 23940 27338 23992 27344
rect 22928 27328 22980 27334
rect 22928 27270 22980 27276
rect 22940 27130 22968 27270
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 22848 26302 22968 26330
rect 22836 25968 22888 25974
rect 22836 25910 22888 25916
rect 22848 25498 22876 25910
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 22940 24818 22968 26302
rect 24044 26042 24072 29106
rect 24400 28960 24452 28966
rect 24400 28902 24452 28908
rect 24412 28150 24440 28902
rect 24492 28484 24544 28490
rect 24492 28426 24544 28432
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24504 27062 24532 28426
rect 24596 28422 24624 29106
rect 24584 28416 24636 28422
rect 24584 28358 24636 28364
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 24688 27674 24716 28018
rect 24768 28008 24820 28014
rect 24768 27950 24820 27956
rect 24676 27668 24728 27674
rect 24676 27610 24728 27616
rect 24492 27056 24544 27062
rect 24492 26998 24544 27004
rect 24780 26994 24808 27950
rect 24952 27940 25004 27946
rect 24952 27882 25004 27888
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24676 26512 24728 26518
rect 24676 26454 24728 26460
rect 24032 26036 24084 26042
rect 24032 25978 24084 25984
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23400 25294 23428 25842
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23400 24954 23428 25230
rect 23388 24948 23440 24954
rect 23388 24890 23440 24896
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22940 24206 22968 24754
rect 23020 24608 23072 24614
rect 23020 24550 23072 24556
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22112 22982 22140 23598
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 21928 22066 22048 22094
rect 21730 21584 21786 21593
rect 21928 21554 21956 22066
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 21730 21519 21786 21528
rect 21916 21548 21968 21554
rect 21744 21486 21772 21519
rect 21916 21490 21968 21496
rect 21732 21480 21784 21486
rect 21732 21422 21784 21428
rect 22020 20466 22048 21966
rect 22112 21962 22140 22918
rect 22192 22500 22244 22506
rect 22284 22500 22336 22506
rect 22244 22460 22284 22488
rect 22192 22442 22244 22448
rect 22284 22442 22336 22448
rect 22100 21956 22152 21962
rect 22100 21898 22152 21904
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22296 21554 22324 21898
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 22020 18698 22048 20402
rect 22112 20262 22140 20810
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 22008 18692 22060 18698
rect 22008 18634 22060 18640
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 22112 17882 22140 18158
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22284 17808 22336 17814
rect 22284 17750 22336 17756
rect 22192 17264 22244 17270
rect 21652 17224 21772 17252
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21652 15502 21680 16050
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21560 14618 21588 15030
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21560 14074 21588 14554
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21560 13326 21588 14010
rect 21652 13394 21680 14214
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21744 2310 21772 17224
rect 22192 17206 22244 17212
rect 21916 16992 21968 16998
rect 21916 16934 21968 16940
rect 21928 16726 21956 16934
rect 21916 16720 21968 16726
rect 21916 16662 21968 16668
rect 22204 16454 22232 17206
rect 22296 17202 22324 17750
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 22112 15706 22140 15982
rect 22204 15910 22232 16390
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 21824 15360 21876 15366
rect 21824 15302 21876 15308
rect 21836 13938 21864 15302
rect 21928 15094 21956 15370
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 21928 14482 21956 15030
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 22020 14414 22048 14758
rect 22204 14550 22232 15846
rect 22296 15638 22324 16458
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21836 13530 21864 13670
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22296 11354 22324 11630
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21836 3058 21864 3878
rect 21928 3194 21956 4558
rect 22204 4010 22232 11086
rect 22388 6914 22416 23598
rect 22756 23186 22784 24006
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22836 22976 22888 22982
rect 22836 22918 22888 22924
rect 22756 22778 22784 22918
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 22848 22710 22876 22918
rect 22836 22704 22888 22710
rect 22466 22672 22522 22681
rect 22836 22646 22888 22652
rect 22466 22607 22468 22616
rect 22520 22607 22522 22616
rect 22468 22578 22520 22584
rect 22652 22500 22704 22506
rect 22652 22442 22704 22448
rect 22664 22030 22692 22442
rect 23032 22386 23060 24550
rect 23400 24206 23428 24890
rect 24688 24750 24716 26454
rect 24780 26314 24808 26930
rect 24872 26382 24900 27814
rect 24964 27470 24992 27882
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 24952 27328 25004 27334
rect 24952 27270 25004 27276
rect 24964 26926 24992 27270
rect 24952 26920 25004 26926
rect 24952 26862 25004 26868
rect 24952 26444 25004 26450
rect 24952 26386 25004 26392
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24768 26308 24820 26314
rect 24768 26250 24820 26256
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 23124 23118 23152 23462
rect 23204 23180 23256 23186
rect 23204 23122 23256 23128
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 22848 22358 23060 22386
rect 22652 22024 22704 22030
rect 22466 21992 22522 22001
rect 22652 21966 22704 21972
rect 22466 21927 22522 21936
rect 22480 21894 22508 21927
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22572 20874 22600 21286
rect 22560 20868 22612 20874
rect 22560 20810 22612 20816
rect 22664 20398 22692 21966
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 22744 19984 22796 19990
rect 22744 19926 22796 19932
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22664 19378 22692 19722
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22756 19310 22784 19926
rect 22848 19514 22876 22358
rect 23112 22024 23164 22030
rect 23110 21992 23112 22001
rect 23164 21992 23166 22001
rect 23110 21927 23166 21936
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 23124 21554 23152 21830
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 23216 20942 23244 23122
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23308 21876 23336 22918
rect 23572 22636 23624 22642
rect 23624 22596 23704 22624
rect 23572 22578 23624 22584
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23492 22030 23520 22374
rect 23480 22024 23532 22030
rect 23480 21966 23532 21972
rect 23388 21888 23440 21894
rect 23308 21848 23388 21876
rect 23388 21830 23440 21836
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23584 21554 23612 21830
rect 23676 21554 23704 22596
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 23952 21554 23980 22170
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23308 21146 23336 21490
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22560 18352 22612 18358
rect 22560 18294 22612 18300
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22480 18086 22508 18158
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22572 17882 22600 18294
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22664 17746 22692 18022
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22664 17134 22692 17682
rect 22652 17128 22704 17134
rect 22652 17070 22704 17076
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22480 11830 22508 17002
rect 22664 16794 22692 17070
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22572 15706 22600 16118
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22468 11824 22520 11830
rect 22468 11766 22520 11772
rect 22756 6914 22784 19246
rect 22848 18766 22876 19450
rect 24136 19378 24164 24006
rect 24492 22568 24544 22574
rect 24492 22510 24544 22516
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24504 22234 24532 22510
rect 24492 22228 24544 22234
rect 24492 22170 24544 22176
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24308 21956 24360 21962
rect 24308 21898 24360 21904
rect 24320 21690 24348 21898
rect 24308 21684 24360 21690
rect 24308 21626 24360 21632
rect 24688 21146 24716 21966
rect 24780 21690 24808 22510
rect 24964 22094 24992 26386
rect 25056 24750 25084 31758
rect 25240 31686 25268 34326
rect 25700 34202 25728 35566
rect 25688 34196 25740 34202
rect 25688 34138 25740 34144
rect 25504 33992 25556 33998
rect 25504 33934 25556 33940
rect 25412 32768 25464 32774
rect 25412 32710 25464 32716
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25228 31680 25280 31686
rect 25228 31622 25280 31628
rect 25240 30734 25268 31622
rect 25228 30728 25280 30734
rect 25228 30670 25280 30676
rect 25332 30666 25360 32166
rect 25424 31278 25452 32710
rect 25516 31346 25544 33934
rect 25688 33108 25740 33114
rect 25688 33050 25740 33056
rect 25596 32496 25648 32502
rect 25596 32438 25648 32444
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25412 31272 25464 31278
rect 25412 31214 25464 31220
rect 25516 30938 25544 31282
rect 25504 30932 25556 30938
rect 25504 30874 25556 30880
rect 25320 30660 25372 30666
rect 25320 30602 25372 30608
rect 25332 30258 25360 30602
rect 25608 30598 25636 32438
rect 25596 30592 25648 30598
rect 25596 30534 25648 30540
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 25504 30252 25556 30258
rect 25504 30194 25556 30200
rect 25412 30184 25464 30190
rect 25412 30126 25464 30132
rect 25320 30048 25372 30054
rect 25320 29990 25372 29996
rect 25136 29096 25188 29102
rect 25136 29038 25188 29044
rect 25148 27946 25176 29038
rect 25136 27940 25188 27946
rect 25136 27882 25188 27888
rect 25136 27056 25188 27062
rect 25136 26998 25188 27004
rect 25148 26586 25176 26998
rect 25136 26580 25188 26586
rect 25136 26522 25188 26528
rect 25136 25696 25188 25702
rect 25136 25638 25188 25644
rect 25148 25226 25176 25638
rect 25136 25220 25188 25226
rect 25136 25162 25188 25168
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 25332 22094 25360 29990
rect 25424 29306 25452 30126
rect 25412 29300 25464 29306
rect 25412 29242 25464 29248
rect 25424 28558 25452 29242
rect 25516 28966 25544 30194
rect 25596 29640 25648 29646
rect 25596 29582 25648 29588
rect 25504 28960 25556 28966
rect 25504 28902 25556 28908
rect 25516 28626 25544 28902
rect 25504 28620 25556 28626
rect 25504 28562 25556 28568
rect 25412 28552 25464 28558
rect 25412 28494 25464 28500
rect 25608 28218 25636 29582
rect 25700 29102 25728 33050
rect 25792 30054 25820 43726
rect 26240 37188 26292 37194
rect 26240 37130 26292 37136
rect 26252 36922 26280 37130
rect 26240 36916 26292 36922
rect 26240 36858 26292 36864
rect 26240 36780 26292 36786
rect 26240 36722 26292 36728
rect 25964 36168 26016 36174
rect 25964 36110 26016 36116
rect 25872 34944 25924 34950
rect 25872 34886 25924 34892
rect 25884 33930 25912 34886
rect 25976 34610 26004 36110
rect 26252 35630 26280 36722
rect 26240 35624 26292 35630
rect 26240 35566 26292 35572
rect 26332 35556 26384 35562
rect 26332 35498 26384 35504
rect 26148 35488 26200 35494
rect 26148 35430 26200 35436
rect 25964 34604 26016 34610
rect 25964 34546 26016 34552
rect 26056 34536 26108 34542
rect 26056 34478 26108 34484
rect 25964 34468 26016 34474
rect 25964 34410 26016 34416
rect 25872 33924 25924 33930
rect 25872 33866 25924 33872
rect 25976 33862 26004 34410
rect 25964 33856 26016 33862
rect 25964 33798 26016 33804
rect 25872 32496 25924 32502
rect 25872 32438 25924 32444
rect 25884 31890 25912 32438
rect 25964 32360 26016 32366
rect 25964 32302 26016 32308
rect 25872 31884 25924 31890
rect 25872 31826 25924 31832
rect 25976 31754 26004 32302
rect 25884 31726 26004 31754
rect 25884 31142 25912 31726
rect 25872 31136 25924 31142
rect 25872 31078 25924 31084
rect 25780 30048 25832 30054
rect 25780 29990 25832 29996
rect 25688 29096 25740 29102
rect 25688 29038 25740 29044
rect 25596 28212 25648 28218
rect 25596 28154 25648 28160
rect 25608 27606 25636 28154
rect 25596 27600 25648 27606
rect 25596 27542 25648 27548
rect 25780 27600 25832 27606
rect 25780 27542 25832 27548
rect 25596 27464 25648 27470
rect 25596 27406 25648 27412
rect 25504 27328 25556 27334
rect 25504 27270 25556 27276
rect 25516 25906 25544 27270
rect 25608 26296 25636 27406
rect 25792 27062 25820 27542
rect 25780 27056 25832 27062
rect 25686 27024 25742 27033
rect 25780 26998 25832 27004
rect 25686 26959 25742 26968
rect 25700 26926 25728 26959
rect 25688 26920 25740 26926
rect 25884 26897 25912 31078
rect 25964 30592 26016 30598
rect 25964 30534 26016 30540
rect 25976 30258 26004 30534
rect 25964 30252 26016 30258
rect 25964 30194 26016 30200
rect 25976 27334 26004 30194
rect 25964 27328 26016 27334
rect 25964 27270 26016 27276
rect 25688 26862 25740 26868
rect 25870 26888 25926 26897
rect 25870 26823 25926 26832
rect 25688 26784 25740 26790
rect 25688 26726 25740 26732
rect 25780 26784 25832 26790
rect 25884 26772 25912 26823
rect 25964 26784 26016 26790
rect 25884 26744 25964 26772
rect 25780 26726 25832 26732
rect 25964 26726 26016 26732
rect 25700 26518 25728 26726
rect 25688 26512 25740 26518
rect 25688 26454 25740 26460
rect 25688 26308 25740 26314
rect 25608 26268 25688 26296
rect 25688 26250 25740 26256
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 25412 25696 25464 25702
rect 25412 25638 25464 25644
rect 25424 24886 25452 25638
rect 25700 25430 25728 26250
rect 25792 25498 25820 26726
rect 25780 25492 25832 25498
rect 25780 25434 25832 25440
rect 25688 25424 25740 25430
rect 25688 25366 25740 25372
rect 25412 24880 25464 24886
rect 25412 24822 25464 24828
rect 26068 24698 26096 34478
rect 26160 33114 26188 35430
rect 26344 35290 26372 35498
rect 26332 35284 26384 35290
rect 26332 35226 26384 35232
rect 26332 35080 26384 35086
rect 26332 35022 26384 35028
rect 26344 34678 26372 35022
rect 26332 34672 26384 34678
rect 26332 34614 26384 34620
rect 26332 34536 26384 34542
rect 26332 34478 26384 34484
rect 26148 33108 26200 33114
rect 26148 33050 26200 33056
rect 26344 32978 26372 34478
rect 26332 32972 26384 32978
rect 26332 32914 26384 32920
rect 26240 32836 26292 32842
rect 26240 32778 26292 32784
rect 26252 32502 26280 32778
rect 26240 32496 26292 32502
rect 26240 32438 26292 32444
rect 26344 30870 26372 32914
rect 26332 30864 26384 30870
rect 26332 30806 26384 30812
rect 26344 28082 26372 30806
rect 26332 28076 26384 28082
rect 26332 28018 26384 28024
rect 26344 27470 26372 28018
rect 26332 27464 26384 27470
rect 26332 27406 26384 27412
rect 26148 27396 26200 27402
rect 26148 27338 26200 27344
rect 26160 26314 26188 27338
rect 26330 27024 26386 27033
rect 26330 26959 26386 26968
rect 26344 26858 26372 26959
rect 26240 26852 26292 26858
rect 26240 26794 26292 26800
rect 26332 26852 26384 26858
rect 26332 26794 26384 26800
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 26160 24954 26188 26250
rect 26148 24948 26200 24954
rect 26148 24890 26200 24896
rect 26068 24670 26188 24698
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 25596 23860 25648 23866
rect 25596 23802 25648 23808
rect 25608 23594 25636 23802
rect 26068 23798 26096 24006
rect 26056 23792 26108 23798
rect 26056 23734 26108 23740
rect 25596 23588 25648 23594
rect 25596 23530 25648 23536
rect 25412 23520 25464 23526
rect 25412 23462 25464 23468
rect 25424 23186 25452 23462
rect 25412 23180 25464 23186
rect 25412 23122 25464 23128
rect 25964 23180 26016 23186
rect 25964 23122 26016 23128
rect 25780 22704 25832 22710
rect 25780 22646 25832 22652
rect 25792 22098 25820 22646
rect 24964 22066 25084 22094
rect 25332 22066 25452 22094
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24676 21140 24728 21146
rect 24676 21082 24728 21088
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24504 19514 24532 19790
rect 24492 19508 24544 19514
rect 24492 19450 24544 19456
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23676 18970 23704 19246
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 22928 18692 22980 18698
rect 22928 18634 22980 18640
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 22848 15026 22876 15438
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22836 14816 22888 14822
rect 22836 14758 22888 14764
rect 22848 14006 22876 14758
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22296 6886 22416 6914
rect 22664 6886 22784 6914
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22296 3602 22324 6886
rect 22376 4480 22428 4486
rect 22376 4422 22428 4428
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 21916 3188 21968 3194
rect 21916 3130 21968 3136
rect 22006 3088 22062 3097
rect 21824 3052 21876 3058
rect 22006 3023 22062 3032
rect 21824 2994 21876 3000
rect 22020 2922 22048 3023
rect 22008 2916 22060 2922
rect 22008 2858 22060 2864
rect 22112 2650 22140 3470
rect 22388 3058 22416 4422
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22572 3194 22600 4014
rect 22664 3670 22692 6886
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22652 3664 22704 3670
rect 22652 3606 22704 3612
rect 22848 3534 22876 3878
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22940 3126 22968 18634
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 23032 17678 23060 18566
rect 23584 18222 23612 18702
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 23572 18216 23624 18222
rect 23572 18158 23624 18164
rect 23584 17678 23612 18158
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23112 17264 23164 17270
rect 23112 17206 23164 17212
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23032 16794 23060 17138
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23124 14618 23152 17206
rect 23204 17060 23256 17066
rect 23204 17002 23256 17008
rect 23216 16726 23244 17002
rect 23400 16726 23428 17614
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24136 17202 24164 17478
rect 24780 17338 24808 18226
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24872 17746 24900 18022
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 23940 16992 23992 16998
rect 23940 16934 23992 16940
rect 23952 16794 23980 16934
rect 24044 16794 24072 17070
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 23204 16720 23256 16726
rect 23204 16662 23256 16668
rect 23388 16720 23440 16726
rect 23388 16662 23440 16668
rect 23400 15026 23428 16662
rect 23952 16658 23980 16730
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23768 15094 23796 16594
rect 24044 16182 24072 16730
rect 24872 16590 24900 17682
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24032 16176 24084 16182
rect 24032 16118 24084 16124
rect 24964 15978 24992 17478
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24400 15360 24452 15366
rect 24400 15302 24452 15308
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23400 14006 23428 14962
rect 23768 14482 23796 15030
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 24308 14408 24360 14414
rect 24308 14350 24360 14356
rect 24320 14074 24348 14350
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 24412 13938 24440 15302
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24412 13462 24440 13874
rect 24400 13456 24452 13462
rect 24400 13398 24452 13404
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 22928 3120 22980 3126
rect 22928 3062 22980 3068
rect 23216 3058 23244 3470
rect 23400 3126 23428 3878
rect 23388 3120 23440 3126
rect 23480 3120 23532 3126
rect 23388 3062 23440 3068
rect 23478 3088 23480 3097
rect 23532 3088 23534 3097
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 23204 3052 23256 3058
rect 23478 3023 23534 3032
rect 23204 2994 23256 3000
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 23480 2916 23532 2922
rect 23480 2858 23532 2864
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 21732 2304 21784 2310
rect 21732 2246 21784 2252
rect 21180 2032 21232 2038
rect 21180 1974 21232 1980
rect 21928 800 21956 2314
rect 22572 800 22600 2858
rect 23492 2650 23520 2858
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 23952 2514 23980 11630
rect 24308 4072 24360 4078
rect 24308 4014 24360 4020
rect 24320 3670 24348 4014
rect 24860 3936 24912 3942
rect 24860 3878 24912 3884
rect 24308 3664 24360 3670
rect 24308 3606 24360 3612
rect 24872 3602 24900 3878
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 25056 2582 25084 22066
rect 25228 21548 25280 21554
rect 25228 21490 25280 21496
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 25148 19718 25176 20402
rect 25240 20330 25268 21490
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25332 20534 25360 20878
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 25228 20324 25280 20330
rect 25228 20266 25280 20272
rect 25240 19786 25268 20266
rect 25228 19780 25280 19786
rect 25228 19722 25280 19728
rect 25136 19712 25188 19718
rect 25136 19654 25188 19660
rect 25424 17542 25452 22066
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25872 22092 25924 22098
rect 25872 22034 25924 22040
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 25516 21554 25544 21966
rect 25884 21962 25912 22034
rect 25872 21956 25924 21962
rect 25872 21898 25924 21904
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25516 21010 25544 21286
rect 25504 21004 25556 21010
rect 25504 20946 25556 20952
rect 25596 20256 25648 20262
rect 25596 20198 25648 20204
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25608 19922 25636 20198
rect 25596 19916 25648 19922
rect 25596 19858 25648 19864
rect 25884 19786 25912 20198
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 25780 19712 25832 19718
rect 25780 19654 25832 19660
rect 25792 18290 25820 19654
rect 25780 18284 25832 18290
rect 25780 18226 25832 18232
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 25412 17536 25464 17542
rect 25412 17478 25464 17484
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 25148 15978 25176 17070
rect 25424 16454 25452 17478
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25516 16794 25544 17138
rect 25608 16998 25636 17682
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25136 15972 25188 15978
rect 25136 15914 25188 15920
rect 25792 15502 25820 18226
rect 25872 17604 25924 17610
rect 25872 17546 25924 17552
rect 25884 17202 25912 17546
rect 25872 17196 25924 17202
rect 25872 17138 25924 17144
rect 25780 15496 25832 15502
rect 25780 15438 25832 15444
rect 25136 14340 25188 14346
rect 25136 14282 25188 14288
rect 25148 14074 25176 14282
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25596 3936 25648 3942
rect 25596 3878 25648 3884
rect 25608 3670 25636 3878
rect 25700 3670 25728 4082
rect 25976 3942 26004 23122
rect 26160 22094 26188 24670
rect 26252 23186 26280 26794
rect 26436 24682 26464 45526
rect 26976 38412 27028 38418
rect 26976 38354 27028 38360
rect 26988 37874 27016 38354
rect 26976 37868 27028 37874
rect 26976 37810 27028 37816
rect 27620 37664 27672 37670
rect 27620 37606 27672 37612
rect 29460 37664 29512 37670
rect 29460 37606 29512 37612
rect 27632 37194 27660 37606
rect 28540 37256 28592 37262
rect 28540 37198 28592 37204
rect 28724 37256 28776 37262
rect 28724 37198 28776 37204
rect 27620 37188 27672 37194
rect 27620 37130 27672 37136
rect 27528 37120 27580 37126
rect 27528 37062 27580 37068
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 28448 37120 28500 37126
rect 28448 37062 28500 37068
rect 27540 36786 27568 37062
rect 27528 36780 27580 36786
rect 27528 36722 27580 36728
rect 27344 36236 27396 36242
rect 27344 36178 27396 36184
rect 27436 36236 27488 36242
rect 27436 36178 27488 36184
rect 26700 36168 26752 36174
rect 26700 36110 26752 36116
rect 26608 36032 26660 36038
rect 26608 35974 26660 35980
rect 26516 35692 26568 35698
rect 26516 35634 26568 35640
rect 26528 35086 26556 35634
rect 26620 35222 26648 35974
rect 26608 35216 26660 35222
rect 26608 35158 26660 35164
rect 26620 35086 26648 35158
rect 26516 35080 26568 35086
rect 26516 35022 26568 35028
rect 26608 35080 26660 35086
rect 26608 35022 26660 35028
rect 26528 30666 26556 35022
rect 26712 34678 26740 36110
rect 26792 35760 26844 35766
rect 26792 35702 26844 35708
rect 26700 34672 26752 34678
rect 26700 34614 26752 34620
rect 26804 34542 26832 35702
rect 27356 35562 27384 36178
rect 27448 35698 27476 36178
rect 27540 35766 27568 36722
rect 27724 36038 27752 37062
rect 28460 36854 28488 37062
rect 28448 36848 28500 36854
rect 28448 36790 28500 36796
rect 28552 36378 28580 37198
rect 28736 36922 28764 37198
rect 28724 36916 28776 36922
rect 28724 36858 28776 36864
rect 29472 36854 29500 37606
rect 29920 37324 29972 37330
rect 29920 37266 29972 37272
rect 29644 37256 29696 37262
rect 29644 37198 29696 37204
rect 29460 36848 29512 36854
rect 29460 36790 29512 36796
rect 28540 36372 28592 36378
rect 28540 36314 28592 36320
rect 27896 36168 27948 36174
rect 27896 36110 27948 36116
rect 29000 36168 29052 36174
rect 29000 36110 29052 36116
rect 27712 36032 27764 36038
rect 27712 35974 27764 35980
rect 27528 35760 27580 35766
rect 27528 35702 27580 35708
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27344 35556 27396 35562
rect 27344 35498 27396 35504
rect 27252 35148 27304 35154
rect 27252 35090 27304 35096
rect 26884 35080 26936 35086
rect 26884 35022 26936 35028
rect 26896 34610 26924 35022
rect 26884 34604 26936 34610
rect 26884 34546 26936 34552
rect 26792 34536 26844 34542
rect 26792 34478 26844 34484
rect 26884 32292 26936 32298
rect 26884 32234 26936 32240
rect 26896 31958 26924 32234
rect 26884 31952 26936 31958
rect 26884 31894 26936 31900
rect 27160 31476 27212 31482
rect 27160 31418 27212 31424
rect 26974 31240 27030 31249
rect 26974 31175 27030 31184
rect 26988 30870 27016 31175
rect 26976 30864 27028 30870
rect 26976 30806 27028 30812
rect 26516 30660 26568 30666
rect 26516 30602 26568 30608
rect 26792 30660 26844 30666
rect 26792 30602 26844 30608
rect 26804 30190 26832 30602
rect 26792 30184 26844 30190
rect 26792 30126 26844 30132
rect 27068 29640 27120 29646
rect 27068 29582 27120 29588
rect 26976 28756 27028 28762
rect 26976 28698 27028 28704
rect 26516 27668 26568 27674
rect 26516 27610 26568 27616
rect 26528 26994 26556 27610
rect 26988 27334 27016 28698
rect 27080 27826 27108 29582
rect 27172 28762 27200 31418
rect 27160 28756 27212 28762
rect 27160 28698 27212 28704
rect 27080 27798 27200 27826
rect 26884 27328 26936 27334
rect 26884 27270 26936 27276
rect 26976 27328 27028 27334
rect 26976 27270 27028 27276
rect 26516 26988 26568 26994
rect 26516 26930 26568 26936
rect 26896 26586 26924 27270
rect 26988 27130 27016 27270
rect 26976 27124 27028 27130
rect 26976 27066 27028 27072
rect 26884 26580 26936 26586
rect 26884 26522 26936 26528
rect 26988 26382 27016 27066
rect 27172 26382 27200 27798
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 27160 26376 27212 26382
rect 27160 26318 27212 26324
rect 27172 25362 27200 26318
rect 27160 25356 27212 25362
rect 27160 25298 27212 25304
rect 26424 24676 26476 24682
rect 26424 24618 26476 24624
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 26240 23180 26292 23186
rect 26240 23122 26292 23128
rect 27172 22778 27200 24142
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 27160 22772 27212 22778
rect 27160 22714 27212 22720
rect 26068 22066 26188 22094
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 25596 3664 25648 3670
rect 25596 3606 25648 3612
rect 25688 3664 25740 3670
rect 25688 3606 25740 3612
rect 25136 3596 25188 3602
rect 25136 3538 25188 3544
rect 25228 3596 25280 3602
rect 25228 3538 25280 3544
rect 25044 2576 25096 2582
rect 25044 2518 25096 2524
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23216 800 23244 2382
rect 24492 2372 24544 2378
rect 24492 2314 24544 2320
rect 24504 800 24532 2314
rect 25148 800 25176 3538
rect 25240 3398 25268 3538
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 26068 3126 26096 22066
rect 26252 22001 26280 22714
rect 27264 22094 27292 35090
rect 27356 34610 27384 35498
rect 27436 34944 27488 34950
rect 27436 34886 27488 34892
rect 27344 34604 27396 34610
rect 27344 34546 27396 34552
rect 27448 33930 27476 34886
rect 27540 34066 27568 35702
rect 27712 35080 27764 35086
rect 27712 35022 27764 35028
rect 27724 34746 27752 35022
rect 27712 34740 27764 34746
rect 27712 34682 27764 34688
rect 27528 34060 27580 34066
rect 27528 34002 27580 34008
rect 27436 33924 27488 33930
rect 27436 33866 27488 33872
rect 27344 33312 27396 33318
rect 27344 33254 27396 33260
rect 27356 32910 27384 33254
rect 27540 33114 27568 34002
rect 27908 33862 27936 36110
rect 28172 35692 28224 35698
rect 28172 35634 28224 35640
rect 28184 35018 28212 35634
rect 28632 35624 28684 35630
rect 28632 35566 28684 35572
rect 28264 35488 28316 35494
rect 28264 35430 28316 35436
rect 28448 35488 28500 35494
rect 28448 35430 28500 35436
rect 28276 35222 28304 35430
rect 28460 35290 28488 35430
rect 28448 35284 28500 35290
rect 28448 35226 28500 35232
rect 28264 35216 28316 35222
rect 28264 35158 28316 35164
rect 28644 35154 28672 35566
rect 29012 35290 29040 36110
rect 29656 36106 29684 37198
rect 29932 36582 29960 37266
rect 29920 36576 29972 36582
rect 29920 36518 29972 36524
rect 29932 36174 29960 36518
rect 29920 36168 29972 36174
rect 29920 36110 29972 36116
rect 29092 36100 29144 36106
rect 29092 36042 29144 36048
rect 29644 36100 29696 36106
rect 29644 36042 29696 36048
rect 29104 35698 29132 36042
rect 29460 36032 29512 36038
rect 29460 35974 29512 35980
rect 29092 35692 29144 35698
rect 29092 35634 29144 35640
rect 29000 35284 29052 35290
rect 29000 35226 29052 35232
rect 28908 35216 28960 35222
rect 28908 35158 28960 35164
rect 28632 35148 28684 35154
rect 28632 35090 28684 35096
rect 28172 35012 28224 35018
rect 28172 34954 28224 34960
rect 28540 35012 28592 35018
rect 28540 34954 28592 34960
rect 27896 33856 27948 33862
rect 27896 33798 27948 33804
rect 27620 33380 27672 33386
rect 27620 33322 27672 33328
rect 27528 33108 27580 33114
rect 27528 33050 27580 33056
rect 27344 32904 27396 32910
rect 27344 32846 27396 32852
rect 27356 31414 27384 32846
rect 27540 32450 27568 33050
rect 27632 32978 27660 33322
rect 27620 32972 27672 32978
rect 27620 32914 27672 32920
rect 27448 32422 27568 32450
rect 27448 31890 27476 32422
rect 27436 31884 27488 31890
rect 27436 31826 27488 31832
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 27724 31482 27752 31690
rect 27712 31476 27764 31482
rect 27712 31418 27764 31424
rect 27344 31408 27396 31414
rect 27344 31350 27396 31356
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27436 30048 27488 30054
rect 27436 29990 27488 29996
rect 27448 29714 27476 29990
rect 27436 29708 27488 29714
rect 27436 29650 27488 29656
rect 27436 29572 27488 29578
rect 27436 29514 27488 29520
rect 27448 29306 27476 29514
rect 27436 29300 27488 29306
rect 27436 29242 27488 29248
rect 27632 28937 27660 31282
rect 27804 30252 27856 30258
rect 27804 30194 27856 30200
rect 27712 30048 27764 30054
rect 27712 29990 27764 29996
rect 27724 29170 27752 29990
rect 27712 29164 27764 29170
rect 27712 29106 27764 29112
rect 27816 29034 27844 30194
rect 27804 29028 27856 29034
rect 27804 28970 27856 28976
rect 27618 28928 27674 28937
rect 27618 28863 27674 28872
rect 27632 27130 27660 28863
rect 27908 27470 27936 33798
rect 28448 33652 28500 33658
rect 28448 33594 28500 33600
rect 28264 32836 28316 32842
rect 28264 32778 28316 32784
rect 28172 32428 28224 32434
rect 28276 32416 28304 32778
rect 28460 32774 28488 33594
rect 28552 33318 28580 34954
rect 28644 34678 28672 35090
rect 28724 34944 28776 34950
rect 28724 34886 28776 34892
rect 28632 34672 28684 34678
rect 28632 34614 28684 34620
rect 28644 34202 28672 34614
rect 28736 34610 28764 34886
rect 28920 34610 28948 35158
rect 29000 35080 29052 35086
rect 29000 35022 29052 35028
rect 28724 34604 28776 34610
rect 28724 34546 28776 34552
rect 28908 34604 28960 34610
rect 28908 34546 28960 34552
rect 28816 34536 28868 34542
rect 28816 34478 28868 34484
rect 28632 34196 28684 34202
rect 28632 34138 28684 34144
rect 28644 33522 28672 34138
rect 28632 33516 28684 33522
rect 28632 33458 28684 33464
rect 28630 33416 28686 33425
rect 28630 33351 28686 33360
rect 28540 33312 28592 33318
rect 28540 33254 28592 33260
rect 28540 32972 28592 32978
rect 28540 32914 28592 32920
rect 28448 32768 28500 32774
rect 28448 32710 28500 32716
rect 28552 32434 28580 32914
rect 28644 32570 28672 33351
rect 28724 33312 28776 33318
rect 28724 33254 28776 33260
rect 28632 32564 28684 32570
rect 28632 32506 28684 32512
rect 28448 32428 28500 32434
rect 28276 32388 28448 32416
rect 28172 32370 28224 32376
rect 28448 32370 28500 32376
rect 28540 32428 28592 32434
rect 28540 32370 28592 32376
rect 28080 32224 28132 32230
rect 28080 32166 28132 32172
rect 28092 31890 28120 32166
rect 28184 32026 28212 32370
rect 28264 32224 28316 32230
rect 28264 32166 28316 32172
rect 28172 32020 28224 32026
rect 28172 31962 28224 31968
rect 28080 31884 28132 31890
rect 28080 31826 28132 31832
rect 28276 31278 28304 32166
rect 28264 31272 28316 31278
rect 28264 31214 28316 31220
rect 28264 30592 28316 30598
rect 28264 30534 28316 30540
rect 27988 29504 28040 29510
rect 27988 29446 28040 29452
rect 28000 29170 28028 29446
rect 27988 29164 28040 29170
rect 27988 29106 28040 29112
rect 27988 29028 28040 29034
rect 27988 28970 28040 28976
rect 27896 27464 27948 27470
rect 27896 27406 27948 27412
rect 27620 27124 27672 27130
rect 27620 27066 27672 27072
rect 27528 26988 27580 26994
rect 27528 26930 27580 26936
rect 27540 26042 27568 26930
rect 27528 26036 27580 26042
rect 27528 25978 27580 25984
rect 27344 24608 27396 24614
rect 27344 24550 27396 24556
rect 27356 24274 27384 24550
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27804 23656 27856 23662
rect 27804 23598 27856 23604
rect 27816 23118 27844 23598
rect 27896 23180 27948 23186
rect 27896 23122 27948 23128
rect 27804 23112 27856 23118
rect 27804 23054 27856 23060
rect 27528 22568 27580 22574
rect 27528 22510 27580 22516
rect 27540 22234 27568 22510
rect 27528 22228 27580 22234
rect 27528 22170 27580 22176
rect 27264 22066 27476 22094
rect 26976 22024 27028 22030
rect 26238 21992 26294 22001
rect 26976 21966 27028 21972
rect 26238 21927 26294 21936
rect 26988 21434 27016 21966
rect 26896 21406 27016 21434
rect 27344 21412 27396 21418
rect 26896 20466 26924 21406
rect 27344 21354 27396 21360
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26884 20460 26936 20466
rect 26884 20402 26936 20408
rect 26896 19718 26924 20402
rect 26988 19854 27016 21286
rect 27160 20800 27212 20806
rect 27160 20742 27212 20748
rect 27172 20398 27200 20742
rect 27356 20534 27384 21354
rect 27344 20528 27396 20534
rect 27344 20470 27396 20476
rect 27160 20392 27212 20398
rect 27160 20334 27212 20340
rect 27356 20058 27384 20470
rect 27344 20052 27396 20058
rect 27344 19994 27396 20000
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 26884 19712 26936 19718
rect 26884 19654 26936 19660
rect 27252 18760 27304 18766
rect 27252 18702 27304 18708
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26148 17876 26200 17882
rect 26148 17818 26200 17824
rect 26160 17270 26188 17818
rect 26792 17604 26844 17610
rect 26792 17546 26844 17552
rect 26148 17264 26200 17270
rect 26148 17206 26200 17212
rect 26804 16998 26832 17546
rect 26988 17338 27016 18158
rect 27172 17882 27200 18226
rect 27264 18222 27292 18702
rect 27252 18216 27304 18222
rect 27252 18158 27304 18164
rect 27160 17876 27212 17882
rect 27160 17818 27212 17824
rect 26976 17332 27028 17338
rect 26976 17274 27028 17280
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 26804 16590 26832 16934
rect 26988 16658 27016 17274
rect 27068 17128 27120 17134
rect 27068 17070 27120 17076
rect 27080 16794 27108 17070
rect 27068 16788 27120 16794
rect 27068 16730 27120 16736
rect 26976 16652 27028 16658
rect 26976 16594 27028 16600
rect 26792 16584 26844 16590
rect 26792 16526 26844 16532
rect 27448 6914 27476 22066
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27816 21554 27844 21966
rect 27908 21690 27936 23122
rect 28000 22094 28028 28970
rect 28276 28966 28304 30534
rect 28460 30394 28488 32370
rect 28736 31890 28764 33254
rect 28828 33046 28856 34478
rect 28920 33590 28948 34546
rect 28908 33584 28960 33590
rect 28908 33526 28960 33532
rect 28816 33040 28868 33046
rect 28816 32982 28868 32988
rect 29012 32434 29040 35022
rect 29104 33658 29132 35634
rect 29472 34610 29500 35974
rect 29828 35012 29880 35018
rect 29828 34954 29880 34960
rect 29460 34604 29512 34610
rect 29460 34546 29512 34552
rect 29644 33924 29696 33930
rect 29644 33866 29696 33872
rect 29092 33652 29144 33658
rect 29092 33594 29144 33600
rect 29656 33114 29684 33866
rect 29736 33856 29788 33862
rect 29736 33798 29788 33804
rect 29644 33108 29696 33114
rect 29644 33050 29696 33056
rect 29552 32904 29604 32910
rect 29552 32846 29604 32852
rect 29564 32774 29592 32846
rect 29552 32768 29604 32774
rect 29552 32710 29604 32716
rect 29000 32428 29052 32434
rect 29000 32370 29052 32376
rect 28908 32020 28960 32026
rect 28908 31962 28960 31968
rect 28724 31884 28776 31890
rect 28724 31826 28776 31832
rect 28920 31482 28948 31962
rect 29012 31754 29040 32370
rect 29368 32020 29420 32026
rect 29368 31962 29420 31968
rect 29380 31822 29408 31962
rect 29564 31822 29592 32710
rect 29368 31816 29420 31822
rect 29368 31758 29420 31764
rect 29552 31816 29604 31822
rect 29552 31758 29604 31764
rect 29012 31726 29132 31754
rect 28908 31476 28960 31482
rect 28908 31418 28960 31424
rect 28632 31340 28684 31346
rect 28632 31282 28684 31288
rect 28816 31340 28868 31346
rect 28816 31282 28868 31288
rect 28540 30728 28592 30734
rect 28540 30670 28592 30676
rect 28448 30388 28500 30394
rect 28448 30330 28500 30336
rect 28356 29572 28408 29578
rect 28356 29514 28408 29520
rect 28264 28960 28316 28966
rect 28264 28902 28316 28908
rect 28276 28558 28304 28902
rect 28368 28762 28396 29514
rect 28356 28756 28408 28762
rect 28356 28698 28408 28704
rect 28552 28626 28580 30670
rect 28540 28620 28592 28626
rect 28540 28562 28592 28568
rect 28264 28552 28316 28558
rect 28264 28494 28316 28500
rect 28264 27328 28316 27334
rect 28264 27270 28316 27276
rect 28276 26994 28304 27270
rect 28264 26988 28316 26994
rect 28264 26930 28316 26936
rect 28552 25838 28580 28562
rect 28540 25832 28592 25838
rect 28540 25774 28592 25780
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 28276 23866 28304 24754
rect 28356 24608 28408 24614
rect 28356 24550 28408 24556
rect 28264 23860 28316 23866
rect 28264 23802 28316 23808
rect 28080 23180 28132 23186
rect 28080 23122 28132 23128
rect 28092 22710 28120 23122
rect 28080 22704 28132 22710
rect 28080 22646 28132 22652
rect 28000 22066 28120 22094
rect 27896 21684 27948 21690
rect 27896 21626 27948 21632
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27804 21140 27856 21146
rect 27804 21082 27856 21088
rect 27816 20942 27844 21082
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 27908 20874 27936 21490
rect 27988 21344 28040 21350
rect 27988 21286 28040 21292
rect 27896 20868 27948 20874
rect 27896 20810 27948 20816
rect 27908 19854 27936 20810
rect 28000 20534 28028 21286
rect 27988 20528 28040 20534
rect 27988 20470 28040 20476
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 27712 18692 27764 18698
rect 27712 18634 27764 18640
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27632 16794 27660 17478
rect 27724 17338 27752 18634
rect 27896 18148 27948 18154
rect 27896 18090 27948 18096
rect 27804 18080 27856 18086
rect 27804 18022 27856 18028
rect 27816 17746 27844 18022
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 27712 17332 27764 17338
rect 27712 17274 27764 17280
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27908 16590 27936 18090
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 28092 6914 28120 22066
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28184 21146 28212 21422
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 28184 20874 28212 20946
rect 28172 20868 28224 20874
rect 28172 20810 28224 20816
rect 28276 19378 28304 23802
rect 28368 23798 28396 24550
rect 28356 23792 28408 23798
rect 28356 23734 28408 23740
rect 28448 23112 28500 23118
rect 28448 23054 28500 23060
rect 28460 22778 28488 23054
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 28448 21684 28500 21690
rect 28448 21626 28500 21632
rect 28460 21593 28488 21626
rect 28446 21584 28502 21593
rect 28356 21548 28408 21554
rect 28446 21519 28502 21528
rect 28356 21490 28408 21496
rect 28368 21010 28396 21490
rect 28448 21140 28500 21146
rect 28448 21082 28500 21088
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 28368 19854 28396 20946
rect 28460 20942 28488 21082
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28356 19848 28408 19854
rect 28356 19790 28408 19796
rect 28460 19718 28488 20878
rect 28448 19712 28500 19718
rect 28448 19654 28500 19660
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28552 8838 28580 25774
rect 28540 8832 28592 8838
rect 28540 8774 28592 8780
rect 27356 6886 27476 6914
rect 28000 6886 28120 6914
rect 27160 4208 27212 4214
rect 27160 4150 27212 4156
rect 27172 4049 27200 4150
rect 26974 4040 27030 4049
rect 26974 3975 27030 3984
rect 27158 4040 27214 4049
rect 27158 3975 27214 3984
rect 26620 3466 26832 3482
rect 26608 3460 26844 3466
rect 26660 3454 26792 3460
rect 26608 3402 26660 3408
rect 26792 3402 26844 3408
rect 26884 3392 26936 3398
rect 26884 3334 26936 3340
rect 26896 3126 26924 3334
rect 26056 3120 26108 3126
rect 26056 3062 26108 3068
rect 26884 3120 26936 3126
rect 26884 3062 26936 3068
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 26436 800 26464 2994
rect 26988 2446 27016 3975
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 27080 3074 27108 3130
rect 27080 3046 27200 3074
rect 27172 2990 27200 3046
rect 27160 2984 27212 2990
rect 27160 2926 27212 2932
rect 26976 2440 27028 2446
rect 26976 2382 27028 2388
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 27080 800 27108 2314
rect 27356 2310 27384 6886
rect 27436 3528 27488 3534
rect 27436 3470 27488 3476
rect 27448 2650 27476 3470
rect 27436 2644 27488 2650
rect 27436 2586 27488 2592
rect 28000 2514 28028 6886
rect 28080 4072 28132 4078
rect 28080 4014 28132 4020
rect 28092 3126 28120 4014
rect 28644 3126 28672 31282
rect 28828 30394 28856 31282
rect 28816 30388 28868 30394
rect 28816 30330 28868 30336
rect 28828 29170 28856 30330
rect 28920 30326 28948 31418
rect 29000 31340 29052 31346
rect 29000 31282 29052 31288
rect 29012 30734 29040 31282
rect 29000 30728 29052 30734
rect 29000 30670 29052 30676
rect 28908 30320 28960 30326
rect 28908 30262 28960 30268
rect 29012 30258 29040 30670
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 29012 29850 29040 30194
rect 29104 30122 29132 31726
rect 29748 31686 29776 33798
rect 29736 31680 29788 31686
rect 29736 31622 29788 31628
rect 29748 30394 29776 31622
rect 29736 30388 29788 30394
rect 29736 30330 29788 30336
rect 29460 30252 29512 30258
rect 29460 30194 29512 30200
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 29092 30116 29144 30122
rect 29092 30058 29144 30064
rect 29000 29844 29052 29850
rect 29000 29786 29052 29792
rect 28816 29164 28868 29170
rect 28816 29106 28868 29112
rect 29012 29102 29040 29786
rect 29000 29096 29052 29102
rect 29000 29038 29052 29044
rect 29472 28490 29500 30194
rect 29656 29034 29684 30194
rect 29840 30138 29868 34954
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29932 30258 29960 34546
rect 30010 32328 30066 32337
rect 30010 32263 30066 32272
rect 30024 31958 30052 32263
rect 30012 31952 30064 31958
rect 30012 31894 30064 31900
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 30012 30184 30064 30190
rect 29840 30110 29960 30138
rect 30012 30126 30064 30132
rect 29932 29850 29960 30110
rect 29920 29844 29972 29850
rect 29920 29786 29972 29792
rect 30024 29646 30052 30126
rect 29736 29640 29788 29646
rect 29736 29582 29788 29588
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 29748 29306 29776 29582
rect 30024 29510 30052 29582
rect 30012 29504 30064 29510
rect 30012 29446 30064 29452
rect 29736 29300 29788 29306
rect 29736 29242 29788 29248
rect 29644 29028 29696 29034
rect 29644 28970 29696 28976
rect 30012 29028 30064 29034
rect 30012 28970 30064 28976
rect 29460 28484 29512 28490
rect 29460 28426 29512 28432
rect 29472 28150 29500 28426
rect 29552 28416 29604 28422
rect 29552 28358 29604 28364
rect 29564 28150 29592 28358
rect 29460 28144 29512 28150
rect 29460 28086 29512 28092
rect 29552 28144 29604 28150
rect 29552 28086 29604 28092
rect 28908 27532 28960 27538
rect 28908 27474 28960 27480
rect 28920 26586 28948 27474
rect 28908 26580 28960 26586
rect 28908 26522 28960 26528
rect 29472 26518 29500 28086
rect 30024 28082 30052 28970
rect 30012 28076 30064 28082
rect 30012 28018 30064 28024
rect 30012 27872 30064 27878
rect 30012 27814 30064 27820
rect 29736 26920 29788 26926
rect 29736 26862 29788 26868
rect 29460 26512 29512 26518
rect 29460 26454 29512 26460
rect 29092 26308 29144 26314
rect 29092 26250 29144 26256
rect 29104 26042 29132 26250
rect 29092 26036 29144 26042
rect 29092 25978 29144 25984
rect 29472 25974 29500 26454
rect 29748 26382 29776 26862
rect 29920 26512 29972 26518
rect 29920 26454 29972 26460
rect 29736 26376 29788 26382
rect 29736 26318 29788 26324
rect 29460 25968 29512 25974
rect 29460 25910 29512 25916
rect 29932 25786 29960 26454
rect 30024 25974 30052 27814
rect 30116 26908 30144 47126
rect 30760 47122 30788 49286
rect 30902 49200 31014 49286
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49200 40030 50000
rect 40562 49200 40674 50000
rect 41206 49200 41318 50000
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 43782 49200 43894 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49200 46470 50000
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 30748 47116 30800 47122
rect 30748 47058 30800 47064
rect 30840 47048 30892 47054
rect 30840 46990 30892 46996
rect 30656 37868 30708 37874
rect 30656 37810 30708 37816
rect 30668 36786 30696 37810
rect 30656 36780 30708 36786
rect 30656 36722 30708 36728
rect 30748 36576 30800 36582
rect 30748 36518 30800 36524
rect 30760 35766 30788 36518
rect 30748 35760 30800 35766
rect 30748 35702 30800 35708
rect 30748 35624 30800 35630
rect 30748 35566 30800 35572
rect 30564 35488 30616 35494
rect 30564 35430 30616 35436
rect 30576 35154 30604 35430
rect 30760 35290 30788 35566
rect 30748 35284 30800 35290
rect 30748 35226 30800 35232
rect 30564 35148 30616 35154
rect 30564 35090 30616 35096
rect 30288 35080 30340 35086
rect 30288 35022 30340 35028
rect 30300 34746 30328 35022
rect 30288 34740 30340 34746
rect 30288 34682 30340 34688
rect 30576 34678 30604 35090
rect 30564 34672 30616 34678
rect 30564 34614 30616 34620
rect 30380 34400 30432 34406
rect 30380 34342 30432 34348
rect 30392 33930 30420 34342
rect 30852 33998 30880 46990
rect 32232 46594 32260 49200
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 34796 47184 34848 47190
rect 34796 47126 34848 47132
rect 34612 46980 34664 46986
rect 34612 46922 34664 46928
rect 32232 46566 32352 46594
rect 32220 46504 32272 46510
rect 32220 46446 32272 46452
rect 32232 46170 32260 46446
rect 32324 46442 32352 46566
rect 32404 46504 32456 46510
rect 32404 46446 32456 46452
rect 32312 46436 32364 46442
rect 32312 46378 32364 46384
rect 32220 46164 32272 46170
rect 32220 46106 32272 46112
rect 32416 45626 32444 46446
rect 32404 45620 32456 45626
rect 32404 45562 32456 45568
rect 31024 35828 31076 35834
rect 31024 35770 31076 35776
rect 30932 35148 30984 35154
rect 30932 35090 30984 35096
rect 30472 33992 30524 33998
rect 30472 33934 30524 33940
rect 30840 33992 30892 33998
rect 30840 33934 30892 33940
rect 30380 33924 30432 33930
rect 30380 33866 30432 33872
rect 30392 32586 30420 33866
rect 30484 33522 30512 33934
rect 30472 33516 30524 33522
rect 30472 33458 30524 33464
rect 30840 33448 30892 33454
rect 30840 33390 30892 33396
rect 30564 32836 30616 32842
rect 30564 32778 30616 32784
rect 30300 32558 30420 32586
rect 30196 32224 30248 32230
rect 30196 32166 30248 32172
rect 30208 32026 30236 32166
rect 30196 32020 30248 32026
rect 30196 31962 30248 31968
rect 30208 30938 30236 31962
rect 30300 31770 30328 32558
rect 30472 32292 30524 32298
rect 30472 32234 30524 32240
rect 30484 32026 30512 32234
rect 30576 32230 30604 32778
rect 30656 32768 30708 32774
rect 30656 32710 30708 32716
rect 30564 32224 30616 32230
rect 30564 32166 30616 32172
rect 30472 32020 30524 32026
rect 30472 31962 30524 31968
rect 30472 31816 30524 31822
rect 30300 31742 30420 31770
rect 30472 31758 30524 31764
rect 30196 30932 30248 30938
rect 30196 30874 30248 30880
rect 30288 30796 30340 30802
rect 30288 30738 30340 30744
rect 30300 30666 30328 30738
rect 30392 30682 30420 31742
rect 30484 31278 30512 31758
rect 30472 31272 30524 31278
rect 30472 31214 30524 31220
rect 30668 30734 30696 32710
rect 30852 32366 30880 33390
rect 30840 32360 30892 32366
rect 30840 32302 30892 32308
rect 30748 31952 30800 31958
rect 30746 31920 30748 31929
rect 30800 31920 30802 31929
rect 30746 31855 30802 31864
rect 30760 31686 30788 31855
rect 30748 31680 30800 31686
rect 30748 31622 30800 31628
rect 30852 31346 30880 32302
rect 30944 31754 30972 35090
rect 31036 35086 31064 35770
rect 31024 35080 31076 35086
rect 31024 35022 31076 35028
rect 31036 34082 31064 35022
rect 31036 34054 31248 34082
rect 31024 33516 31076 33522
rect 31024 33458 31076 33464
rect 31036 32774 31064 33458
rect 31116 32972 31168 32978
rect 31116 32914 31168 32920
rect 31024 32768 31076 32774
rect 31024 32710 31076 32716
rect 31024 32360 31076 32366
rect 31024 32302 31076 32308
rect 31036 31890 31064 32302
rect 31128 31890 31156 32914
rect 31024 31884 31076 31890
rect 31024 31826 31076 31832
rect 31116 31884 31168 31890
rect 31116 31826 31168 31832
rect 30944 31726 31064 31754
rect 30840 31340 30892 31346
rect 30840 31282 30892 31288
rect 30852 30938 30880 31282
rect 30840 30932 30892 30938
rect 30840 30874 30892 30880
rect 30656 30728 30708 30734
rect 30288 30660 30340 30666
rect 30392 30654 30604 30682
rect 30656 30670 30708 30676
rect 30288 30602 30340 30608
rect 30300 30190 30328 30602
rect 30380 30592 30432 30598
rect 30380 30534 30432 30540
rect 30288 30184 30340 30190
rect 30288 30126 30340 30132
rect 30196 29844 30248 29850
rect 30196 29786 30248 29792
rect 30208 28694 30236 29786
rect 30288 29164 30340 29170
rect 30288 29106 30340 29112
rect 30196 28688 30248 28694
rect 30196 28630 30248 28636
rect 30300 28490 30328 29106
rect 30392 28558 30420 30534
rect 30576 29170 30604 30654
rect 30668 30054 30696 30670
rect 30852 30258 30880 30874
rect 30840 30252 30892 30258
rect 30840 30194 30892 30200
rect 30656 30048 30708 30054
rect 30656 29990 30708 29996
rect 30564 29164 30616 29170
rect 30564 29106 30616 29112
rect 30748 29164 30800 29170
rect 30748 29106 30800 29112
rect 30380 28552 30432 28558
rect 30380 28494 30432 28500
rect 30288 28484 30340 28490
rect 30288 28426 30340 28432
rect 30196 28076 30248 28082
rect 30196 28018 30248 28024
rect 30208 27470 30236 28018
rect 30380 27668 30432 27674
rect 30380 27610 30432 27616
rect 30196 27464 30248 27470
rect 30196 27406 30248 27412
rect 30392 26994 30420 27610
rect 30576 27146 30604 29106
rect 30656 29028 30708 29034
rect 30656 28970 30708 28976
rect 30668 28150 30696 28970
rect 30760 28762 30788 29106
rect 30748 28756 30800 28762
rect 30748 28698 30800 28704
rect 30656 28144 30708 28150
rect 30656 28086 30708 28092
rect 30484 27130 30604 27146
rect 30472 27124 30604 27130
rect 30524 27118 30604 27124
rect 30472 27066 30524 27072
rect 30576 26994 30604 27118
rect 30668 27062 30696 28086
rect 30656 27056 30708 27062
rect 30656 26998 30708 27004
rect 30380 26988 30432 26994
rect 30380 26930 30432 26936
rect 30564 26988 30616 26994
rect 30564 26930 30616 26936
rect 30472 26920 30524 26926
rect 30116 26880 30236 26908
rect 30104 26240 30156 26246
rect 30104 26182 30156 26188
rect 30012 25968 30064 25974
rect 30012 25910 30064 25916
rect 30116 25906 30144 26182
rect 30104 25900 30156 25906
rect 30104 25842 30156 25848
rect 29932 25758 30052 25786
rect 29920 25696 29972 25702
rect 29920 25638 29972 25644
rect 29932 25362 29960 25638
rect 29920 25356 29972 25362
rect 29920 25298 29972 25304
rect 28816 22704 28868 22710
rect 28816 22646 28868 22652
rect 28828 21894 28856 22646
rect 28908 22500 28960 22506
rect 28908 22442 28960 22448
rect 28816 21888 28868 21894
rect 28816 21830 28868 21836
rect 28816 21548 28868 21554
rect 28816 21490 28868 21496
rect 28828 20058 28856 21490
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28920 19938 28948 22442
rect 29368 22024 29420 22030
rect 29736 22024 29788 22030
rect 29420 21984 29736 22012
rect 29368 21966 29420 21972
rect 29736 21966 29788 21972
rect 29000 21548 29052 21554
rect 29000 21490 29052 21496
rect 29012 20806 29040 21490
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 29380 20466 29408 21966
rect 29460 21888 29512 21894
rect 29460 21830 29512 21836
rect 29472 21554 29500 21830
rect 29460 21548 29512 21554
rect 29460 21490 29512 21496
rect 29368 20460 29420 20466
rect 29368 20402 29420 20408
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 28736 19910 28948 19938
rect 29472 19922 29500 20198
rect 30024 20058 30052 25758
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 30116 21146 30144 21422
rect 30104 21140 30156 21146
rect 30104 21082 30156 21088
rect 30208 20806 30236 26880
rect 30472 26862 30524 26868
rect 30380 26444 30432 26450
rect 30380 26386 30432 26392
rect 30288 25832 30340 25838
rect 30288 25774 30340 25780
rect 30300 24818 30328 25774
rect 30392 25498 30420 26386
rect 30380 25492 30432 25498
rect 30380 25434 30432 25440
rect 30288 24812 30340 24818
rect 30288 24754 30340 24760
rect 30196 20800 30248 20806
rect 30196 20742 30248 20748
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 29460 19916 29512 19922
rect 28736 18306 28764 19910
rect 29460 19858 29512 19864
rect 28908 19780 28960 19786
rect 28908 19722 28960 19728
rect 28920 19514 28948 19722
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 30300 19446 30328 24754
rect 30380 21888 30432 21894
rect 30380 21830 30432 21836
rect 30392 21622 30420 21830
rect 30380 21616 30432 21622
rect 30380 21558 30432 21564
rect 29000 19440 29052 19446
rect 29000 19382 29052 19388
rect 30288 19440 30340 19446
rect 30288 19382 30340 19388
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 28816 18352 28868 18358
rect 28736 18300 28816 18306
rect 28736 18294 28868 18300
rect 28736 18278 28856 18294
rect 28736 17882 28764 18278
rect 28816 18080 28868 18086
rect 28816 18022 28868 18028
rect 28724 17876 28776 17882
rect 28724 17818 28776 17824
rect 28828 17610 28856 18022
rect 28816 17604 28868 17610
rect 28816 17546 28868 17552
rect 28920 6914 28948 19314
rect 29012 18290 29040 19382
rect 30380 18352 30432 18358
rect 30380 18294 30432 18300
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 29012 17678 29040 18226
rect 30392 17678 30420 18294
rect 29000 17672 29052 17678
rect 29000 17614 29052 17620
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 29644 17536 29696 17542
rect 29644 17478 29696 17484
rect 29656 17270 29684 17478
rect 29644 17264 29696 17270
rect 29644 17206 29696 17212
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30392 13394 30420 14214
rect 30380 13388 30432 13394
rect 30380 13330 30432 13336
rect 30484 12646 30512 26862
rect 30932 25220 30984 25226
rect 30932 25162 30984 25168
rect 30944 24818 30972 25162
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30932 18964 30984 18970
rect 30932 18906 30984 18912
rect 30944 18766 30972 18906
rect 30932 18760 30984 18766
rect 30932 18702 30984 18708
rect 30656 18284 30708 18290
rect 30656 18226 30708 18232
rect 30668 17678 30696 18226
rect 30656 17672 30708 17678
rect 30656 17614 30708 17620
rect 30564 14272 30616 14278
rect 30564 14214 30616 14220
rect 30576 13394 30604 14214
rect 30564 13388 30616 13394
rect 30564 13330 30616 13336
rect 30472 12640 30524 12646
rect 30472 12582 30524 12588
rect 28828 6886 28948 6914
rect 28828 4010 28856 6886
rect 28816 4004 28868 4010
rect 28816 3946 28868 3952
rect 28080 3120 28132 3126
rect 28080 3062 28132 3068
rect 28632 3120 28684 3126
rect 28632 3062 28684 3068
rect 30668 2854 30696 17614
rect 30944 17610 30972 18702
rect 30932 17604 30984 17610
rect 30932 17546 30984 17552
rect 31036 4146 31064 31726
rect 31220 31414 31248 34054
rect 31300 33856 31352 33862
rect 31300 33798 31352 33804
rect 31312 32434 31340 33798
rect 31576 33380 31628 33386
rect 31576 33322 31628 33328
rect 31392 32836 31444 32842
rect 31392 32778 31444 32784
rect 31404 32570 31432 32778
rect 31392 32564 31444 32570
rect 31392 32506 31444 32512
rect 31588 32434 31616 33322
rect 33692 32836 33744 32842
rect 33692 32778 33744 32784
rect 31668 32768 31720 32774
rect 31668 32710 31720 32716
rect 31680 32450 31708 32710
rect 33704 32570 33732 32778
rect 33692 32564 33744 32570
rect 33692 32506 33744 32512
rect 31680 32434 31800 32450
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 31484 32428 31536 32434
rect 31484 32370 31536 32376
rect 31576 32428 31628 32434
rect 31680 32428 31812 32434
rect 31680 32422 31760 32428
rect 31576 32370 31628 32376
rect 31760 32370 31812 32376
rect 33692 32428 33744 32434
rect 33692 32370 33744 32376
rect 31496 32337 31524 32370
rect 32680 32360 32732 32366
rect 31482 32328 31538 32337
rect 31300 32292 31352 32298
rect 32680 32302 32732 32308
rect 31482 32263 31538 32272
rect 31300 32234 31352 32240
rect 31312 31822 31340 32234
rect 31300 31816 31352 31822
rect 31496 31804 31524 32263
rect 31576 31816 31628 31822
rect 31496 31776 31576 31804
rect 31300 31758 31352 31764
rect 31576 31758 31628 31764
rect 32404 31680 32456 31686
rect 32404 31622 32456 31628
rect 31208 31408 31260 31414
rect 31208 31350 31260 31356
rect 32416 31346 32444 31622
rect 32692 31346 32720 32302
rect 33140 31884 33192 31890
rect 33140 31826 33192 31832
rect 33152 31482 33180 31826
rect 33140 31476 33192 31482
rect 33140 31418 33192 31424
rect 33704 31346 33732 32370
rect 34152 32360 34204 32366
rect 34152 32302 34204 32308
rect 34164 31958 34192 32302
rect 34152 31952 34204 31958
rect 34152 31894 34204 31900
rect 33784 31816 33836 31822
rect 33784 31758 33836 31764
rect 33796 31482 33824 31758
rect 33784 31476 33836 31482
rect 33784 31418 33836 31424
rect 32404 31340 32456 31346
rect 32404 31282 32456 31288
rect 32588 31340 32640 31346
rect 32588 31282 32640 31288
rect 32680 31340 32732 31346
rect 32680 31282 32732 31288
rect 32956 31340 33008 31346
rect 32956 31282 33008 31288
rect 33692 31340 33744 31346
rect 33692 31282 33744 31288
rect 31116 31272 31168 31278
rect 31116 31214 31168 31220
rect 32496 31272 32548 31278
rect 32496 31214 32548 31220
rect 31128 27606 31156 31214
rect 32404 30728 32456 30734
rect 32404 30670 32456 30676
rect 31300 30184 31352 30190
rect 31300 30126 31352 30132
rect 31312 29850 31340 30126
rect 32416 30122 32444 30670
rect 32404 30116 32456 30122
rect 32404 30058 32456 30064
rect 31392 30048 31444 30054
rect 31392 29990 31444 29996
rect 31760 30048 31812 30054
rect 31760 29990 31812 29996
rect 31300 29844 31352 29850
rect 31300 29786 31352 29792
rect 31404 27606 31432 29990
rect 31484 28076 31536 28082
rect 31484 28018 31536 28024
rect 31116 27600 31168 27606
rect 31116 27542 31168 27548
rect 31392 27600 31444 27606
rect 31392 27542 31444 27548
rect 31208 27532 31260 27538
rect 31208 27474 31260 27480
rect 31220 27062 31248 27474
rect 31392 27328 31444 27334
rect 31392 27270 31444 27276
rect 31208 27056 31260 27062
rect 31208 26998 31260 27004
rect 31404 26994 31432 27270
rect 31496 27130 31524 28018
rect 31772 27470 31800 29990
rect 32128 29572 32180 29578
rect 32128 29514 32180 29520
rect 32140 29306 32168 29514
rect 32128 29300 32180 29306
rect 32128 29242 32180 29248
rect 31760 27464 31812 27470
rect 31760 27406 31812 27412
rect 31944 27464 31996 27470
rect 31944 27406 31996 27412
rect 32312 27464 32364 27470
rect 32312 27406 32364 27412
rect 31484 27124 31536 27130
rect 31484 27066 31536 27072
rect 31392 26988 31444 26994
rect 31392 26930 31444 26936
rect 31576 26988 31628 26994
rect 31576 26930 31628 26936
rect 31300 26784 31352 26790
rect 31300 26726 31352 26732
rect 31312 26450 31340 26726
rect 31300 26444 31352 26450
rect 31300 26386 31352 26392
rect 31588 26314 31616 26930
rect 31956 26926 31984 27406
rect 32324 26994 32352 27406
rect 32312 26988 32364 26994
rect 32312 26930 32364 26936
rect 31944 26920 31996 26926
rect 31944 26862 31996 26868
rect 32324 26586 32352 26930
rect 32312 26580 32364 26586
rect 32312 26522 32364 26528
rect 31576 26308 31628 26314
rect 31576 26250 31628 26256
rect 31760 26308 31812 26314
rect 31760 26250 31812 26256
rect 31588 25498 31616 26250
rect 31772 26042 31800 26250
rect 31760 26036 31812 26042
rect 31760 25978 31812 25984
rect 31576 25492 31628 25498
rect 31576 25434 31628 25440
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31220 21486 31248 21966
rect 32404 21956 32456 21962
rect 32404 21898 32456 21904
rect 31208 21480 31260 21486
rect 31208 21422 31260 21428
rect 31116 21004 31168 21010
rect 31116 20946 31168 20952
rect 31128 20874 31156 20946
rect 31220 20942 31248 21422
rect 32312 21412 32364 21418
rect 32312 21354 32364 21360
rect 32220 21072 32272 21078
rect 32220 21014 32272 21020
rect 31576 21004 31628 21010
rect 31576 20946 31628 20952
rect 31208 20936 31260 20942
rect 31208 20878 31260 20884
rect 31588 20874 31616 20946
rect 32232 20874 32260 21014
rect 32324 20942 32352 21354
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 31116 20868 31168 20874
rect 31116 20810 31168 20816
rect 31576 20868 31628 20874
rect 31576 20810 31628 20816
rect 32220 20868 32272 20874
rect 32220 20810 32272 20816
rect 31300 19984 31352 19990
rect 31300 19926 31352 19932
rect 31116 18896 31168 18902
rect 31116 18838 31168 18844
rect 31128 18766 31156 18838
rect 31312 18766 31340 19926
rect 31392 19780 31444 19786
rect 31392 19722 31444 19728
rect 31116 18760 31168 18766
rect 31116 18702 31168 18708
rect 31300 18760 31352 18766
rect 31300 18702 31352 18708
rect 31128 17678 31156 18702
rect 31208 18624 31260 18630
rect 31208 18566 31260 18572
rect 31220 18358 31248 18566
rect 31300 18420 31352 18426
rect 31300 18362 31352 18368
rect 31208 18352 31260 18358
rect 31208 18294 31260 18300
rect 31312 18222 31340 18362
rect 31300 18216 31352 18222
rect 31300 18158 31352 18164
rect 31312 17882 31340 18158
rect 31300 17876 31352 17882
rect 31300 17818 31352 17824
rect 31116 17672 31168 17678
rect 31116 17614 31168 17620
rect 31300 17672 31352 17678
rect 31300 17614 31352 17620
rect 31024 4140 31076 4146
rect 31024 4082 31076 4088
rect 31128 4078 31156 17614
rect 31116 4072 31168 4078
rect 31116 4014 31168 4020
rect 30932 3596 30984 3602
rect 30932 3538 30984 3544
rect 30656 2848 30708 2854
rect 30656 2790 30708 2796
rect 27988 2508 28040 2514
rect 27988 2450 28040 2456
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 27344 2304 27396 2310
rect 27344 2246 27396 2252
rect 28368 800 28396 2382
rect 29656 800 29684 2382
rect 29736 2304 29788 2310
rect 29736 2246 29788 2252
rect 29748 1902 29776 2246
rect 29736 1896 29788 1902
rect 29736 1838 29788 1844
rect 30944 800 30972 3538
rect 31312 3534 31340 17614
rect 31404 12434 31432 19722
rect 31484 18964 31536 18970
rect 31484 18906 31536 18912
rect 31496 18766 31524 18906
rect 31484 18760 31536 18766
rect 31484 18702 31536 18708
rect 31588 18578 31616 20810
rect 32218 20632 32274 20641
rect 32218 20567 32220 20576
rect 32272 20567 32274 20576
rect 32220 20538 32272 20544
rect 32220 19984 32272 19990
rect 32220 19926 32272 19932
rect 32232 19786 32260 19926
rect 32324 19854 32352 20878
rect 32416 20602 32444 21898
rect 32404 20596 32456 20602
rect 32404 20538 32456 20544
rect 32312 19848 32364 19854
rect 32312 19790 32364 19796
rect 32220 19780 32272 19786
rect 32220 19722 32272 19728
rect 31668 18896 31720 18902
rect 31668 18838 31720 18844
rect 31680 18698 31708 18838
rect 32324 18748 32352 19790
rect 32404 18760 32456 18766
rect 32324 18720 32404 18748
rect 31668 18692 31720 18698
rect 31668 18634 31720 18640
rect 32324 18630 32352 18720
rect 32404 18702 32456 18708
rect 32312 18624 32364 18630
rect 31588 18550 31708 18578
rect 32312 18566 32364 18572
rect 31484 18420 31536 18426
rect 31484 18362 31536 18368
rect 31496 18086 31524 18362
rect 31576 18284 31628 18290
rect 31576 18226 31628 18232
rect 31484 18080 31536 18086
rect 31484 18022 31536 18028
rect 31588 17746 31616 18226
rect 31576 17740 31628 17746
rect 31576 17682 31628 17688
rect 31484 17672 31536 17678
rect 31484 17614 31536 17620
rect 31496 17338 31524 17614
rect 31484 17332 31536 17338
rect 31484 17274 31536 17280
rect 31588 17218 31616 17682
rect 31496 17202 31616 17218
rect 31484 17196 31616 17202
rect 31536 17190 31616 17196
rect 31484 17138 31536 17144
rect 31404 12406 31524 12434
rect 31300 3528 31352 3534
rect 31300 3470 31352 3476
rect 31496 3398 31524 12406
rect 31680 6914 31708 18550
rect 32312 18080 32364 18086
rect 32312 18022 32364 18028
rect 32324 17678 32352 18022
rect 32312 17672 32364 17678
rect 32312 17614 32364 17620
rect 32220 13252 32272 13258
rect 32220 13194 32272 13200
rect 31588 6886 31708 6914
rect 31588 4146 31616 6886
rect 31576 4140 31628 4146
rect 31576 4082 31628 4088
rect 32232 3602 32260 13194
rect 32220 3596 32272 3602
rect 32220 3538 32272 3544
rect 31484 3392 31536 3398
rect 31484 3334 31536 3340
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 32232 800 32260 2926
rect 32508 2310 32536 31214
rect 32600 30870 32628 31282
rect 32588 30864 32640 30870
rect 32588 30806 32640 30812
rect 32968 30734 32996 31282
rect 32680 30728 32732 30734
rect 32680 30670 32732 30676
rect 32956 30728 33008 30734
rect 32956 30670 33008 30676
rect 32692 30054 32720 30670
rect 33140 30592 33192 30598
rect 33140 30534 33192 30540
rect 33152 30326 33180 30534
rect 33140 30320 33192 30326
rect 33140 30262 33192 30268
rect 32864 30184 32916 30190
rect 32864 30126 32916 30132
rect 32680 30048 32732 30054
rect 32680 29990 32732 29996
rect 32876 29714 32904 30126
rect 32864 29708 32916 29714
rect 32864 29650 32916 29656
rect 33704 29646 33732 31282
rect 33784 30320 33836 30326
rect 33784 30262 33836 30268
rect 33796 29850 33824 30262
rect 33784 29844 33836 29850
rect 33784 29786 33836 29792
rect 33692 29640 33744 29646
rect 33692 29582 33744 29588
rect 33704 29170 33732 29582
rect 33692 29164 33744 29170
rect 33692 29106 33744 29112
rect 34520 22432 34572 22438
rect 34520 22374 34572 22380
rect 34532 21690 34560 22374
rect 34520 21684 34572 21690
rect 34520 21626 34572 21632
rect 34624 21622 34652 46922
rect 34704 22636 34756 22642
rect 34704 22578 34756 22584
rect 34716 22234 34744 22578
rect 34808 22234 34836 47126
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 38028 41414 38056 49200
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 38120 46578 38148 46990
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 39960 46866 39988 49200
rect 41248 47138 41276 49200
rect 40144 47110 41276 47138
rect 39960 46838 40080 46866
rect 38292 46504 38344 46510
rect 38292 46446 38344 46452
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 38304 46170 38332 46446
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38200 45960 38252 45966
rect 38200 45902 38252 45908
rect 38212 45830 38240 45902
rect 38200 45824 38252 45830
rect 38200 45766 38252 45772
rect 37292 41386 38056 41414
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 37292 24274 37320 41386
rect 37280 24268 37332 24274
rect 37280 24210 37332 24216
rect 37740 23724 37792 23730
rect 37740 23666 37792 23672
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 37752 23118 37780 23666
rect 36452 23112 36504 23118
rect 36452 23054 36504 23060
rect 37740 23112 37792 23118
rect 37740 23054 37792 23060
rect 36464 22642 36492 23054
rect 37752 22982 37780 23054
rect 37740 22976 37792 22982
rect 37740 22918 37792 22924
rect 37752 22778 37780 22918
rect 37740 22772 37792 22778
rect 37740 22714 37792 22720
rect 36452 22636 36504 22642
rect 36452 22578 36504 22584
rect 36636 22432 36688 22438
rect 36636 22374 36688 22380
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34704 22228 34756 22234
rect 34704 22170 34756 22176
rect 34796 22228 34848 22234
rect 34796 22170 34848 22176
rect 36648 22030 36676 22374
rect 37752 22030 37780 22714
rect 35348 22024 35400 22030
rect 35348 21966 35400 21972
rect 36360 22024 36412 22030
rect 36360 21966 36412 21972
rect 36636 22024 36688 22030
rect 36636 21966 36688 21972
rect 37740 22024 37792 22030
rect 37740 21966 37792 21972
rect 33416 21616 33468 21622
rect 33416 21558 33468 21564
rect 34612 21616 34664 21622
rect 34612 21558 34664 21564
rect 34796 21616 34848 21622
rect 34796 21558 34848 21564
rect 32864 21480 32916 21486
rect 32864 21422 32916 21428
rect 32680 21140 32732 21146
rect 32680 21082 32732 21088
rect 32588 19304 32640 19310
rect 32588 19246 32640 19252
rect 32600 18970 32628 19246
rect 32588 18964 32640 18970
rect 32588 18906 32640 18912
rect 32692 2514 32720 21082
rect 32876 20874 32904 21422
rect 33428 21146 33456 21558
rect 33416 21140 33468 21146
rect 33416 21082 33468 21088
rect 34808 20874 34836 21558
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35360 20874 35388 21966
rect 36372 21554 36400 21966
rect 37004 21956 37056 21962
rect 37004 21898 37056 21904
rect 36360 21548 36412 21554
rect 36360 21490 36412 21496
rect 35532 21480 35584 21486
rect 35532 21422 35584 21428
rect 36268 21480 36320 21486
rect 36268 21422 36320 21428
rect 35544 21078 35572 21422
rect 36280 21146 36308 21422
rect 37016 21350 37044 21898
rect 37752 21554 37780 21966
rect 38212 21622 38240 45766
rect 38752 45484 38804 45490
rect 38752 45426 38804 45432
rect 38660 44328 38712 44334
rect 38660 44270 38712 44276
rect 38672 43654 38700 44270
rect 38660 43648 38712 43654
rect 38660 43590 38712 43596
rect 38660 38752 38712 38758
rect 38660 38694 38712 38700
rect 38672 38350 38700 38694
rect 38660 38344 38712 38350
rect 38660 38286 38712 38292
rect 38672 37942 38700 38286
rect 38660 37936 38712 37942
rect 38660 37878 38712 37884
rect 38764 37874 38792 45426
rect 40052 44334 40080 46838
rect 38844 44328 38896 44334
rect 38844 44270 38896 44276
rect 40040 44328 40092 44334
rect 40040 44270 40092 44276
rect 38856 43994 38884 44270
rect 38844 43988 38896 43994
rect 38844 43930 38896 43936
rect 38936 43784 38988 43790
rect 38936 43726 38988 43732
rect 38948 38554 38976 43726
rect 39856 38888 39908 38894
rect 39856 38830 39908 38836
rect 38936 38548 38988 38554
rect 38936 38490 38988 38496
rect 38752 37868 38804 37874
rect 38752 37810 38804 37816
rect 38764 27878 38792 37810
rect 38752 27872 38804 27878
rect 38752 27814 38804 27820
rect 38764 24818 38792 27814
rect 38752 24812 38804 24818
rect 38752 24754 38804 24760
rect 38476 23656 38528 23662
rect 38476 23598 38528 23604
rect 38384 23180 38436 23186
rect 38384 23122 38436 23128
rect 38292 21888 38344 21894
rect 38292 21830 38344 21836
rect 38200 21616 38252 21622
rect 38200 21558 38252 21564
rect 37740 21548 37792 21554
rect 37740 21490 37792 21496
rect 38304 21486 38332 21830
rect 38292 21480 38344 21486
rect 38292 21422 38344 21428
rect 36636 21344 36688 21350
rect 36636 21286 36688 21292
rect 37004 21344 37056 21350
rect 37004 21286 37056 21292
rect 36268 21140 36320 21146
rect 36268 21082 36320 21088
rect 35532 21072 35584 21078
rect 35532 21014 35584 21020
rect 36280 20874 36308 21082
rect 32864 20868 32916 20874
rect 32864 20810 32916 20816
rect 34796 20868 34848 20874
rect 34796 20810 34848 20816
rect 35348 20868 35400 20874
rect 35348 20810 35400 20816
rect 36268 20868 36320 20874
rect 36268 20810 36320 20816
rect 32876 17678 32904 20810
rect 35254 20632 35310 20641
rect 35254 20567 35310 20576
rect 35268 20398 35296 20567
rect 34704 20392 34756 20398
rect 34704 20334 34756 20340
rect 35256 20392 35308 20398
rect 35256 20334 35308 20340
rect 33508 20256 33560 20262
rect 33508 20198 33560 20204
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 32956 19780 33008 19786
rect 32956 19722 33008 19728
rect 32968 18766 32996 19722
rect 33060 19378 33088 19790
rect 33520 19446 33548 20198
rect 34716 19990 34744 20334
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34704 19984 34756 19990
rect 34704 19926 34756 19932
rect 34716 19786 34744 19926
rect 34704 19780 34756 19786
rect 34704 19722 34756 19728
rect 33508 19440 33560 19446
rect 33508 19382 33560 19388
rect 33048 19372 33100 19378
rect 33048 19314 33100 19320
rect 33324 19372 33376 19378
rect 33324 19314 33376 19320
rect 33060 18902 33088 19314
rect 33048 18896 33100 18902
rect 33048 18838 33100 18844
rect 32956 18760 33008 18766
rect 32956 18702 33008 18708
rect 33336 18290 33364 19314
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 33600 18760 33652 18766
rect 33600 18702 33652 18708
rect 33324 18284 33376 18290
rect 33324 18226 33376 18232
rect 33612 18222 33640 18702
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 34796 18148 34848 18154
rect 34796 18090 34848 18096
rect 33048 18080 33100 18086
rect 33048 18022 33100 18028
rect 32864 17672 32916 17678
rect 32864 17614 32916 17620
rect 32876 14414 32904 17614
rect 33060 17202 33088 18022
rect 34808 17882 34836 18090
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34796 17876 34848 17882
rect 34796 17818 34848 17824
rect 33048 17196 33100 17202
rect 33048 17138 33100 17144
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 32864 14408 32916 14414
rect 32864 14350 32916 14356
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 32956 3596 33008 3602
rect 32956 3538 33008 3544
rect 32968 3058 32996 3538
rect 33140 3392 33192 3398
rect 33140 3334 33192 3340
rect 33152 3126 33180 3334
rect 33140 3120 33192 3126
rect 33140 3062 33192 3068
rect 32956 3052 33008 3058
rect 32956 2994 33008 3000
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 32680 2508 32732 2514
rect 32680 2450 32732 2456
rect 32496 2304 32548 2310
rect 32496 2246 32548 2252
rect 33520 800 33548 2926
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35360 2650 35388 20810
rect 36648 20602 36676 21286
rect 36820 20800 36872 20806
rect 36820 20742 36872 20748
rect 36636 20596 36688 20602
rect 36636 20538 36688 20544
rect 36544 20324 36596 20330
rect 36544 20266 36596 20272
rect 36556 20058 36584 20266
rect 36544 20052 36596 20058
rect 36544 19994 36596 20000
rect 35900 19916 35952 19922
rect 35900 19858 35952 19864
rect 35624 19168 35676 19174
rect 35624 19110 35676 19116
rect 35636 18358 35664 19110
rect 35624 18352 35676 18358
rect 35624 18294 35676 18300
rect 35912 18222 35940 19858
rect 36648 19446 36676 20538
rect 36832 20534 36860 20742
rect 36820 20528 36872 20534
rect 36820 20470 36872 20476
rect 36636 19440 36688 19446
rect 36636 19382 36688 19388
rect 36912 18692 36964 18698
rect 36912 18634 36964 18640
rect 35900 18216 35952 18222
rect 35900 18158 35952 18164
rect 36924 18086 36952 18634
rect 36912 18080 36964 18086
rect 36912 18022 36964 18028
rect 35440 17808 35492 17814
rect 35440 17750 35492 17756
rect 35452 17678 35480 17750
rect 35440 17672 35492 17678
rect 35440 17614 35492 17620
rect 36176 17672 36228 17678
rect 36176 17614 36228 17620
rect 36188 17134 36216 17614
rect 36176 17128 36228 17134
rect 36176 17070 36228 17076
rect 36544 4072 36596 4078
rect 36544 4014 36596 4020
rect 36556 3602 36584 4014
rect 37016 3670 37044 21286
rect 37372 19712 37424 19718
rect 37372 19654 37424 19660
rect 37096 19372 37148 19378
rect 37096 19314 37148 19320
rect 37108 18426 37136 19314
rect 37384 18766 37412 19654
rect 37372 18760 37424 18766
rect 37372 18702 37424 18708
rect 37384 18426 37412 18702
rect 37464 18624 37516 18630
rect 37464 18566 37516 18572
rect 37096 18420 37148 18426
rect 37096 18362 37148 18368
rect 37372 18420 37424 18426
rect 37372 18362 37424 18368
rect 37476 18358 37504 18566
rect 37464 18352 37516 18358
rect 37464 18294 37516 18300
rect 37556 18352 37608 18358
rect 37556 18294 37608 18300
rect 37188 18216 37240 18222
rect 37464 18216 37516 18222
rect 37240 18164 37464 18170
rect 37568 18170 37596 18294
rect 37516 18164 37596 18170
rect 37188 18158 37596 18164
rect 37096 18148 37148 18154
rect 37200 18142 37596 18158
rect 37096 18090 37148 18096
rect 37108 17746 37136 18090
rect 37464 18080 37516 18086
rect 37464 18022 37516 18028
rect 37476 17882 37504 18022
rect 37464 17876 37516 17882
rect 37464 17818 37516 17824
rect 37096 17740 37148 17746
rect 37096 17682 37148 17688
rect 37108 17202 37136 17682
rect 37096 17196 37148 17202
rect 37096 17138 37148 17144
rect 37280 5636 37332 5642
rect 37280 5578 37332 5584
rect 37292 4826 37320 5578
rect 37740 5296 37792 5302
rect 37740 5238 37792 5244
rect 37648 5160 37700 5166
rect 37648 5102 37700 5108
rect 37280 4820 37332 4826
rect 37280 4762 37332 4768
rect 37280 4616 37332 4622
rect 37280 4558 37332 4564
rect 37292 4282 37320 4558
rect 37280 4276 37332 4282
rect 37280 4218 37332 4224
rect 37660 4214 37688 5102
rect 37648 4208 37700 4214
rect 37648 4150 37700 4156
rect 37752 4146 37780 5238
rect 37740 4140 37792 4146
rect 37740 4082 37792 4088
rect 38200 4140 38252 4146
rect 38200 4082 38252 4088
rect 37372 3936 37424 3942
rect 37372 3878 37424 3884
rect 37004 3664 37056 3670
rect 37004 3606 37056 3612
rect 36544 3596 36596 3602
rect 36544 3538 36596 3544
rect 35348 2644 35400 2650
rect 35348 2586 35400 2592
rect 35900 2644 35952 2650
rect 35900 2586 35952 2592
rect 35912 2514 35940 2586
rect 35900 2508 35952 2514
rect 35900 2450 35952 2456
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35452 800 35480 2382
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 36096 800 36124 2314
rect 37384 1970 37412 3878
rect 38212 2446 38240 4082
rect 38304 3534 38332 21422
rect 38396 18222 38424 23122
rect 38384 18216 38436 18222
rect 38384 18158 38436 18164
rect 38292 3528 38344 3534
rect 38292 3470 38344 3476
rect 38304 2854 38332 3470
rect 38396 2922 38424 18158
rect 38488 5642 38516 23598
rect 38568 23520 38620 23526
rect 38568 23462 38620 23468
rect 38580 21894 38608 23462
rect 38568 21888 38620 21894
rect 38568 21830 38620 21836
rect 38580 20942 38608 21830
rect 38568 20936 38620 20942
rect 38568 20878 38620 20884
rect 38764 20262 38792 24754
rect 38948 23186 38976 38490
rect 39868 32026 39896 38830
rect 39948 37936 40000 37942
rect 39948 37878 40000 37884
rect 39856 32020 39908 32026
rect 39856 31962 39908 31968
rect 39212 24132 39264 24138
rect 39212 24074 39264 24080
rect 39224 23730 39252 24074
rect 39212 23724 39264 23730
rect 39212 23666 39264 23672
rect 39488 23316 39540 23322
rect 39488 23258 39540 23264
rect 38936 23180 38988 23186
rect 38936 23122 38988 23128
rect 39500 22778 39528 23258
rect 39488 22772 39540 22778
rect 39488 22714 39540 22720
rect 39500 22438 39528 22714
rect 39764 22636 39816 22642
rect 39764 22578 39816 22584
rect 39488 22432 39540 22438
rect 39488 22374 39540 22380
rect 39776 22030 39804 22578
rect 38844 22024 38896 22030
rect 38844 21966 38896 21972
rect 39764 22024 39816 22030
rect 39764 21966 39816 21972
rect 38856 20806 38884 21966
rect 39776 21457 39804 21966
rect 39762 21448 39818 21457
rect 39762 21383 39818 21392
rect 38844 20800 38896 20806
rect 38844 20742 38896 20748
rect 38752 20256 38804 20262
rect 38752 20198 38804 20204
rect 38856 11150 38884 20742
rect 39960 16250 39988 37878
rect 40040 23044 40092 23050
rect 40144 23032 40172 47110
rect 41512 47048 41564 47054
rect 41512 46990 41564 46996
rect 40408 46980 40460 46986
rect 40408 46922 40460 46928
rect 40224 45484 40276 45490
rect 40224 45426 40276 45432
rect 40236 37942 40264 45426
rect 40224 37936 40276 37942
rect 40224 37878 40276 37884
rect 40420 30802 40448 46922
rect 41524 46578 41552 46990
rect 41512 46572 41564 46578
rect 41512 46514 41564 46520
rect 41892 46442 41920 49200
rect 41880 46436 41932 46442
rect 41880 46378 41932 46384
rect 41052 46368 41104 46374
rect 41052 46310 41104 46316
rect 41064 46034 41092 46310
rect 42536 46034 42564 49200
rect 42708 47048 42760 47054
rect 42708 46990 42760 46996
rect 42616 46504 42668 46510
rect 42616 46446 42668 46452
rect 41052 46028 41104 46034
rect 41052 45970 41104 45976
rect 42524 46028 42576 46034
rect 42524 45970 42576 45976
rect 41236 45892 41288 45898
rect 41236 45834 41288 45840
rect 41248 45626 41276 45834
rect 42628 45626 42656 46446
rect 41236 45620 41288 45626
rect 41236 45562 41288 45568
rect 42616 45620 42668 45626
rect 42616 45562 42668 45568
rect 42720 45490 42748 46990
rect 42708 45484 42760 45490
rect 42708 45426 42760 45432
rect 43180 45422 43208 49200
rect 43824 47054 43852 49200
rect 44468 47122 44496 49200
rect 45112 47410 45140 49200
rect 45112 47382 45508 47410
rect 44456 47116 44508 47122
rect 44456 47058 44508 47064
rect 43812 47048 43864 47054
rect 43812 46990 43864 46996
rect 45100 47048 45152 47054
rect 45100 46990 45152 46996
rect 43352 46980 43404 46986
rect 43352 46922 43404 46928
rect 43168 45416 43220 45422
rect 43168 45358 43220 45364
rect 43260 45348 43312 45354
rect 43260 45290 43312 45296
rect 43272 45082 43300 45290
rect 43260 45076 43312 45082
rect 43260 45018 43312 45024
rect 43168 44872 43220 44878
rect 43168 44814 43220 44820
rect 41144 38820 41196 38826
rect 41144 38762 41196 38768
rect 40684 38412 40736 38418
rect 40684 38354 40736 38360
rect 40696 36310 40724 38354
rect 40684 36304 40736 36310
rect 40684 36246 40736 36252
rect 40408 30796 40460 30802
rect 40408 30738 40460 30744
rect 40592 24744 40644 24750
rect 40592 24686 40644 24692
rect 40960 24744 41012 24750
rect 40960 24686 41012 24692
rect 40604 23866 40632 24686
rect 40972 24614 41000 24686
rect 40960 24608 41012 24614
rect 40960 24550 41012 24556
rect 40592 23860 40644 23866
rect 40592 23802 40644 23808
rect 40604 23186 40632 23802
rect 41156 23730 41184 38762
rect 43180 38418 43208 44814
rect 43168 38412 43220 38418
rect 43168 38354 43220 38360
rect 41420 33312 41472 33318
rect 41420 33254 41472 33260
rect 41432 32502 41460 33254
rect 41420 32496 41472 32502
rect 41420 32438 41472 32444
rect 43364 29238 43392 46922
rect 43444 45824 43496 45830
rect 43444 45766 43496 45772
rect 43456 45558 43484 45766
rect 43444 45552 43496 45558
rect 43444 45494 43496 45500
rect 44824 45552 44876 45558
rect 44824 45494 44876 45500
rect 43352 29232 43404 29238
rect 43352 29174 43404 29180
rect 42432 27668 42484 27674
rect 42432 27610 42484 27616
rect 41236 24064 41288 24070
rect 41236 24006 41288 24012
rect 41248 23730 41276 24006
rect 41144 23724 41196 23730
rect 41144 23666 41196 23672
rect 41236 23724 41288 23730
rect 41236 23666 41288 23672
rect 41156 23254 41184 23666
rect 41144 23248 41196 23254
rect 41144 23190 41196 23196
rect 40592 23180 40644 23186
rect 40592 23122 40644 23128
rect 40092 23004 40172 23032
rect 40776 23044 40828 23050
rect 40040 22986 40092 22992
rect 40776 22986 40828 22992
rect 41788 23044 41840 23050
rect 41788 22986 41840 22992
rect 40788 22778 40816 22986
rect 40776 22772 40828 22778
rect 40776 22714 40828 22720
rect 40040 22432 40092 22438
rect 40040 22374 40092 22380
rect 40052 22030 40080 22374
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 40316 21956 40368 21962
rect 40316 21898 40368 21904
rect 39948 16244 40000 16250
rect 39948 16186 40000 16192
rect 38844 11144 38896 11150
rect 38844 11086 38896 11092
rect 38476 5636 38528 5642
rect 38476 5578 38528 5584
rect 38488 5166 38516 5578
rect 38476 5160 38528 5166
rect 38476 5102 38528 5108
rect 39120 5024 39172 5030
rect 39120 4966 39172 4972
rect 39948 5024 40000 5030
rect 39948 4966 40000 4972
rect 39132 4622 39160 4966
rect 39960 4690 39988 4966
rect 39948 4684 40000 4690
rect 39948 4626 40000 4632
rect 39120 4616 39172 4622
rect 39120 4558 39172 4564
rect 40132 4548 40184 4554
rect 40132 4490 40184 4496
rect 39304 4140 39356 4146
rect 39304 4082 39356 4088
rect 40040 4140 40092 4146
rect 40040 4082 40092 4088
rect 39316 2990 39344 4082
rect 39856 3460 39908 3466
rect 39856 3402 39908 3408
rect 39868 3194 39896 3402
rect 39856 3188 39908 3194
rect 39856 3130 39908 3136
rect 39948 3052 40000 3058
rect 39948 2994 40000 3000
rect 39304 2984 39356 2990
rect 39304 2926 39356 2932
rect 38384 2916 38436 2922
rect 38384 2858 38436 2864
rect 38292 2848 38344 2854
rect 38292 2790 38344 2796
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 38200 2440 38252 2446
rect 38200 2382 38252 2388
rect 37372 1964 37424 1970
rect 37372 1906 37424 1912
rect 38028 800 38056 2382
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 39316 800 39344 2314
rect 39960 800 39988 2994
rect 40052 2922 40080 4082
rect 40144 3670 40172 4490
rect 40328 4214 40356 21898
rect 41694 21584 41750 21593
rect 41694 21519 41696 21528
rect 41748 21519 41750 21528
rect 41696 21490 41748 21496
rect 41800 18358 41828 22986
rect 42444 22030 42472 27610
rect 42984 24200 43036 24206
rect 42984 24142 43036 24148
rect 42800 24132 42852 24138
rect 42800 24074 42852 24080
rect 42524 23656 42576 23662
rect 42524 23598 42576 23604
rect 42536 23050 42564 23598
rect 42812 23118 42840 24074
rect 42996 23526 43024 24142
rect 43168 24064 43220 24070
rect 43168 24006 43220 24012
rect 42984 23520 43036 23526
rect 42984 23462 43036 23468
rect 42800 23112 42852 23118
rect 42800 23054 42852 23060
rect 42524 23044 42576 23050
rect 42524 22986 42576 22992
rect 42536 22778 42564 22986
rect 42524 22772 42576 22778
rect 42524 22714 42576 22720
rect 42812 22574 42840 23054
rect 42996 22642 43024 23462
rect 43180 23322 43208 24006
rect 44836 23730 44864 45494
rect 45008 45416 45060 45422
rect 45008 45358 45060 45364
rect 45020 45082 45048 45358
rect 45008 45076 45060 45082
rect 45008 45018 45060 45024
rect 45112 44402 45140 46990
rect 45376 46980 45428 46986
rect 45376 46922 45428 46928
rect 45192 46504 45244 46510
rect 45192 46446 45244 46452
rect 45204 45082 45232 46446
rect 45192 45076 45244 45082
rect 45192 45018 45244 45024
rect 45388 44538 45416 46922
rect 45480 46866 45508 47382
rect 45480 46838 45600 46866
rect 45468 45824 45520 45830
rect 45468 45766 45520 45772
rect 45480 45234 45508 45766
rect 45572 45422 45600 46838
rect 45652 46504 45704 46510
rect 45652 46446 45704 46452
rect 45560 45416 45612 45422
rect 45560 45358 45612 45364
rect 45480 45206 45600 45234
rect 45572 44878 45600 45206
rect 45664 45082 45692 46446
rect 45756 45966 45784 49200
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 45836 45960 45888 45966
rect 45836 45902 45888 45908
rect 45652 45076 45704 45082
rect 45652 45018 45704 45024
rect 45560 44872 45612 44878
rect 45560 44814 45612 44820
rect 45376 44532 45428 44538
rect 45376 44474 45428 44480
rect 45848 44402 45876 45902
rect 46020 45824 46072 45830
rect 46020 45766 46072 45772
rect 45100 44396 45152 44402
rect 45100 44338 45152 44344
rect 45836 44396 45888 44402
rect 45836 44338 45888 44344
rect 46032 39302 46060 45766
rect 46400 45626 46428 49200
rect 46846 47696 46902 47705
rect 46846 47631 46902 47640
rect 46478 47016 46534 47025
rect 46478 46951 46534 46960
rect 46388 45620 46440 45626
rect 46388 45562 46440 45568
rect 46204 44396 46256 44402
rect 46204 44338 46256 44344
rect 46020 39296 46072 39302
rect 46020 39238 46072 39244
rect 46216 38894 46244 44338
rect 46492 44146 46520 46951
rect 46860 46510 46888 47631
rect 46848 46504 46900 46510
rect 46848 46446 46900 46452
rect 46848 46164 46900 46170
rect 46848 46106 46900 46112
rect 46756 45280 46808 45286
rect 46756 45222 46808 45228
rect 46400 44118 46520 44146
rect 46204 38888 46256 38894
rect 46204 38830 46256 38836
rect 46216 32434 46244 38830
rect 46296 38344 46348 38350
rect 46296 38286 46348 38292
rect 46308 37942 46336 38286
rect 46296 37936 46348 37942
rect 46296 37878 46348 37884
rect 46296 32904 46348 32910
rect 46296 32846 46348 32852
rect 46204 32428 46256 32434
rect 46204 32370 46256 32376
rect 46308 32026 46336 32846
rect 46296 32020 46348 32026
rect 46296 31962 46348 31968
rect 46400 31754 46428 44118
rect 46572 42220 46624 42226
rect 46572 42162 46624 42168
rect 46480 42016 46532 42022
rect 46480 41958 46532 41964
rect 46492 41682 46520 41958
rect 46480 41676 46532 41682
rect 46480 41618 46532 41624
rect 46480 39840 46532 39846
rect 46480 39782 46532 39788
rect 46492 39506 46520 39782
rect 46480 39500 46532 39506
rect 46480 39442 46532 39448
rect 46584 35894 46612 42162
rect 46768 40050 46796 45222
rect 46860 42226 46888 46106
rect 47044 46034 47072 49200
rect 47400 47184 47452 47190
rect 47400 47126 47452 47132
rect 47032 46028 47084 46034
rect 47032 45970 47084 45976
rect 47032 44940 47084 44946
rect 47032 44882 47084 44888
rect 46940 44192 46992 44198
rect 46940 44134 46992 44140
rect 46952 43858 46980 44134
rect 46940 43852 46992 43858
rect 46940 43794 46992 43800
rect 47044 43314 47072 44882
rect 47032 43308 47084 43314
rect 47032 43250 47084 43256
rect 46940 42628 46992 42634
rect 46940 42570 46992 42576
rect 46952 42362 46980 42570
rect 46940 42356 46992 42362
rect 46940 42298 46992 42304
rect 46848 42220 46900 42226
rect 46848 42162 46900 42168
rect 46756 40044 46808 40050
rect 46756 39986 46808 39992
rect 46662 39536 46718 39545
rect 46662 39471 46718 39480
rect 46216 31726 46428 31754
rect 46492 35866 46612 35894
rect 46020 30660 46072 30666
rect 46020 30602 46072 30608
rect 45650 30016 45706 30025
rect 45650 29951 45706 29960
rect 45558 28656 45614 28665
rect 45558 28591 45614 28600
rect 45572 27674 45600 28591
rect 45560 27668 45612 27674
rect 45560 27610 45612 27616
rect 45192 26376 45244 26382
rect 45192 26318 45244 26324
rect 45204 24818 45232 26318
rect 45192 24812 45244 24818
rect 45192 24754 45244 24760
rect 45376 24744 45428 24750
rect 45376 24686 45428 24692
rect 45388 23866 45416 24686
rect 45560 24676 45612 24682
rect 45560 24618 45612 24624
rect 45572 23905 45600 24618
rect 45664 24342 45692 29951
rect 45742 26616 45798 26625
rect 45742 26551 45798 26560
rect 45652 24336 45704 24342
rect 45652 24278 45704 24284
rect 45558 23896 45614 23905
rect 45376 23860 45428 23866
rect 45558 23831 45614 23840
rect 45376 23802 45428 23808
rect 43352 23724 43404 23730
rect 43352 23666 43404 23672
rect 44824 23724 44876 23730
rect 44824 23666 44876 23672
rect 43168 23316 43220 23322
rect 43168 23258 43220 23264
rect 43364 23186 43392 23666
rect 43628 23316 43680 23322
rect 43628 23258 43680 23264
rect 43352 23180 43404 23186
rect 43352 23122 43404 23128
rect 43168 22976 43220 22982
rect 43168 22918 43220 22924
rect 43180 22642 43208 22918
rect 42984 22636 43036 22642
rect 42984 22578 43036 22584
rect 43168 22636 43220 22642
rect 43168 22578 43220 22584
rect 42800 22568 42852 22574
rect 42800 22510 42852 22516
rect 42432 22024 42484 22030
rect 42432 21966 42484 21972
rect 42708 21956 42760 21962
rect 42708 21898 42760 21904
rect 41880 21548 41932 21554
rect 41880 21490 41932 21496
rect 41892 21418 41920 21490
rect 42720 21486 42748 21898
rect 42812 21690 42840 22510
rect 43076 22160 43128 22166
rect 43076 22102 43128 22108
rect 42800 21684 42852 21690
rect 42800 21626 42852 21632
rect 42892 21684 42944 21690
rect 42892 21626 42944 21632
rect 42708 21480 42760 21486
rect 42708 21422 42760 21428
rect 41880 21412 41932 21418
rect 41880 21354 41932 21360
rect 41788 18352 41840 18358
rect 41788 18294 41840 18300
rect 41800 18154 41828 18294
rect 41788 18148 41840 18154
rect 41788 18090 41840 18096
rect 40408 5228 40460 5234
rect 40408 5170 40460 5176
rect 40420 4826 40448 5170
rect 41236 5160 41288 5166
rect 41236 5102 41288 5108
rect 40408 4820 40460 4826
rect 40408 4762 40460 4768
rect 40316 4208 40368 4214
rect 40316 4150 40368 4156
rect 40224 3936 40276 3942
rect 40224 3878 40276 3884
rect 40132 3664 40184 3670
rect 40132 3606 40184 3612
rect 40236 3534 40264 3878
rect 40224 3528 40276 3534
rect 40224 3470 40276 3476
rect 40040 2916 40092 2922
rect 40040 2858 40092 2864
rect 40052 2446 40080 2858
rect 40328 2650 40356 4150
rect 41248 4146 41276 5102
rect 41512 4752 41564 4758
rect 41512 4694 41564 4700
rect 41236 4140 41288 4146
rect 41236 4082 41288 4088
rect 41420 3936 41472 3942
rect 41420 3878 41472 3884
rect 41052 3528 41104 3534
rect 41052 3470 41104 3476
rect 41064 3194 41092 3470
rect 41328 3460 41380 3466
rect 41328 3402 41380 3408
rect 41052 3188 41104 3194
rect 41052 3130 41104 3136
rect 40592 3052 40644 3058
rect 40592 2994 40644 3000
rect 41236 3052 41288 3058
rect 41236 2994 41288 3000
rect 40604 2650 40632 2994
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40316 2644 40368 2650
rect 40316 2586 40368 2592
rect 40592 2644 40644 2650
rect 40592 2586 40644 2592
rect 40696 2514 40724 2926
rect 40684 2508 40736 2514
rect 40684 2450 40736 2456
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 40592 2440 40644 2446
rect 40592 2382 40644 2388
rect 40604 800 40632 2382
rect 41248 800 41276 2994
rect 41340 2854 41368 3402
rect 41328 2848 41380 2854
rect 41328 2790 41380 2796
rect 41432 1902 41460 3878
rect 41524 2922 41552 4694
rect 41800 4690 41828 18090
rect 41788 4684 41840 4690
rect 41788 4626 41840 4632
rect 41800 3602 41828 4626
rect 41788 3596 41840 3602
rect 41788 3538 41840 3544
rect 41512 2916 41564 2922
rect 41512 2858 41564 2864
rect 41892 2582 41920 21354
rect 42904 21350 42932 21626
rect 43088 21554 43116 22102
rect 43168 21888 43220 21894
rect 43168 21830 43220 21836
rect 43076 21548 43128 21554
rect 43076 21490 43128 21496
rect 43180 21434 43208 21830
rect 42996 21406 43208 21434
rect 42892 21344 42944 21350
rect 42892 21286 42944 21292
rect 42708 21140 42760 21146
rect 42708 21082 42760 21088
rect 42720 20466 42748 21082
rect 42892 21072 42944 21078
rect 42892 21014 42944 21020
rect 42904 20806 42932 21014
rect 42996 20942 43024 21406
rect 43076 21344 43128 21350
rect 43076 21286 43128 21292
rect 43088 20942 43116 21286
rect 42984 20936 43036 20942
rect 42984 20878 43036 20884
rect 43076 20936 43128 20942
rect 43076 20878 43128 20884
rect 42892 20800 42944 20806
rect 42892 20742 42944 20748
rect 42708 20460 42760 20466
rect 42708 20402 42760 20408
rect 43260 20460 43312 20466
rect 43260 20402 43312 20408
rect 42720 19786 42748 20402
rect 43272 19854 43300 20402
rect 43260 19848 43312 19854
rect 43260 19790 43312 19796
rect 42708 19780 42760 19786
rect 42708 19722 42760 19728
rect 42720 19378 42748 19722
rect 42708 19372 42760 19378
rect 42708 19314 42760 19320
rect 42800 18692 42852 18698
rect 42800 18634 42852 18640
rect 42812 18426 42840 18634
rect 42800 18420 42852 18426
rect 42800 18362 42852 18368
rect 43364 6914 43392 23122
rect 43640 21593 43668 23258
rect 44836 23118 44864 23666
rect 45192 23656 45244 23662
rect 45192 23598 45244 23604
rect 45652 23656 45704 23662
rect 45652 23598 45704 23604
rect 45204 23254 45232 23598
rect 45192 23248 45244 23254
rect 45192 23190 45244 23196
rect 44824 23112 44876 23118
rect 44824 23054 44876 23060
rect 44272 23044 44324 23050
rect 44272 22986 44324 22992
rect 44284 22778 44312 22986
rect 45100 22976 45152 22982
rect 45100 22918 45152 22924
rect 44272 22772 44324 22778
rect 44272 22714 44324 22720
rect 45112 22642 45140 22918
rect 45664 22778 45692 23598
rect 45652 22772 45704 22778
rect 45652 22714 45704 22720
rect 45756 22710 45784 26551
rect 45836 25288 45888 25294
rect 45836 25230 45888 25236
rect 45744 22704 45796 22710
rect 45744 22646 45796 22652
rect 45100 22636 45152 22642
rect 45100 22578 45152 22584
rect 45560 22636 45612 22642
rect 45560 22578 45612 22584
rect 45192 22228 45244 22234
rect 45192 22170 45244 22176
rect 45204 22030 45232 22170
rect 45192 22024 45244 22030
rect 45192 21966 45244 21972
rect 45376 22024 45428 22030
rect 45376 21966 45428 21972
rect 45388 21622 45416 21966
rect 45572 21962 45600 22578
rect 45848 22030 45876 25230
rect 45928 24200 45980 24206
rect 45928 24142 45980 24148
rect 45940 23225 45968 24142
rect 45926 23216 45982 23225
rect 45926 23151 45982 23160
rect 45928 22432 45980 22438
rect 45928 22374 45980 22380
rect 45940 22166 45968 22374
rect 45928 22160 45980 22166
rect 45928 22102 45980 22108
rect 45836 22024 45888 22030
rect 45836 21966 45888 21972
rect 45560 21956 45612 21962
rect 45744 21956 45796 21962
rect 45612 21916 45692 21944
rect 45560 21898 45612 21904
rect 45376 21616 45428 21622
rect 43626 21584 43682 21593
rect 45376 21558 45428 21564
rect 43626 21519 43628 21528
rect 43680 21519 43682 21528
rect 43812 21548 43864 21554
rect 43628 21490 43680 21496
rect 43812 21490 43864 21496
rect 44272 21548 44324 21554
rect 44272 21490 44324 21496
rect 43640 21459 43668 21490
rect 43824 21418 43852 21490
rect 43812 21412 43864 21418
rect 43812 21354 43864 21360
rect 43628 21140 43680 21146
rect 43628 21082 43680 21088
rect 43640 20806 43668 21082
rect 43720 20936 43772 20942
rect 43720 20878 43772 20884
rect 43628 20800 43680 20806
rect 43628 20742 43680 20748
rect 43732 20534 43760 20878
rect 43812 20800 43864 20806
rect 43812 20742 43864 20748
rect 43720 20528 43772 20534
rect 43720 20470 43772 20476
rect 43824 20398 43852 20742
rect 44284 20466 44312 21490
rect 45008 21480 45060 21486
rect 45008 21422 45060 21428
rect 43904 20460 43956 20466
rect 43904 20402 43956 20408
rect 44272 20460 44324 20466
rect 44272 20402 44324 20408
rect 43812 20392 43864 20398
rect 43812 20334 43864 20340
rect 43824 18834 43852 20334
rect 43916 19990 43944 20402
rect 43904 19984 43956 19990
rect 43904 19926 43956 19932
rect 43916 19514 43944 19926
rect 43996 19848 44048 19854
rect 43996 19790 44048 19796
rect 43904 19508 43956 19514
rect 43904 19450 43956 19456
rect 44008 19378 44036 19790
rect 43996 19372 44048 19378
rect 43996 19314 44048 19320
rect 43812 18828 43864 18834
rect 43812 18770 43864 18776
rect 43904 18216 43956 18222
rect 43904 18158 43956 18164
rect 43916 17746 43944 18158
rect 44284 17882 44312 20402
rect 45020 20058 45048 21422
rect 45560 20392 45612 20398
rect 45560 20334 45612 20340
rect 45008 20052 45060 20058
rect 45008 19994 45060 20000
rect 45468 19168 45520 19174
rect 45468 19110 45520 19116
rect 45480 18834 45508 19110
rect 45468 18828 45520 18834
rect 45468 18770 45520 18776
rect 45100 18760 45152 18766
rect 45100 18702 45152 18708
rect 45376 18760 45428 18766
rect 45376 18702 45428 18708
rect 44456 18692 44508 18698
rect 44456 18634 44508 18640
rect 44364 18624 44416 18630
rect 44364 18566 44416 18572
rect 44376 18290 44404 18566
rect 44364 18284 44416 18290
rect 44364 18226 44416 18232
rect 44272 17876 44324 17882
rect 44272 17818 44324 17824
rect 44180 17808 44232 17814
rect 44180 17750 44232 17756
rect 43904 17740 43956 17746
rect 43904 17682 43956 17688
rect 43904 17128 43956 17134
rect 43904 17070 43956 17076
rect 43916 16794 43944 17070
rect 43904 16788 43956 16794
rect 43904 16730 43956 16736
rect 44192 13938 44220 17750
rect 44180 13932 44232 13938
rect 44180 13874 44232 13880
rect 43180 6886 43392 6914
rect 43180 5778 43208 6886
rect 43168 5772 43220 5778
rect 43168 5714 43220 5720
rect 42248 5636 42300 5642
rect 42248 5578 42300 5584
rect 42260 5370 42288 5578
rect 42248 5364 42300 5370
rect 42248 5306 42300 5312
rect 42892 5228 42944 5234
rect 42892 5170 42944 5176
rect 42524 4480 42576 4486
rect 42524 4422 42576 4428
rect 42536 4146 42564 4422
rect 42524 4140 42576 4146
rect 42524 4082 42576 4088
rect 42432 3596 42484 3602
rect 42432 3538 42484 3544
rect 42340 3392 42392 3398
rect 42340 3334 42392 3340
rect 41880 2576 41932 2582
rect 41880 2518 41932 2524
rect 41420 1896 41472 1902
rect 41420 1838 41472 1844
rect 42352 1714 42380 3334
rect 42444 3058 42472 3538
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 42536 2514 42564 4082
rect 42904 4078 42932 5170
rect 43180 4690 43208 5714
rect 43168 4684 43220 4690
rect 43168 4626 43220 4632
rect 42892 4072 42944 4078
rect 42892 4014 42944 4020
rect 44468 3738 44496 18634
rect 45112 18426 45140 18702
rect 45100 18420 45152 18426
rect 45100 18362 45152 18368
rect 44732 18216 44784 18222
rect 44732 18158 44784 18164
rect 44744 16114 44772 18158
rect 45112 17678 45140 18362
rect 45388 17678 45416 18702
rect 45572 18154 45600 20334
rect 45560 18148 45612 18154
rect 45560 18090 45612 18096
rect 45100 17672 45152 17678
rect 45100 17614 45152 17620
rect 45376 17672 45428 17678
rect 45376 17614 45428 17620
rect 45388 17338 45416 17614
rect 45376 17332 45428 17338
rect 45376 17274 45428 17280
rect 45376 17128 45428 17134
rect 45376 17070 45428 17076
rect 44732 16108 44784 16114
rect 44732 16050 44784 16056
rect 45100 16040 45152 16046
rect 45100 15982 45152 15988
rect 45112 15706 45140 15982
rect 45100 15700 45152 15706
rect 45100 15642 45152 15648
rect 45008 14408 45060 14414
rect 45008 14350 45060 14356
rect 45020 13870 45048 14350
rect 45192 14340 45244 14346
rect 45192 14282 45244 14288
rect 45204 14074 45232 14282
rect 45192 14068 45244 14074
rect 45192 14010 45244 14016
rect 45008 13864 45060 13870
rect 45008 13806 45060 13812
rect 45388 6914 45416 17070
rect 45664 16658 45692 21916
rect 45744 21898 45796 21904
rect 45756 21554 45784 21898
rect 45848 21690 45876 21966
rect 45836 21684 45888 21690
rect 45836 21626 45888 21632
rect 45744 21548 45796 21554
rect 45744 21490 45796 21496
rect 46032 21434 46060 30602
rect 46216 25786 46244 31726
rect 46492 31482 46520 35866
rect 46480 31476 46532 31482
rect 46480 31418 46532 31424
rect 46478 31376 46534 31385
rect 46478 31311 46534 31320
rect 46296 28076 46348 28082
rect 46296 28018 46348 28024
rect 46308 25906 46336 28018
rect 46296 25900 46348 25906
rect 46296 25842 46348 25848
rect 46492 25786 46520 31311
rect 46572 26920 46624 26926
rect 46572 26862 46624 26868
rect 46216 25758 46336 25786
rect 46204 22568 46256 22574
rect 46202 22536 46204 22545
rect 46256 22536 46258 22545
rect 46202 22471 46258 22480
rect 45940 21406 46060 21434
rect 45940 21078 45968 21406
rect 46020 21344 46072 21350
rect 46020 21286 46072 21292
rect 45928 21072 45980 21078
rect 45928 21014 45980 21020
rect 46032 20534 46060 21286
rect 46020 20528 46072 20534
rect 46020 20470 46072 20476
rect 45836 19848 45888 19854
rect 45836 19790 45888 19796
rect 46112 19848 46164 19854
rect 46112 19790 46164 19796
rect 45744 19780 45796 19786
rect 45744 19722 45796 19728
rect 45756 19242 45784 19722
rect 45744 19236 45796 19242
rect 45744 19178 45796 19184
rect 45756 18698 45784 19178
rect 45744 18692 45796 18698
rect 45744 18634 45796 18640
rect 45652 16652 45704 16658
rect 45652 16594 45704 16600
rect 45558 15736 45614 15745
rect 45558 15671 45614 15680
rect 45572 15638 45600 15671
rect 45560 15632 45612 15638
rect 45560 15574 45612 15580
rect 45664 15502 45692 16594
rect 45652 15496 45704 15502
rect 45652 15438 45704 15444
rect 45664 15026 45692 15438
rect 45652 15020 45704 15026
rect 45652 14962 45704 14968
rect 45756 12434 45784 18634
rect 45848 18465 45876 19790
rect 45928 19712 45980 19718
rect 45928 19654 45980 19660
rect 45940 19378 45968 19654
rect 46020 19508 46072 19514
rect 46020 19450 46072 19456
rect 45928 19372 45980 19378
rect 45928 19314 45980 19320
rect 45834 18456 45890 18465
rect 45834 18391 45890 18400
rect 45756 12406 45968 12434
rect 45468 7812 45520 7818
rect 45468 7754 45520 7760
rect 45560 7812 45612 7818
rect 45560 7754 45612 7760
rect 45112 6886 45416 6914
rect 44456 3732 44508 3738
rect 44456 3674 44508 3680
rect 42616 3392 42668 3398
rect 42616 3334 42668 3340
rect 42628 3126 42656 3334
rect 42616 3120 42668 3126
rect 42616 3062 42668 3068
rect 43168 2984 43220 2990
rect 43168 2926 43220 2932
rect 42524 2508 42576 2514
rect 42524 2450 42576 2456
rect 42352 1686 42564 1714
rect 42536 800 42564 1686
rect 43180 800 43208 2926
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 45112 800 45140 6886
rect 45480 4758 45508 7754
rect 45572 7410 45600 7754
rect 45560 7404 45612 7410
rect 45560 7346 45612 7352
rect 45940 5370 45968 12406
rect 46032 11082 46060 19450
rect 46124 19378 46152 19790
rect 46112 19372 46164 19378
rect 46112 19314 46164 19320
rect 46124 18902 46152 19314
rect 46204 19168 46256 19174
rect 46204 19110 46256 19116
rect 46112 18896 46164 18902
rect 46112 18838 46164 18844
rect 46216 18358 46244 19110
rect 46204 18352 46256 18358
rect 46204 18294 46256 18300
rect 46308 17610 46336 25758
rect 46400 25758 46520 25786
rect 46400 20505 46428 25758
rect 46480 25696 46532 25702
rect 46480 25638 46532 25644
rect 46492 25362 46520 25638
rect 46480 25356 46532 25362
rect 46480 25298 46532 25304
rect 46480 24608 46532 24614
rect 46480 24550 46532 24556
rect 46492 24274 46520 24550
rect 46480 24268 46532 24274
rect 46480 24210 46532 24216
rect 46480 22568 46532 22574
rect 46480 22510 46532 22516
rect 46492 21146 46520 22510
rect 46584 21962 46612 26862
rect 46676 23662 46704 39471
rect 46768 38706 46796 39986
rect 46768 38678 46888 38706
rect 46756 38548 46808 38554
rect 46756 38490 46808 38496
rect 46768 37874 46796 38490
rect 46860 38434 46888 38678
rect 46860 38406 46980 38434
rect 46848 38276 46900 38282
rect 46848 38218 46900 38224
rect 46860 38010 46888 38218
rect 46848 38004 46900 38010
rect 46848 37946 46900 37952
rect 46952 37890 46980 38406
rect 47308 38208 47360 38214
rect 47308 38150 47360 38156
rect 46756 37868 46808 37874
rect 46756 37810 46808 37816
rect 46860 37862 46980 37890
rect 46860 35894 46888 37862
rect 46768 35866 46888 35894
rect 46768 26926 46796 35866
rect 47124 35488 47176 35494
rect 47124 35430 47176 35436
rect 47136 34066 47164 35430
rect 47216 34400 47268 34406
rect 47216 34342 47268 34348
rect 47124 34060 47176 34066
rect 47124 34002 47176 34008
rect 47228 33930 47256 34342
rect 47216 33924 47268 33930
rect 47216 33866 47268 33872
rect 46848 33516 46900 33522
rect 46848 33458 46900 33464
rect 46860 33425 46888 33458
rect 46846 33416 46902 33425
rect 46846 33351 46902 33360
rect 47032 32972 47084 32978
rect 47032 32914 47084 32920
rect 46940 32836 46992 32842
rect 46940 32778 46992 32784
rect 46952 32570 46980 32778
rect 47044 32570 47072 32914
rect 46940 32564 46992 32570
rect 46940 32506 46992 32512
rect 47032 32564 47084 32570
rect 47032 32506 47084 32512
rect 46848 31476 46900 31482
rect 46848 31418 46900 31424
rect 46756 26920 46808 26926
rect 46756 26862 46808 26868
rect 46860 25378 46888 31418
rect 47032 30796 47084 30802
rect 47032 30738 47084 30744
rect 46940 27872 46992 27878
rect 46940 27814 46992 27820
rect 46952 27538 46980 27814
rect 46940 27532 46992 27538
rect 46940 27474 46992 27480
rect 46768 25350 46888 25378
rect 46768 24818 46796 25350
rect 46846 25256 46902 25265
rect 46846 25191 46902 25200
rect 46756 24812 46808 24818
rect 46756 24754 46808 24760
rect 46860 24750 46888 25191
rect 46848 24744 46900 24750
rect 46848 24686 46900 24692
rect 46664 23656 46716 23662
rect 46664 23598 46716 23604
rect 47044 23322 47072 30738
rect 47032 23316 47084 23322
rect 47032 23258 47084 23264
rect 47216 23044 47268 23050
rect 47216 22986 47268 22992
rect 46664 22432 46716 22438
rect 46664 22374 46716 22380
rect 46572 21956 46624 21962
rect 46572 21898 46624 21904
rect 46676 21894 46704 22374
rect 47228 21962 47256 22986
rect 47216 21956 47268 21962
rect 47216 21898 47268 21904
rect 46664 21888 46716 21894
rect 46664 21830 46716 21836
rect 46676 21622 46704 21830
rect 46664 21616 46716 21622
rect 46664 21558 46716 21564
rect 46480 21140 46532 21146
rect 46480 21082 46532 21088
rect 46386 20496 46442 20505
rect 47228 20466 47256 21898
rect 46386 20431 46442 20440
rect 47216 20460 47268 20466
rect 47216 20402 47268 20408
rect 47320 20346 47348 38150
rect 47412 32366 47440 47126
rect 47688 47054 47716 49200
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47952 46572 48004 46578
rect 47952 46514 48004 46520
rect 47964 46345 47992 46514
rect 48044 46368 48096 46374
rect 47950 46336 48006 46345
rect 48044 46310 48096 46316
rect 47950 46271 48006 46280
rect 47584 46096 47636 46102
rect 47584 46038 47636 46044
rect 47596 42226 47624 46038
rect 47676 44804 47728 44810
rect 47676 44746 47728 44752
rect 47688 44538 47716 44746
rect 47676 44532 47728 44538
rect 47676 44474 47728 44480
rect 47768 43104 47820 43110
rect 47768 43046 47820 43052
rect 47780 42770 47808 43046
rect 47768 42764 47820 42770
rect 47768 42706 47820 42712
rect 47584 42220 47636 42226
rect 47584 42162 47636 42168
rect 47492 40928 47544 40934
rect 47492 40870 47544 40876
rect 47400 32360 47452 32366
rect 47400 32302 47452 32308
rect 47504 24410 47532 40870
rect 47596 38214 47624 42162
rect 47676 41540 47728 41546
rect 47676 41482 47728 41488
rect 47688 40730 47716 41482
rect 47952 41132 48004 41138
rect 47952 41074 48004 41080
rect 47964 40905 47992 41074
rect 47950 40896 48006 40905
rect 47950 40831 48006 40840
rect 47676 40724 47728 40730
rect 47676 40666 47728 40672
rect 47768 39840 47820 39846
rect 47768 39782 47820 39788
rect 47780 39574 47808 39782
rect 47768 39568 47820 39574
rect 47768 39510 47820 39516
rect 47860 38956 47912 38962
rect 47860 38898 47912 38904
rect 47872 38865 47900 38898
rect 47858 38856 47914 38865
rect 47858 38791 47914 38800
rect 47584 38208 47636 38214
rect 47584 38150 47636 38156
rect 47860 34944 47912 34950
rect 47860 34886 47912 34892
rect 47768 34604 47820 34610
rect 47768 34546 47820 34552
rect 47676 34060 47728 34066
rect 47676 34002 47728 34008
rect 47688 30802 47716 34002
rect 47780 33658 47808 34546
rect 47768 33652 47820 33658
rect 47768 33594 47820 33600
rect 47768 33516 47820 33522
rect 47768 33458 47820 33464
rect 47676 30796 47728 30802
rect 47676 30738 47728 30744
rect 47780 30666 47808 33458
rect 47872 33318 47900 34886
rect 47860 33312 47912 33318
rect 47860 33254 47912 33260
rect 47952 32428 48004 32434
rect 47952 32370 48004 32376
rect 47964 32065 47992 32370
rect 47950 32056 48006 32065
rect 47950 31991 48006 32000
rect 47768 30660 47820 30666
rect 47768 30602 47820 30608
rect 47780 30394 47808 30602
rect 47768 30388 47820 30394
rect 47768 30330 47820 30336
rect 47952 29504 48004 29510
rect 47952 29446 48004 29452
rect 47768 27872 47820 27878
rect 47768 27814 47820 27820
rect 47780 27606 47808 27814
rect 47768 27600 47820 27606
rect 47768 27542 47820 27548
rect 47768 25696 47820 25702
rect 47768 25638 47820 25644
rect 47584 24812 47636 24818
rect 47584 24754 47636 24760
rect 47492 24404 47544 24410
rect 47492 24346 47544 24352
rect 47596 24290 47624 24754
rect 47780 24342 47808 25638
rect 47504 24262 47624 24290
rect 47768 24336 47820 24342
rect 47768 24278 47820 24284
rect 47504 23798 47532 24262
rect 47584 24064 47636 24070
rect 47584 24006 47636 24012
rect 47492 23792 47544 23798
rect 47492 23734 47544 23740
rect 47400 23588 47452 23594
rect 47400 23530 47452 23536
rect 47136 20318 47348 20346
rect 47032 19984 47084 19990
rect 47032 19926 47084 19932
rect 46940 19916 46992 19922
rect 46940 19858 46992 19864
rect 46952 19718 46980 19858
rect 46572 19712 46624 19718
rect 46572 19654 46624 19660
rect 46940 19712 46992 19718
rect 46940 19654 46992 19660
rect 46584 19378 46612 19654
rect 46572 19372 46624 19378
rect 46572 19314 46624 19320
rect 46664 19372 46716 19378
rect 46664 19314 46716 19320
rect 46296 17604 46348 17610
rect 46296 17546 46348 17552
rect 46112 16040 46164 16046
rect 46112 15982 46164 15988
rect 46020 11076 46072 11082
rect 46020 11018 46072 11024
rect 46124 6914 46152 15982
rect 46480 14816 46532 14822
rect 46480 14758 46532 14764
rect 46492 13394 46520 14758
rect 46480 13388 46532 13394
rect 46480 13330 46532 13336
rect 46296 12232 46348 12238
rect 46296 12174 46348 12180
rect 46308 11218 46336 12174
rect 46296 11212 46348 11218
rect 46296 11154 46348 11160
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46308 10130 46336 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 46204 7404 46256 7410
rect 46204 7346 46256 7352
rect 46032 6886 46152 6914
rect 45928 5364 45980 5370
rect 45928 5306 45980 5312
rect 45468 4752 45520 4758
rect 45468 4694 45520 4700
rect 45192 3528 45244 3534
rect 46032 3505 46060 6886
rect 46216 4758 46244 7346
rect 46676 6458 46704 19314
rect 47044 18358 47072 19926
rect 47032 18352 47084 18358
rect 47032 18294 47084 18300
rect 46756 18284 46808 18290
rect 46756 18226 46808 18232
rect 46768 17134 46796 18226
rect 46940 17604 46992 17610
rect 46940 17546 46992 17552
rect 46952 17338 46980 17546
rect 46940 17332 46992 17338
rect 46940 17274 46992 17280
rect 47044 17270 47072 18294
rect 47136 17270 47164 20318
rect 47412 20074 47440 23530
rect 47228 20046 47440 20074
rect 47032 17264 47084 17270
rect 47032 17206 47084 17212
rect 47124 17264 47176 17270
rect 47124 17206 47176 17212
rect 47228 17202 47256 20046
rect 47504 19938 47532 23734
rect 47596 22642 47624 24006
rect 47964 23322 47992 29446
rect 47768 23316 47820 23322
rect 47768 23258 47820 23264
rect 47952 23316 48004 23322
rect 47952 23258 48004 23264
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 47596 21690 47624 22578
rect 47780 21842 47808 23258
rect 47860 22568 47912 22574
rect 47860 22510 47912 22516
rect 47688 21814 47808 21842
rect 47584 21684 47636 21690
rect 47584 21626 47636 21632
rect 47688 21554 47716 21814
rect 47872 21554 47900 22510
rect 47950 21856 48006 21865
rect 47950 21791 48006 21800
rect 47676 21548 47728 21554
rect 47676 21490 47728 21496
rect 47860 21548 47912 21554
rect 47860 21490 47912 21496
rect 47768 21480 47820 21486
rect 47768 21422 47820 21428
rect 47780 20058 47808 21422
rect 47768 20052 47820 20058
rect 47768 19994 47820 20000
rect 47412 19910 47532 19938
rect 47412 19854 47440 19910
rect 47400 19848 47452 19854
rect 47400 19790 47452 19796
rect 47216 17196 47268 17202
rect 47216 17138 47268 17144
rect 46756 17128 46808 17134
rect 47228 17082 47256 17138
rect 46756 17070 46808 17076
rect 46768 7954 46796 17070
rect 47136 17054 47256 17082
rect 46848 14340 46900 14346
rect 46848 14282 46900 14288
rect 46860 8265 46888 14282
rect 47136 10674 47164 17054
rect 47216 16788 47268 16794
rect 47216 16730 47268 16736
rect 47124 10668 47176 10674
rect 47124 10610 47176 10616
rect 46940 8492 46992 8498
rect 46940 8434 46992 8440
rect 46846 8256 46902 8265
rect 46846 8191 46902 8200
rect 46756 7948 46808 7954
rect 46756 7890 46808 7896
rect 46952 7546 46980 8434
rect 47124 8356 47176 8362
rect 47124 8298 47176 8304
rect 47136 7818 47164 8298
rect 47032 7812 47084 7818
rect 47032 7754 47084 7760
rect 47124 7812 47176 7818
rect 47124 7754 47176 7760
rect 47044 7546 47072 7754
rect 46940 7540 46992 7546
rect 46940 7482 46992 7488
rect 47032 7540 47084 7546
rect 47032 7482 47084 7488
rect 47228 6798 47256 16730
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47320 6866 47348 7511
rect 47308 6860 47360 6866
rect 47308 6802 47360 6808
rect 47216 6792 47268 6798
rect 47216 6734 47268 6740
rect 46664 6452 46716 6458
rect 46664 6394 46716 6400
rect 46204 4752 46256 4758
rect 46204 4694 46256 4700
rect 47412 4690 47440 19790
rect 47492 19712 47544 19718
rect 47492 19654 47544 19660
rect 47504 18834 47532 19654
rect 47492 18828 47544 18834
rect 47492 18770 47544 18776
rect 47492 17740 47544 17746
rect 47492 17682 47544 17688
rect 47504 15706 47532 17682
rect 47676 16992 47728 16998
rect 47676 16934 47728 16940
rect 47688 16522 47716 16934
rect 47872 16794 47900 21490
rect 47964 20534 47992 21791
rect 47952 20528 48004 20534
rect 47952 20470 48004 20476
rect 47952 19916 48004 19922
rect 47952 19858 48004 19864
rect 47964 19666 47992 19858
rect 48056 19786 48084 46310
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 48240 43858 48268 44911
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 48136 41608 48188 41614
rect 48134 41576 48136 41585
rect 48188 41576 48190 41585
rect 48134 41511 48190 41520
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48148 39506 48176 40151
rect 48136 39500 48188 39506
rect 48136 39442 48188 39448
rect 48136 38276 48188 38282
rect 48136 38218 48188 38224
rect 48148 38185 48176 38218
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48136 35692 48188 35698
rect 48136 35634 48188 35640
rect 48148 34785 48176 35634
rect 48228 35080 48280 35086
rect 48228 35022 48280 35028
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48240 34105 48268 35022
rect 48226 34096 48282 34105
rect 48226 34031 48282 34040
rect 48136 32836 48188 32842
rect 48136 32778 48188 32784
rect 48148 32745 48176 32778
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48228 30388 48280 30394
rect 48228 30330 48280 30336
rect 48136 29640 48188 29646
rect 48136 29582 48188 29588
rect 48148 29345 48176 29582
rect 48134 29336 48190 29345
rect 48134 29271 48190 29280
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48134 25936 48190 25945
rect 48134 25871 48190 25880
rect 48148 25362 48176 25871
rect 48136 25356 48188 25362
rect 48136 25298 48188 25304
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48148 24274 48176 24511
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 48136 23112 48188 23118
rect 48136 23054 48188 23060
rect 48148 22234 48176 23054
rect 48136 22228 48188 22234
rect 48136 22170 48188 22176
rect 48148 21690 48176 22170
rect 48136 21684 48188 21690
rect 48136 21626 48188 21632
rect 48134 21448 48190 21457
rect 48134 21383 48136 21392
rect 48188 21383 48190 21392
rect 48136 21354 48188 21360
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48044 19780 48096 19786
rect 48044 19722 48096 19728
rect 47964 19638 48084 19666
rect 47860 16788 47912 16794
rect 47860 16730 47912 16736
rect 47768 16652 47820 16658
rect 47768 16594 47820 16600
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 47780 16114 47808 16594
rect 47768 16108 47820 16114
rect 47768 16050 47820 16056
rect 47492 15700 47544 15706
rect 47492 15642 47544 15648
rect 47768 13728 47820 13734
rect 47768 13670 47820 13676
rect 47780 13462 47808 13670
rect 47768 13456 47820 13462
rect 47768 13398 47820 13404
rect 47492 10668 47544 10674
rect 47492 10610 47544 10616
rect 47400 4684 47452 4690
rect 47400 4626 47452 4632
rect 46848 4616 46900 4622
rect 46848 4558 46900 4564
rect 46480 4480 46532 4486
rect 46480 4422 46532 4428
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46308 3602 46336 3878
rect 46492 3602 46520 4422
rect 46664 4208 46716 4214
rect 46860 4185 46888 4558
rect 46664 4150 46716 4156
rect 46846 4176 46902 4185
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 46676 3505 46704 4150
rect 46846 4111 46902 4120
rect 45192 3470 45244 3476
rect 46018 3496 46074 3505
rect 45204 3058 45232 3470
rect 46018 3431 46074 3440
rect 46662 3496 46718 3505
rect 47504 3466 47532 10610
rect 47676 10464 47728 10470
rect 47676 10406 47728 10412
rect 47688 10130 47716 10406
rect 47676 10124 47728 10130
rect 47676 10066 47728 10072
rect 47858 9616 47914 9625
rect 47858 9551 47860 9560
rect 47912 9551 47914 9560
rect 47860 9522 47912 9528
rect 47766 8936 47822 8945
rect 47766 8871 47768 8880
rect 47820 8871 47822 8880
rect 47768 8842 47820 8848
rect 47952 6316 48004 6322
rect 47952 6258 48004 6264
rect 47964 6225 47992 6258
rect 47950 6216 48006 6225
rect 47950 6151 48006 6160
rect 47768 4208 47820 4214
rect 47768 4150 47820 4156
rect 46662 3431 46718 3440
rect 47492 3460 47544 3466
rect 47492 3402 47544 3408
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45388 3126 45416 3334
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 46756 3052 46808 3058
rect 46756 2994 46808 3000
rect 46388 2372 46440 2378
rect 46388 2314 46440 2320
rect 45468 2304 45520 2310
rect 45468 2246 45520 2252
rect 45480 2038 45508 2246
rect 45468 2032 45520 2038
rect 45468 1974 45520 1980
rect 46400 800 46428 2314
rect 18892 734 19104 762
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46768 105 46796 2994
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 47044 800 47072 2382
rect 47688 800 47716 2926
rect 47780 1465 47808 4150
rect 47860 3936 47912 3942
rect 47860 3878 47912 3884
rect 47872 3670 47900 3878
rect 47860 3664 47912 3670
rect 47860 3606 47912 3612
rect 48056 2650 48084 19638
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48148 18834 48176 19071
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 48136 17604 48188 17610
rect 48136 17546 48188 17552
rect 48148 17105 48176 17546
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48136 16516 48188 16522
rect 48136 16458 48188 16464
rect 48148 16425 48176 16458
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48136 13252 48188 13258
rect 48136 13194 48188 13200
rect 48148 12345 48176 13194
rect 48134 12336 48190 12345
rect 48134 12271 48190 12280
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 48240 9450 48268 30330
rect 48228 9444 48280 9450
rect 48228 9386 48280 9392
rect 48136 7404 48188 7410
rect 48136 7346 48188 7352
rect 48148 6905 48176 7346
rect 48134 6896 48190 6905
rect 48134 6831 48190 6840
rect 48320 5228 48372 5234
rect 48320 5170 48372 5176
rect 48044 2644 48096 2650
rect 48044 2586 48096 2592
rect 48044 2372 48096 2378
rect 48044 2314 48096 2320
rect 47766 1456 47822 1465
rect 47766 1391 47822 1400
rect 46754 96 46810 105
rect 46754 31 46810 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48056 785 48084 2314
rect 48332 800 48360 5170
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48976 800 49004 3402
rect 48042 776 48098 785
rect 48042 711 48098 720
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1858 47640 1914 47696
rect 1398 42880 1454 42936
rect 1582 35400 1638 35456
rect 1398 33396 1400 33416
rect 1400 33396 1452 33416
rect 1452 33396 1454 33416
rect 1398 33360 1454 33396
rect 1582 32680 1638 32736
rect 1858 41520 1914 41576
rect 1858 40160 1914 40216
rect 3422 46960 3478 47016
rect 2778 46280 2834 46336
rect 2778 36760 2834 36816
rect 3238 32000 3294 32056
rect 1858 25220 1914 25256
rect 1858 25200 1860 25220
rect 1860 25200 1912 25220
rect 1912 25200 1914 25220
rect 1858 23160 1914 23216
rect 1398 17720 1454 17776
rect 1858 16360 1914 16416
rect 1398 12280 1454 12336
rect 2226 19080 2282 19136
rect 3330 28600 3386 28656
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3514 44920 3570 44976
rect 3698 43560 3754 43616
rect 3606 31320 3662 31376
rect 3882 39480 3938 39536
rect 3514 19760 3570 19816
rect 3422 18400 3478 18456
rect 3054 17040 3110 17096
rect 2778 15000 2834 15056
rect 3422 13640 3478 13696
rect 3146 10240 3202 10296
rect 3146 7520 3202 7576
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3422 6860 3478 6896
rect 3422 6840 3424 6860
rect 3424 6840 3476 6860
rect 3476 6840 3478 6860
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 2962 3440 3018 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4066 1400 4122 1456
rect 10322 21020 10324 21040
rect 10324 21020 10376 21040
rect 10376 21020 10378 21040
rect 10322 20984 10378 21020
rect 14370 21020 14372 21040
rect 14372 21020 14424 21040
rect 14424 21020 14426 21040
rect 14370 20984 14426 21020
rect 14002 20848 14058 20904
rect 12806 20304 12862 20360
rect 14462 20304 14518 20360
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19522 33360 19578 33416
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19430 31184 19486 31240
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 20074 31184 20130 31240
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19982 22616 20038 22672
rect 18418 20848 18474 20904
rect 17406 3440 17462 3496
rect 17682 3032 17738 3088
rect 2778 720 2834 776
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19982 20476 19984 20496
rect 19984 20476 20036 20496
rect 20036 20476 20038 20496
rect 19982 20440 20038 20476
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19982 2896 20038 2952
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20166 3032 20222 3088
rect 20994 29008 21050 29064
rect 20626 3984 20682 4040
rect 20626 2896 20682 2952
rect 22098 26832 22154 26888
rect 22558 29008 22614 29064
rect 22558 28872 22614 28928
rect 23386 31864 23442 31920
rect 21730 21528 21786 21584
rect 22466 22636 22522 22672
rect 22466 22616 22468 22636
rect 22468 22616 22520 22636
rect 22520 22616 22522 22636
rect 22466 21936 22522 21992
rect 23110 21972 23112 21992
rect 23112 21972 23164 21992
rect 23164 21972 23166 21992
rect 23110 21936 23166 21972
rect 25686 26968 25742 27024
rect 25870 26832 25926 26888
rect 26330 26968 26386 27024
rect 22006 3032 22062 3088
rect 23478 3068 23480 3088
rect 23480 3068 23532 3088
rect 23532 3068 23534 3088
rect 23478 3032 23534 3068
rect 26974 31184 27030 31240
rect 27618 28872 27674 28928
rect 28630 33360 28686 33416
rect 26238 21936 26294 21992
rect 28446 21528 28502 21584
rect 26974 3984 27030 4040
rect 27158 3984 27214 4040
rect 30010 32272 30066 32328
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 30746 31900 30748 31920
rect 30748 31900 30800 31920
rect 30800 31900 30802 31920
rect 30746 31864 30802 31900
rect 31482 32272 31538 32328
rect 32218 20596 32274 20632
rect 32218 20576 32220 20596
rect 32220 20576 32272 20596
rect 32272 20576 32274 20596
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35254 20576 35310 20632
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 39762 21392 39818 21448
rect 41694 21548 41750 21584
rect 41694 21528 41696 21548
rect 41696 21528 41748 21548
rect 41748 21528 41750 21548
rect 46846 47640 46902 47696
rect 46478 46960 46534 47016
rect 46662 39480 46718 39536
rect 45650 29960 45706 30016
rect 45558 28600 45614 28656
rect 45742 26560 45798 26616
rect 45558 23840 45614 23896
rect 45926 23160 45982 23216
rect 43626 21548 43682 21584
rect 43626 21528 43628 21548
rect 43628 21528 43680 21548
rect 43680 21528 43682 21548
rect 46478 31320 46534 31376
rect 46202 22516 46204 22536
rect 46204 22516 46256 22536
rect 46256 22516 46258 22536
rect 46202 22480 46258 22516
rect 45558 15680 45614 15736
rect 45834 18400 45890 18456
rect 46846 33360 46902 33416
rect 46846 25200 46902 25256
rect 46386 20440 46442 20496
rect 47950 46280 48006 46336
rect 47950 40840 48006 40896
rect 47858 38800 47914 38856
rect 47950 32000 48006 32056
rect 47950 21800 48006 21856
rect 46846 8200 46902 8256
rect 47306 7520 47362 7576
rect 48134 45600 48190 45656
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 48134 41556 48136 41576
rect 48136 41556 48188 41576
rect 48188 41556 48190 41576
rect 48134 41520 48190 41556
rect 48134 40160 48190 40216
rect 48134 38120 48190 38176
rect 48134 34720 48190 34776
rect 48226 34040 48282 34096
rect 48134 32680 48190 32736
rect 48134 29280 48190 29336
rect 48134 27920 48190 27976
rect 48134 25880 48190 25936
rect 48134 24520 48190 24576
rect 48134 21412 48190 21448
rect 48134 21392 48136 21412
rect 48136 21392 48188 21412
rect 48188 21392 48190 21412
rect 48134 21120 48190 21176
rect 46846 4120 46902 4176
rect 46018 3440 46074 3496
rect 46662 3440 46718 3496
rect 47858 9580 47914 9616
rect 47858 9560 47860 9580
rect 47860 9560 47912 9580
rect 47912 9560 47914 9580
rect 47766 8900 47822 8936
rect 47766 8880 47768 8900
rect 47768 8880 47820 8900
rect 47820 8880 47822 8900
rect 47950 6160 48006 6216
rect 48134 19080 48190 19136
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 12280 48190 12336
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 48134 6840 48190 6896
rect 47766 1400 47822 1456
rect 46754 40 46810 96
rect 48042 720 48098 776
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1853 47698 1919 47701
rect 0 47696 1919 47698
rect 0 47640 1858 47696
rect 1914 47640 1919 47696
rect 0 47638 1919 47640
rect 0 47548 800 47638
rect 1853 47635 1919 47638
rect 46841 47698 46907 47701
rect 49200 47698 50000 47788
rect 46841 47696 50000 47698
rect 46841 47640 46846 47696
rect 46902 47640 50000 47696
rect 46841 47638 50000 47640
rect 46841 47635 46907 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3417 47018 3483 47021
rect 0 47016 3483 47018
rect 0 46960 3422 47016
rect 3478 46960 3483 47016
rect 0 46958 3483 46960
rect 0 46868 800 46958
rect 3417 46955 3483 46958
rect 46473 47018 46539 47021
rect 49200 47018 50000 47108
rect 46473 47016 50000 47018
rect 46473 46960 46478 47016
rect 46534 46960 50000 47016
rect 46473 46958 50000 46960
rect 46473 46955 46539 46958
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46188 800 46278
rect 2773 46275 2839 46278
rect 47945 46338 48011 46341
rect 49200 46338 50000 46428
rect 47945 46336 50000 46338
rect 47945 46280 47950 46336
rect 48006 46280 50000 46336
rect 47945 46278 50000 46280
rect 47945 46275 48011 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3509 44978 3575 44981
rect 0 44976 3575 44978
rect 0 44920 3514 44976
rect 3570 44920 3575 44976
rect 0 44918 3575 44920
rect 0 44828 800 44918
rect 3509 44915 3575 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3693 43618 3759 43621
rect 0 43616 3759 43618
rect 0 43560 3698 43616
rect 3754 43560 3759 43616
rect 0 43558 3759 43560
rect 0 43468 800 43558
rect 3693 43555 3759 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42788 800 42878
rect 1393 42875 1459 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 47945 40898 48011 40901
rect 49200 40898 50000 40988
rect 47945 40896 50000 40898
rect 47945 40840 47950 40896
rect 48006 40840 50000 40896
rect 47945 40838 50000 40840
rect 47945 40835 48011 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1853 40218 1919 40221
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40068 800 40158
rect 1853 40155 1919 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40308
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3877 39538 3943 39541
rect 0 39536 3943 39538
rect 0 39480 3882 39536
rect 3938 39480 3943 39536
rect 0 39478 3943 39480
rect 0 39388 800 39478
rect 3877 39475 3943 39478
rect 46657 39538 46723 39541
rect 49200 39538 50000 39628
rect 46657 39536 50000 39538
rect 46657 39480 46662 39536
rect 46718 39480 50000 39536
rect 46657 39478 50000 39480
rect 46657 39475 46723 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47853 38858 47919 38861
rect 49200 38858 50000 38948
rect 47853 38856 50000 38858
rect 47853 38800 47858 38856
rect 47914 38800 50000 38856
rect 47853 38798 50000 38800
rect 47853 38795 47919 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35458 800 35548
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 48221 34098 48287 34101
rect 49200 34098 50000 34188
rect 48221 34096 50000 34098
rect 48221 34040 48226 34096
rect 48282 34040 50000 34096
rect 48221 34038 50000 34040
rect 48221 34035 48287 34038
rect 49200 33948 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 19517 33418 19583 33421
rect 28625 33418 28691 33421
rect 19517 33416 28691 33418
rect 19517 33360 19522 33416
rect 19578 33360 28630 33416
rect 28686 33360 28691 33416
rect 19517 33358 28691 33360
rect 19517 33355 19583 33358
rect 28625 33355 28691 33358
rect 46841 33418 46907 33421
rect 49200 33418 50000 33508
rect 46841 33416 50000 33418
rect 46841 33360 46846 33416
rect 46902 33360 50000 33416
rect 46841 33358 50000 33360
rect 46841 33355 46907 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32828
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32588 800 32678
rect 1577 32675 1643 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 49200 32588 50000 32678
rect 30005 32330 30071 32333
rect 31477 32330 31543 32333
rect 30005 32328 31543 32330
rect 30005 32272 30010 32328
rect 30066 32272 31482 32328
rect 31538 32272 31543 32328
rect 30005 32270 31543 32272
rect 30005 32267 30071 32270
rect 31477 32267 31543 32270
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 3233 32058 3299 32061
rect 0 32056 3299 32058
rect 0 32000 3238 32056
rect 3294 32000 3299 32056
rect 0 31998 3299 32000
rect 0 31908 800 31998
rect 3233 31995 3299 31998
rect 47945 32058 48011 32061
rect 49200 32058 50000 32148
rect 47945 32056 50000 32058
rect 47945 32000 47950 32056
rect 48006 32000 50000 32056
rect 47945 31998 50000 32000
rect 47945 31995 48011 31998
rect 23381 31922 23447 31925
rect 30741 31922 30807 31925
rect 23381 31920 30807 31922
rect 23381 31864 23386 31920
rect 23442 31864 30746 31920
rect 30802 31864 30807 31920
rect 49200 31908 50000 31998
rect 23381 31862 30807 31864
rect 23381 31859 23447 31862
rect 30741 31859 30807 31862
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3601 31378 3667 31381
rect 0 31376 3667 31378
rect 0 31320 3606 31376
rect 3662 31320 3667 31376
rect 0 31318 3667 31320
rect 0 31228 800 31318
rect 3601 31315 3667 31318
rect 46473 31378 46539 31381
rect 49200 31378 50000 31468
rect 46473 31376 50000 31378
rect 46473 31320 46478 31376
rect 46534 31320 50000 31376
rect 46473 31318 50000 31320
rect 46473 31315 46539 31318
rect 19425 31242 19491 31245
rect 20069 31242 20135 31245
rect 26969 31242 27035 31245
rect 19425 31240 27035 31242
rect 19425 31184 19430 31240
rect 19486 31184 20074 31240
rect 20130 31184 26974 31240
rect 27030 31184 27035 31240
rect 49200 31228 50000 31318
rect 19425 31182 27035 31184
rect 19425 31179 19491 31182
rect 20069 31179 20135 31182
rect 26969 31179 27035 31182
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 29868 800 30108
rect 45645 30018 45711 30021
rect 49200 30018 50000 30108
rect 45645 30016 50000 30018
rect 45645 29960 45650 30016
rect 45706 29960 50000 30016
rect 45645 29958 50000 29960
rect 45645 29955 45711 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 48129 29338 48195 29341
rect 49200 29338 50000 29428
rect 48129 29336 50000 29338
rect 48129 29280 48134 29336
rect 48190 29280 50000 29336
rect 48129 29278 50000 29280
rect 48129 29275 48195 29278
rect 49200 29188 50000 29278
rect 20989 29066 21055 29069
rect 22553 29066 22619 29069
rect 20989 29064 22619 29066
rect 20989 29008 20994 29064
rect 21050 29008 22558 29064
rect 22614 29008 22619 29064
rect 20989 29006 22619 29008
rect 20989 29003 21055 29006
rect 22553 29003 22619 29006
rect 22553 28930 22619 28933
rect 27613 28930 27679 28933
rect 22553 28928 27679 28930
rect 22553 28872 22558 28928
rect 22614 28872 27618 28928
rect 27674 28872 27679 28928
rect 22553 28870 27679 28872
rect 22553 28867 22619 28870
rect 27613 28867 27679 28870
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3325 28658 3391 28661
rect 0 28656 3391 28658
rect 0 28600 3330 28656
rect 3386 28600 3391 28656
rect 0 28598 3391 28600
rect 0 28508 800 28598
rect 3325 28595 3391 28598
rect 45553 28658 45619 28661
rect 49200 28658 50000 28748
rect 45553 28656 50000 28658
rect 45553 28600 45558 28656
rect 45614 28600 50000 28656
rect 45553 28598 50000 28600
rect 45553 28595 45619 28598
rect 49200 28508 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 49200 27828 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 25681 27026 25747 27029
rect 26325 27026 26391 27029
rect 25681 27024 26391 27026
rect 25681 26968 25686 27024
rect 25742 26968 26330 27024
rect 26386 26968 26391 27024
rect 25681 26966 26391 26968
rect 25681 26963 25747 26966
rect 26325 26963 26391 26966
rect 22093 26890 22159 26893
rect 25865 26890 25931 26893
rect 22093 26888 25931 26890
rect 22093 26832 22098 26888
rect 22154 26832 25870 26888
rect 25926 26832 25931 26888
rect 22093 26830 25931 26832
rect 22093 26827 22159 26830
rect 25865 26827 25931 26830
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 45737 26618 45803 26621
rect 49200 26618 50000 26708
rect 45737 26616 50000 26618
rect 45737 26560 45742 26616
rect 45798 26560 50000 26616
rect 45737 26558 50000 26560
rect 45737 26555 45803 26558
rect 49200 26468 50000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 48129 25938 48195 25941
rect 49200 25938 50000 26028
rect 48129 25936 50000 25938
rect 48129 25880 48134 25936
rect 48190 25880 50000 25936
rect 48129 25878 50000 25880
rect 48129 25875 48195 25878
rect 49200 25788 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25108 800 25198
rect 1853 25195 1919 25198
rect 46841 25258 46907 25261
rect 49200 25258 50000 25348
rect 46841 25256 50000 25258
rect 46841 25200 46846 25256
rect 46902 25200 50000 25256
rect 46841 25198 50000 25200
rect 46841 25195 46907 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24428 800 24668
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 45553 23898 45619 23901
rect 49200 23898 50000 23988
rect 45553 23896 50000 23898
rect 45553 23840 45558 23896
rect 45614 23840 50000 23896
rect 45553 23838 50000 23840
rect 45553 23835 45619 23838
rect 49200 23748 50000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23068 800 23158
rect 1853 23155 1919 23158
rect 45921 23218 45987 23221
rect 49200 23218 50000 23308
rect 45921 23216 50000 23218
rect 45921 23160 45926 23216
rect 45982 23160 50000 23216
rect 45921 23158 50000 23160
rect 45921 23155 45987 23158
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 19977 22674 20043 22677
rect 22461 22674 22527 22677
rect 19977 22672 22527 22674
rect 0 22388 800 22628
rect 19977 22616 19982 22672
rect 20038 22616 22466 22672
rect 22522 22616 22527 22672
rect 19977 22614 22527 22616
rect 19977 22611 20043 22614
rect 22461 22611 22527 22614
rect 46197 22538 46263 22541
rect 49200 22538 50000 22628
rect 46197 22536 50000 22538
rect 46197 22480 46202 22536
rect 46258 22480 50000 22536
rect 46197 22478 50000 22480
rect 46197 22475 46263 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 22461 21994 22527 21997
rect 23105 21994 23171 21997
rect 26233 21994 26299 21997
rect 22461 21992 26299 21994
rect 0 21708 800 21948
rect 22461 21936 22466 21992
rect 22522 21936 23110 21992
rect 23166 21936 26238 21992
rect 26294 21936 26299 21992
rect 22461 21934 26299 21936
rect 22461 21931 22527 21934
rect 23105 21931 23171 21934
rect 26233 21931 26299 21934
rect 47945 21858 48011 21861
rect 49200 21858 50000 21948
rect 47945 21856 50000 21858
rect 47945 21800 47950 21856
rect 48006 21800 50000 21856
rect 47945 21798 50000 21800
rect 47945 21795 48011 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 21725 21586 21791 21589
rect 28441 21586 28507 21589
rect 21725 21584 28507 21586
rect 21725 21528 21730 21584
rect 21786 21528 28446 21584
rect 28502 21528 28507 21584
rect 21725 21526 28507 21528
rect 21725 21523 21791 21526
rect 28441 21523 28507 21526
rect 41689 21586 41755 21589
rect 43621 21586 43687 21589
rect 41689 21584 43687 21586
rect 41689 21528 41694 21584
rect 41750 21528 43626 21584
rect 43682 21528 43687 21584
rect 41689 21526 43687 21528
rect 41689 21523 41755 21526
rect 43621 21523 43687 21526
rect 39757 21450 39823 21453
rect 48129 21450 48195 21453
rect 39757 21448 48195 21450
rect 39757 21392 39762 21448
rect 39818 21392 48134 21448
rect 48190 21392 48195 21448
rect 39757 21390 48195 21392
rect 39757 21387 39823 21390
rect 48129 21387 48195 21390
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 10317 21042 10383 21045
rect 14365 21042 14431 21045
rect 10317 21040 14431 21042
rect 10317 20984 10322 21040
rect 10378 20984 14370 21040
rect 14426 20984 14431 21040
rect 49200 21028 50000 21118
rect 10317 20982 14431 20984
rect 10317 20979 10383 20982
rect 14365 20979 14431 20982
rect 13997 20906 14063 20909
rect 18413 20906 18479 20909
rect 13997 20904 18479 20906
rect 13997 20848 14002 20904
rect 14058 20848 18418 20904
rect 18474 20848 18479 20904
rect 13997 20846 18479 20848
rect 13997 20843 14063 20846
rect 18413 20843 18479 20846
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 32213 20634 32279 20637
rect 35249 20634 35315 20637
rect 32213 20632 35315 20634
rect 0 20348 800 20588
rect 32213 20576 32218 20632
rect 32274 20576 35254 20632
rect 35310 20576 35315 20632
rect 32213 20574 35315 20576
rect 32213 20571 32279 20574
rect 35249 20571 35315 20574
rect 19977 20498 20043 20501
rect 46381 20498 46447 20501
rect 19977 20496 46447 20498
rect 19977 20440 19982 20496
rect 20038 20440 46386 20496
rect 46442 20440 46447 20496
rect 19977 20438 46447 20440
rect 19977 20435 20043 20438
rect 46381 20435 46447 20438
rect 12801 20362 12867 20365
rect 14457 20362 14523 20365
rect 12801 20360 14523 20362
rect 12801 20304 12806 20360
rect 12862 20304 14462 20360
rect 14518 20304 14523 20360
rect 12801 20302 14523 20304
rect 12801 20299 12867 20302
rect 14457 20299 14523 20302
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 3509 19818 3575 19821
rect 0 19816 3575 19818
rect 0 19760 3514 19816
rect 3570 19760 3575 19816
rect 0 19758 3575 19760
rect 0 19668 800 19758
rect 3509 19755 3575 19758
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3417 18458 3483 18461
rect 0 18456 3483 18458
rect 0 18400 3422 18456
rect 3478 18400 3483 18456
rect 0 18398 3483 18400
rect 0 18308 800 18398
rect 3417 18395 3483 18398
rect 45829 18458 45895 18461
rect 49200 18458 50000 18548
rect 45829 18456 50000 18458
rect 45829 18400 45834 18456
rect 45890 18400 50000 18456
rect 45829 18398 50000 18400
rect 45829 18395 45895 18398
rect 49200 18308 50000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17628 800 17718
rect 1393 17715 1459 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3049 17098 3115 17101
rect 0 17096 3115 17098
rect 0 17040 3054 17096
rect 3110 17040 3115 17096
rect 0 17038 3115 17040
rect 0 16948 800 17038
rect 3049 17035 3115 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16268 800 16358
rect 1853 16355 1919 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16508
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 45553 15738 45619 15741
rect 49200 15738 50000 15828
rect 45553 15736 50000 15738
rect 45553 15680 45558 15736
rect 45614 15680 50000 15736
rect 45553 15678 50000 15680
rect 45553 15675 45619 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3417 13698 3483 13701
rect 0 13696 3483 13698
rect 0 13640 3422 13696
rect 3478 13640 3483 13696
rect 0 13638 3483 13640
rect 0 13548 800 13638
rect 3417 13635 3483 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 3141 10298 3207 10301
rect 0 10296 3207 10298
rect 0 10240 3146 10296
rect 3202 10240 3207 10296
rect 0 10238 3207 10240
rect 0 10148 800 10238
rect 3141 10235 3207 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 47853 9618 47919 9621
rect 49200 9618 50000 9708
rect 47853 9616 50000 9618
rect 47853 9560 47858 9616
rect 47914 9560 50000 9616
rect 47853 9558 50000 9560
rect 47853 9555 47919 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47761 8938 47827 8941
rect 49200 8938 50000 9028
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 46841 8258 46907 8261
rect 49200 8258 50000 8348
rect 46841 8256 50000 8258
rect 46841 8200 46846 8256
rect 46902 8200 50000 8256
rect 46841 8198 50000 8200
rect 46841 8195 46907 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3141 7578 3207 7581
rect 0 7576 3207 7578
rect 0 7520 3146 7576
rect 3202 7520 3207 7576
rect 0 7518 3207 7520
rect 0 7428 800 7518
rect 3141 7515 3207 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 3417 6898 3483 6901
rect 0 6896 3483 6898
rect 0 6840 3422 6896
rect 3478 6840 3483 6896
rect 0 6838 3483 6840
rect 0 6748 800 6838
rect 3417 6835 3483 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 47945 6218 48011 6221
rect 49200 6218 50000 6308
rect 47945 6216 50000 6218
rect 47945 6160 47950 6216
rect 48006 6160 50000 6216
rect 47945 6158 50000 6160
rect 47945 6155 48011 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 46841 4178 46907 4181
rect 49200 4178 50000 4268
rect 46841 4176 50000 4178
rect 46841 4120 46846 4176
rect 46902 4120 50000 4176
rect 46841 4118 50000 4120
rect 46841 4115 46907 4118
rect 20621 4042 20687 4045
rect 26969 4042 27035 4045
rect 27153 4042 27219 4045
rect 20621 4040 27219 4042
rect 20621 3984 20626 4040
rect 20682 3984 26974 4040
rect 27030 3984 27158 4040
rect 27214 3984 27219 4040
rect 49200 4028 50000 4118
rect 20621 3982 27219 3984
rect 20621 3979 20687 3982
rect 26969 3979 27035 3982
rect 27153 3979 27219 3982
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3588
rect 2957 3498 3023 3501
rect 0 3496 3023 3498
rect 0 3440 2962 3496
rect 3018 3440 3023 3496
rect 0 3438 3023 3440
rect 0 3348 800 3438
rect 2957 3435 3023 3438
rect 17401 3498 17467 3501
rect 46013 3498 46079 3501
rect 17401 3496 46079 3498
rect 17401 3440 17406 3496
rect 17462 3440 46018 3496
rect 46074 3440 46079 3496
rect 17401 3438 46079 3440
rect 17401 3435 17467 3438
rect 46013 3435 46079 3438
rect 46657 3498 46723 3501
rect 49200 3498 50000 3588
rect 46657 3496 50000 3498
rect 46657 3440 46662 3496
rect 46718 3440 50000 3496
rect 46657 3438 50000 3440
rect 46657 3435 46723 3438
rect 49200 3348 50000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 17677 3090 17743 3093
rect 20161 3090 20227 3093
rect 17677 3088 20227 3090
rect 17677 3032 17682 3088
rect 17738 3032 20166 3088
rect 20222 3032 20227 3088
rect 17677 3030 20227 3032
rect 17677 3027 17743 3030
rect 20161 3027 20227 3030
rect 22001 3090 22067 3093
rect 23473 3090 23539 3093
rect 22001 3088 23539 3090
rect 22001 3032 22006 3088
rect 22062 3032 23478 3088
rect 23534 3032 23539 3088
rect 22001 3030 23539 3032
rect 22001 3027 22067 3030
rect 23473 3027 23539 3030
rect 19977 2954 20043 2957
rect 20621 2954 20687 2957
rect 19977 2952 20687 2954
rect 0 2668 800 2908
rect 19977 2896 19982 2952
rect 20038 2896 20626 2952
rect 20682 2896 20687 2952
rect 19977 2894 20687 2896
rect 19977 2891 20043 2894
rect 20621 2891 20687 2894
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 4061 1458 4127 1461
rect 0 1456 4127 1458
rect 0 1400 4066 1456
rect 4122 1400 4127 1456
rect 0 1398 4127 1400
rect 0 1308 800 1398
rect 4061 1395 4127 1398
rect 47761 1458 47827 1461
rect 49200 1458 50000 1548
rect 47761 1456 50000 1458
rect 47761 1400 47766 1456
rect 47822 1400 50000 1456
rect 47761 1398 50000 1400
rect 47761 1395 47827 1398
rect 49200 1308 50000 1398
rect 0 778 800 868
rect 2773 778 2839 781
rect 0 776 2839 778
rect 0 720 2778 776
rect 2834 720 2839 776
rect 0 718 2839 720
rect 0 628 800 718
rect 2773 715 2839 718
rect 48037 778 48103 781
rect 49200 778 50000 868
rect 48037 776 50000 778
rect 48037 720 48042 776
rect 48098 720 50000 776
rect 48037 718 50000 720
rect 48037 715 48103 718
rect 49200 628 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 188
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 24564 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 45816 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 29900 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform -1 0 35604 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 41676 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 36708 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform 1 0 32200 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1644511149
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1644511149
transform 1 0 15456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_185
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_200
timestamp 1644511149
transform 1 0 19504 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_212
timestamp 1644511149
transform 1 0 20608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_269
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_287
timestamp 1644511149
transform 1 0 27508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_295
timestamp 1644511149
transform 1 0 28244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_314
timestamp 1644511149
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1644511149
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1644511149
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_430
timestamp 1644511149
transform 1 0 40664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1644511149
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1644511149
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_65
timestamp 1644511149
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1644511149
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_91
timestamp 1644511149
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_95
timestamp 1644511149
transform 1 0 9844 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_103
timestamp 1644511149
transform 1 0 10580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1644511149
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1644511149
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_135
timestamp 1644511149
transform 1 0 13524 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 1644511149
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1644511149
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_189
timestamp 1644511149
transform 1 0 18492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_197
timestamp 1644511149
transform 1 0 19228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1644511149
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_228
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_235
timestamp 1644511149
transform 1 0 22724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_239
timestamp 1644511149
transform 1 0 23092 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_269
timestamp 1644511149
transform 1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_294
timestamp 1644511149
transform 1 0 28152 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_306
timestamp 1644511149
transform 1 0 29256 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_318
timestamp 1644511149
transform 1 0 30360 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_330
timestamp 1644511149
transform 1 0 31464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_345
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1644511149
transform 1 0 35972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_413
timestamp 1644511149
transform 1 0 39100 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1644511149
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_436
timestamp 1644511149
transform 1 0 41216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_443
timestamp 1644511149
transform 1 0 41860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_470
timestamp 1644511149
transform 1 0 44344 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_52
timestamp 1644511149
transform 1 0 5888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1644511149
transform 1 0 6256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_63
timestamp 1644511149
transform 1 0 6900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_70
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1644511149
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_95
timestamp 1644511149
transform 1 0 9844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1644511149
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_151
timestamp 1644511149
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_158
timestamp 1644511149
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_186
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1644511149
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1644511149
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_216
timestamp 1644511149
transform 1 0 20976 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_222
timestamp 1644511149
transform 1 0 21528 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_239
timestamp 1644511149
transform 1 0 23092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_246
timestamp 1644511149
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_284
timestamp 1644511149
transform 1 0 27232 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_296
timestamp 1644511149
transform 1 0 28336 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_350
timestamp 1644511149
transform 1 0 33304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_426
timestamp 1644511149
transform 1 0 40296 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_455
timestamp 1644511149
transform 1 0 42964 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_462
timestamp 1644511149
transform 1 0 43608 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_65
timestamp 1644511149
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_120
timestamp 1644511149
transform 1 0 12144 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1644511149
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1644511149
transform 1 0 14168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1644511149
transform 1 0 15456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1644511149
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1644511149
transform 1 0 17572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_186
timestamp 1644511149
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1644511149
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_214
timestamp 1644511149
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1644511149
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_234
timestamp 1644511149
transform 1 0 22632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_238
timestamp 1644511149
transform 1 0 23000 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_253
timestamp 1644511149
transform 1 0 24380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_260
timestamp 1644511149
transform 1 0 25024 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_267
timestamp 1644511149
transform 1 0 25668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_294
timestamp 1644511149
transform 1 0 28152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_306
timestamp 1644511149
transform 1 0 29256 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_318
timestamp 1644511149
transform 1 0 30360 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1644511149
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_399
timestamp 1644511149
transform 1 0 37812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_411
timestamp 1644511149
transform 1 0 38916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_422
timestamp 1644511149
transform 1 0 39928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_431
timestamp 1644511149
transform 1 0 40756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_438
timestamp 1644511149
transform 1 0 41400 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_446
timestamp 1644511149
transform 1 0 42136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_455
timestamp 1644511149
transform 1 0 42964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_467
timestamp 1644511149
transform 1 0 44068 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_479
timestamp 1644511149
transform 1 0 45172 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_490
timestamp 1644511149
transform 1 0 46184 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_146
timestamp 1644511149
transform 1 0 14536 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_158
timestamp 1644511149
transform 1 0 15640 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_170
timestamp 1644511149
transform 1 0 16744 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_182
timestamp 1644511149
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_186
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_190
timestamp 1644511149
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1644511149
transform 1 0 20884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1644511149
transform 1 0 21988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1644511149
transform 1 0 23092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_394
timestamp 1644511149
transform 1 0 37352 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_406
timestamp 1644511149
transform 1 0 38456 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_412
timestamp 1644511149
transform 1 0 39008 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_416
timestamp 1644511149
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_443
timestamp 1644511149
transform 1 0 41860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_449
timestamp 1644511149
transform 1 0 42412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_463
timestamp 1644511149
transform 1 0 43700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_498
timestamp 1644511149
transform 1 0 46920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_409
timestamp 1644511149
transform 1 0 38732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_423
timestamp 1644511149
transform 1 0 40020 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_430
timestamp 1644511149
transform 1 0 40664 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_442
timestamp 1644511149
transform 1 0 41768 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_452
timestamp 1644511149
transform 1 0 42688 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_464
timestamp 1644511149
transform 1 0 43792 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_476
timestamp 1644511149
transform 1 0 44896 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_488
timestamp 1644511149
transform 1 0 46000 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1644511149
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_385
timestamp 1644511149
transform 1 0 36524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_404
timestamp 1644511149
transform 1 0 38272 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_416
timestamp 1644511149
transform 1 0 39376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_443
timestamp 1644511149
transform 1 0 41860 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_458
timestamp 1644511149
transform 1 0 43240 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_470
timestamp 1644511149
transform 1 0 44344 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1644511149
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_488
timestamp 1644511149
transform 1 0 46000 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_496
timestamp 1644511149
transform 1 0 46736 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1644511149
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_494
timestamp 1644511149
transform 1 0 46552 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_511
timestamp 1644511149
transform 1 0 48116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_515
timestamp 1644511149
transform 1 0 48484 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_493
timestamp 1644511149
transform 1 0 46460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_499
timestamp 1644511149
transform 1 0 47012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1644511149
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_505
timestamp 1644511149
transform 1 0 47564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_512
timestamp 1644511149
transform 1 0 48208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_232
timestamp 1644511149
transform 1 0 22448 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1644511149
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1644511149
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_507
timestamp 1644511149
transform 1 0 47748 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_515
timestamp 1644511149
transform 1 0 48484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1644511149
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1644511149
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_172
timestamp 1644511149
transform 1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_180
timestamp 1644511149
transform 1 0 17664 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1644511149
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1644511149
transform 1 0 19596 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_213
timestamp 1644511149
transform 1 0 20700 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1644511149
transform 1 0 21252 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1644511149
transform 1 0 21988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1644511149
transform 1 0 23092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_317
timestamp 1644511149
transform 1 0 30268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_339
timestamp 1644511149
transform 1 0 32292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_351
timestamp 1644511149
transform 1 0 33396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_155
timestamp 1644511149
transform 1 0 15364 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1644511149
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_177
timestamp 1644511149
transform 1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_202
timestamp 1644511149
transform 1 0 19688 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_214
timestamp 1644511149
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1644511149
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_246
timestamp 1644511149
transform 1 0 23736 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1644511149
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_258
timestamp 1644511149
transform 1 0 24840 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_262
timestamp 1644511149
transform 1 0 25208 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1644511149
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_477
timestamp 1644511149
transform 1 0 44988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_481
timestamp 1644511149
transform 1 0 45356 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_493
timestamp 1644511149
transform 1 0 46460 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_501
timestamp 1644511149
transform 1 0 47196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_508
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_150
timestamp 1644511149
transform 1 0 14904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1644511149
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_186
timestamp 1644511149
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1644511149
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_217
timestamp 1644511149
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_224
timestamp 1644511149
transform 1 0 21712 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_274
timestamp 1644511149
transform 1 0 26312 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_286
timestamp 1644511149
transform 1 0 27416 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_298
timestamp 1644511149
transform 1 0 28520 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1644511149
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_330
timestamp 1644511149
transform 1 0 31464 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_342
timestamp 1644511149
transform 1 0 32568 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_354
timestamp 1644511149
transform 1 0 33672 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1644511149
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_498
timestamp 1644511149
transform 1 0 46920 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_510
timestamp 1644511149
transform 1 0 48024 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_154
timestamp 1644511149
transform 1 0 15272 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1644511149
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_202
timestamp 1644511149
transform 1 0 19688 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_214
timestamp 1644511149
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1644511149
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_230
timestamp 1644511149
transform 1 0 22264 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_239
timestamp 1644511149
transform 1 0 23092 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_251
timestamp 1644511149
transform 1 0 24196 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_263
timestamp 1644511149
transform 1 0 25300 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_275
timestamp 1644511149
transform 1 0 26404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_493
timestamp 1644511149
transform 1 0 46460 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1644511149
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_146
timestamp 1644511149
transform 1 0 14536 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1644511149
transform 1 0 15088 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_174
timestamp 1644511149
transform 1 0 17112 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1644511149
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1644511149
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_200
timestamp 1644511149
transform 1 0 19504 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_212
timestamp 1644511149
transform 1 0 20608 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1644511149
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_227
timestamp 1644511149
transform 1 0 21988 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_234
timestamp 1644511149
transform 1 0 22632 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1644511149
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1644511149
transform 1 0 25300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_275
timestamp 1644511149
transform 1 0 26404 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_287
timestamp 1644511149
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1644511149
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_480
timestamp 1644511149
transform 1 0 45264 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_492
timestamp 1644511149
transform 1 0 46368 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_507
timestamp 1644511149
transform 1 0 47748 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_515
timestamp 1644511149
transform 1 0 48484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 1644511149
transform 1 0 15180 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_157
timestamp 1644511149
transform 1 0 15548 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1644511149
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_187
timestamp 1644511149
transform 1 0 18308 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_194
timestamp 1644511149
transform 1 0 18952 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_202
timestamp 1644511149
transform 1 0 19688 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_206
timestamp 1644511149
transform 1 0 20056 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1644511149
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_245
timestamp 1644511149
transform 1 0 23644 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_259
timestamp 1644511149
transform 1 0 24932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_266
timestamp 1644511149
transform 1 0 25576 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1644511149
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_495
timestamp 1644511149
transform 1 0 46644 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_130
timestamp 1644511149
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1644511149
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1644511149
transform 1 0 14812 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_171
timestamp 1644511149
transform 1 0 16836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_179
timestamp 1644511149
transform 1 0 17572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1644511149
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_201
timestamp 1644511149
transform 1 0 19596 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_223
timestamp 1644511149
transform 1 0 21620 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_231
timestamp 1644511149
transform 1 0 22356 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_237
timestamp 1644511149
transform 1 0 22908 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_261
timestamp 1644511149
transform 1 0 25116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_268
timestamp 1644511149
transform 1 0 25760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1644511149
transform 1 0 26496 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_284
timestamp 1644511149
transform 1 0 27232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_291
timestamp 1644511149
transform 1 0 27876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1644511149
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_463
timestamp 1644511149
transform 1 0 43700 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_467
timestamp 1644511149
transform 1 0 44068 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_144
timestamp 1644511149
transform 1 0 14352 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_154
timestamp 1644511149
transform 1 0 15272 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_160
timestamp 1644511149
transform 1 0 15824 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_175
timestamp 1644511149
transform 1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_199
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_211
timestamp 1644511149
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_229
timestamp 1644511149
transform 1 0 22172 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_242
timestamp 1644511149
transform 1 0 23368 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_271
timestamp 1644511149
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_284
timestamp 1644511149
transform 1 0 27232 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_311
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_323
timestamp 1644511149
transform 1 0 30820 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1644511149
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_484
timestamp 1644511149
transform 1 0 45632 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_493
timestamp 1644511149
transform 1 0 46460 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_129
timestamp 1644511149
transform 1 0 12972 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_162
timestamp 1644511149
transform 1 0 16008 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_170
timestamp 1644511149
transform 1 0 16744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_178
timestamp 1644511149
transform 1 0 17480 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_219
timestamp 1644511149
transform 1 0 21252 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_231
timestamp 1644511149
transform 1 0 22356 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_235
timestamp 1644511149
transform 1 0 22724 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_243
timestamp 1644511149
transform 1 0 23460 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_266
timestamp 1644511149
transform 1 0 25576 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_272
timestamp 1644511149
transform 1 0 26128 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1644511149
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_282
timestamp 1644511149
transform 1 0 27048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_312
timestamp 1644511149
transform 1 0 29808 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_325
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_329
timestamp 1644511149
transform 1 0 31372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_347
timestamp 1644511149
transform 1 0 33028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_359
timestamp 1644511149
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_376
timestamp 1644511149
transform 1 0 35696 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_380
timestamp 1644511149
transform 1 0 36064 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_402
timestamp 1644511149
transform 1 0 38088 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_414
timestamp 1644511149
transform 1 0 39192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_485
timestamp 1644511149
transform 1 0 45724 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_129
timestamp 1644511149
transform 1 0 12972 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_150
timestamp 1644511149
transform 1 0 14904 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1644511149
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_176
timestamp 1644511149
transform 1 0 17296 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_185
timestamp 1644511149
transform 1 0 18124 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_197
timestamp 1644511149
transform 1 0 19228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_209
timestamp 1644511149
transform 1 0 20332 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_246
timestamp 1644511149
transform 1 0 23736 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_254
timestamp 1644511149
transform 1 0 24472 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_260
timestamp 1644511149
transform 1 0 25024 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1644511149
transform 1 0 27416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_294
timestamp 1644511149
transform 1 0 28152 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_303
timestamp 1644511149
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_315
timestamp 1644511149
transform 1 0 30084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_320
timestamp 1644511149
transform 1 0 30544 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_324
timestamp 1644511149
transform 1 0 30912 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_342
timestamp 1644511149
transform 1 0 32568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_414
timestamp 1644511149
transform 1 0 39192 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_426
timestamp 1644511149
transform 1 0 40296 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_438
timestamp 1644511149
transform 1 0 41400 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1644511149
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_455
timestamp 1644511149
transform 1 0 42964 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_475
timestamp 1644511149
transform 1 0 44804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_510
timestamp 1644511149
transform 1 0 48024 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_144
timestamp 1644511149
transform 1 0 14352 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_151
timestamp 1644511149
transform 1 0 14996 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_180
timestamp 1644511149
transform 1 0 17664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1644511149
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_232
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_240
timestamp 1644511149
transform 1 0 23184 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1644511149
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_283
timestamp 1644511149
transform 1 0 27140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_288
timestamp 1644511149
transform 1 0 27600 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_300
timestamp 1644511149
transform 1 0 28704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_331
timestamp 1644511149
transform 1 0 31556 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_340
timestamp 1644511149
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_347
timestamp 1644511149
transform 1 0 33028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_354
timestamp 1644511149
transform 1 0 33672 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1644511149
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_385
timestamp 1644511149
transform 1 0 36524 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_388
timestamp 1644511149
transform 1 0 36800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_396
timestamp 1644511149
transform 1 0 37536 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_408
timestamp 1644511149
transform 1 0 38640 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1644511149
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_481
timestamp 1644511149
transform 1 0 45356 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_119
timestamp 1644511149
transform 1 0 12052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_124
timestamp 1644511149
transform 1 0 12512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_134
timestamp 1644511149
transform 1 0 13432 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_144
timestamp 1644511149
transform 1 0 14352 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_148
timestamp 1644511149
transform 1 0 14720 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_153
timestamp 1644511149
transform 1 0 15180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1644511149
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_177
timestamp 1644511149
transform 1 0 17388 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1644511149
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_212
timestamp 1644511149
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1644511149
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_233
timestamp 1644511149
transform 1 0 22540 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_256
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_268
timestamp 1644511149
transform 1 0 25760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_297
timestamp 1644511149
transform 1 0 28428 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_304
timestamp 1644511149
transform 1 0 29072 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_316
timestamp 1644511149
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1644511149
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_346
timestamp 1644511149
transform 1 0 32936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_371
timestamp 1644511149
transform 1 0 35236 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_378
timestamp 1644511149
transform 1 0 35880 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1644511149
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_468
timestamp 1644511149
transform 1 0 44160 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_483
timestamp 1644511149
transform 1 0 45540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_499
timestamp 1644511149
transform 1 0 47012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_105
timestamp 1644511149
transform 1 0 10764 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_128
timestamp 1644511149
transform 1 0 12880 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1644511149
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_146
timestamp 1644511149
transform 1 0 14536 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_154
timestamp 1644511149
transform 1 0 15272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_178
timestamp 1644511149
transform 1 0 17480 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_186
timestamp 1644511149
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1644511149
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_222
timestamp 1644511149
transform 1 0 21528 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_234
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1644511149
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_257
timestamp 1644511149
transform 1 0 24748 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_286
timestamp 1644511149
transform 1 0 27416 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_298
timestamp 1644511149
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1644511149
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_330
timestamp 1644511149
transform 1 0 31464 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_340
timestamp 1644511149
transform 1 0 32384 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_347
timestamp 1644511149
transform 1 0 33028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 1644511149
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_368
timestamp 1644511149
transform 1 0 34960 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_372
timestamp 1644511149
transform 1 0 35328 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_394
timestamp 1644511149
transform 1 0 37352 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_406
timestamp 1644511149
transform 1 0 38456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1644511149
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_470
timestamp 1644511149
transform 1 0 44344 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_480
timestamp 1644511149
transform 1 0 45264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_487
timestamp 1644511149
transform 1 0 45908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_498
timestamp 1644511149
transform 1 0 46920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_502
timestamp 1644511149
transform 1 0 47288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_506
timestamp 1644511149
transform 1 0 47656 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_514
timestamp 1644511149
transform 1 0 48392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_99
timestamp 1644511149
transform 1 0 10212 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_104
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_117
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_133
timestamp 1644511149
transform 1 0 13340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1644511149
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_150
timestamp 1644511149
transform 1 0 14904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_154
timestamp 1644511149
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_176
timestamp 1644511149
transform 1 0 17296 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_184
timestamp 1644511149
transform 1 0 18032 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_206
timestamp 1644511149
transform 1 0 20056 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1644511149
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1644511149
transform 1 0 22448 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_244
timestamp 1644511149
transform 1 0 23552 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_256
timestamp 1644511149
transform 1 0 24656 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_263
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_274
timestamp 1644511149
transform 1 0 26312 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_285
timestamp 1644511149
transform 1 0 27324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_309
timestamp 1644511149
transform 1 0 29532 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_316
timestamp 1644511149
transform 1 0 30176 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_328
timestamp 1644511149
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_342
timestamp 1644511149
transform 1 0 32568 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_350
timestamp 1644511149
transform 1 0 33304 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_355
timestamp 1644511149
transform 1 0 33764 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1644511149
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_455
timestamp 1644511149
transform 1 0 42964 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_459
timestamp 1644511149
transform 1 0 43332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_469
timestamp 1644511149
transform 1 0 44252 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_477
timestamp 1644511149
transform 1 0 44988 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1644511149
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_512
timestamp 1644511149
transform 1 0 48208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_129
timestamp 1644511149
transform 1 0 12972 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_137
timestamp 1644511149
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_145
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_152
timestamp 1644511149
transform 1 0 15088 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_160
timestamp 1644511149
transform 1 0 15824 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_167
timestamp 1644511149
transform 1 0 16468 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_175
timestamp 1644511149
transform 1 0 17204 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1644511149
transform 1 0 17756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_188
timestamp 1644511149
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_205
timestamp 1644511149
transform 1 0 19964 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_213
timestamp 1644511149
transform 1 0 20700 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_242
timestamp 1644511149
transform 1 0 23368 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1644511149
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_258
timestamp 1644511149
transform 1 0 24840 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_262
timestamp 1644511149
transform 1 0 25208 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_284
timestamp 1644511149
transform 1 0 27232 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_292
timestamp 1644511149
transform 1 0 27968 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_298
timestamp 1644511149
transform 1 0 28520 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1644511149
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_316
timestamp 1644511149
transform 1 0 30176 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_337
timestamp 1644511149
transform 1 0 32108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_347
timestamp 1644511149
transform 1 0 33028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_354
timestamp 1644511149
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1644511149
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_369
timestamp 1644511149
transform 1 0 35052 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_383
timestamp 1644511149
transform 1 0 36340 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_390
timestamp 1644511149
transform 1 0 36984 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_402
timestamp 1644511149
transform 1 0 38088 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_414
timestamp 1644511149
transform 1 0 39192 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_466
timestamp 1644511149
transform 1 0 43976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1644511149
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_480
timestamp 1644511149
transform 1 0 45264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_487
timestamp 1644511149
transform 1 0 45908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_117
timestamp 1644511149
transform 1 0 11868 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_124
timestamp 1644511149
transform 1 0 12512 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_132
timestamp 1644511149
transform 1 0 13248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1644511149
transform 1 0 15456 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_175
timestamp 1644511149
transform 1 0 17204 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1644511149
transform 1 0 18308 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_229
timestamp 1644511149
transform 1 0 22172 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_236
timestamp 1644511149
transform 1 0 22816 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_242
timestamp 1644511149
transform 1 0 23368 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_248
timestamp 1644511149
transform 1 0 23920 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_255
timestamp 1644511149
transform 1 0 24564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_263
timestamp 1644511149
transform 1 0 25300 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_267
timestamp 1644511149
transform 1 0 25668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_284
timestamp 1644511149
transform 1 0 27232 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_297
timestamp 1644511149
transform 1 0 28428 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_304
timestamp 1644511149
transform 1 0 29072 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_346
timestamp 1644511149
transform 1 0 32936 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_359
timestamp 1644511149
transform 1 0 34132 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_376
timestamp 1644511149
transform 1 0 35696 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1644511149
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_408
timestamp 1644511149
transform 1 0 38640 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_420
timestamp 1644511149
transform 1 0 39744 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_432
timestamp 1644511149
transform 1 0 40848 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_440
timestamp 1644511149
transform 1 0 41584 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_444
timestamp 1644511149
transform 1 0 41952 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_458
timestamp 1644511149
transform 1 0 43240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_465
timestamp 1644511149
transform 1 0 43884 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_484
timestamp 1644511149
transform 1 0 45632 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_491
timestamp 1644511149
transform 1 0 46276 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1644511149
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1644511149
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_88
timestamp 1644511149
transform 1 0 9200 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_100
timestamp 1644511149
transform 1 0 10304 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_108
timestamp 1644511149
transform 1 0 11040 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_116
timestamp 1644511149
transform 1 0 11776 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1644511149
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_162
timestamp 1644511149
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_170
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_178
timestamp 1644511149
transform 1 0 17480 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_183
timestamp 1644511149
transform 1 0 17940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_204
timestamp 1644511149
transform 1 0 19872 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1644511149
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_219
timestamp 1644511149
transform 1 0 21252 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_227
timestamp 1644511149
transform 1 0 21988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_235
timestamp 1644511149
transform 1 0 22724 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 1644511149
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_258
timestamp 1644511149
transform 1 0 24840 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_264
timestamp 1644511149
transform 1 0 25392 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_268
timestamp 1644511149
transform 1 0 25760 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_280
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_286
timestamp 1644511149
transform 1 0 27416 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_298
timestamp 1644511149
transform 1 0 28520 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_303
timestamp 1644511149
transform 1 0 28980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_313
timestamp 1644511149
transform 1 0 29900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_320
timestamp 1644511149
transform 1 0 30544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_332
timestamp 1644511149
transform 1 0 31648 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_359
timestamp 1644511149
transform 1 0 34132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_371
timestamp 1644511149
transform 1 0 35236 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_375
timestamp 1644511149
transform 1 0 35604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_379
timestamp 1644511149
transform 1 0 35972 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_392
timestamp 1644511149
transform 1 0 37168 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1644511149
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_426
timestamp 1644511149
transform 1 0 40296 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_438
timestamp 1644511149
transform 1 0 41400 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_450
timestamp 1644511149
transform 1 0 42504 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_458
timestamp 1644511149
transform 1 0 43240 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_470
timestamp 1644511149
transform 1 0 44344 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_482
timestamp 1644511149
transform 1 0 45448 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_507
timestamp 1644511149
transform 1 0 47748 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_515
timestamp 1644511149
transform 1 0 48484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_77
timestamp 1644511149
transform 1 0 8188 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_101
timestamp 1644511149
transform 1 0 10396 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_109
timestamp 1644511149
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_136
timestamp 1644511149
transform 1 0 13616 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_177
timestamp 1644511149
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_200
timestamp 1644511149
transform 1 0 19504 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_212
timestamp 1644511149
transform 1 0 20608 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_232
timestamp 1644511149
transform 1 0 22448 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_241
timestamp 1644511149
transform 1 0 23276 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_248
timestamp 1644511149
transform 1 0 23920 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 1644511149
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_307
timestamp 1644511149
transform 1 0 29348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_319
timestamp 1644511149
transform 1 0 30452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1644511149
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_366
timestamp 1644511149
transform 1 0 34776 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_374
timestamp 1644511149
transform 1 0 35512 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_380
timestamp 1644511149
transform 1 0 36064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1644511149
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_415
timestamp 1644511149
transform 1 0 39284 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_419
timestamp 1644511149
transform 1 0 39652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_427
timestamp 1644511149
transform 1 0 40388 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_434
timestamp 1644511149
transform 1 0 41032 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_446
timestamp 1644511149
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_459
timestamp 1644511149
transform 1 0 43332 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_467
timestamp 1644511149
transform 1 0 44068 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_472
timestamp 1644511149
transform 1 0 44528 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_479
timestamp 1644511149
transform 1 0 45172 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_486
timestamp 1644511149
transform 1 0 45816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1644511149
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_88
timestamp 1644511149
transform 1 0 9200 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_100
timestamp 1644511149
transform 1 0 10304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_108
timestamp 1644511149
transform 1 0 11040 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_120
timestamp 1644511149
transform 1 0 12144 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1644511149
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_151
timestamp 1644511149
transform 1 0 14996 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_158
timestamp 1644511149
transform 1 0 15640 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_171
timestamp 1644511149
transform 1 0 16836 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_179
timestamp 1644511149
transform 1 0 17572 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_184
timestamp 1644511149
transform 1 0 18032 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_203
timestamp 1644511149
transform 1 0 19780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_208
timestamp 1644511149
transform 1 0 20240 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_216
timestamp 1644511149
transform 1 0 20976 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1644511149
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_261
timestamp 1644511149
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_283
timestamp 1644511149
transform 1 0 27140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_287
timestamp 1644511149
transform 1 0 27508 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_295
timestamp 1644511149
transform 1 0 28244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_385
timestamp 1644511149
transform 1 0 36524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_392
timestamp 1644511149
transform 1 0 37168 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_408
timestamp 1644511149
transform 1 0 38640 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_444
timestamp 1644511149
transform 1 0 41952 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_452
timestamp 1644511149
transform 1 0 42688 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_462
timestamp 1644511149
transform 1 0 43608 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_502
timestamp 1644511149
transform 1 0 47288 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_77
timestamp 1644511149
transform 1 0 8188 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_100
timestamp 1644511149
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_145
timestamp 1644511149
transform 1 0 14444 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_150
timestamp 1644511149
transform 1 0 14904 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_162
timestamp 1644511149
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_175
timestamp 1644511149
transform 1 0 17204 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_183
timestamp 1644511149
transform 1 0 17940 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_204
timestamp 1644511149
transform 1 0 19872 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_234
timestamp 1644511149
transform 1 0 22632 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_241
timestamp 1644511149
transform 1 0 23276 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_253
timestamp 1644511149
transform 1 0 24380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_266
timestamp 1644511149
transform 1 0 25576 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_308
timestamp 1644511149
transform 1 0 29440 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_320
timestamp 1644511149
transform 1 0 30544 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_403
timestamp 1644511149
transform 1 0 38180 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_411
timestamp 1644511149
transform 1 0 38916 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_419
timestamp 1644511149
transform 1 0 39652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_430
timestamp 1644511149
transform 1 0 40664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_434
timestamp 1644511149
transform 1 0 41032 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_439
timestamp 1644511149
transform 1 0 41492 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_455
timestamp 1644511149
transform 1 0 42964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_462
timestamp 1644511149
transform 1 0 43608 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_474
timestamp 1644511149
transform 1 0 44712 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_478
timestamp 1644511149
transform 1 0 45080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_120
timestamp 1644511149
transform 1 0 12144 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_127
timestamp 1644511149
transform 1 0 12788 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1644511149
transform 1 0 14352 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_156
timestamp 1644511149
transform 1 0 15456 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_175
timestamp 1644511149
transform 1 0 17204 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_185
timestamp 1644511149
transform 1 0 18124 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1644511149
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_203
timestamp 1644511149
transform 1 0 19780 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_207
timestamp 1644511149
transform 1 0 20148 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_229
timestamp 1644511149
transform 1 0 22172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_237
timestamp 1644511149
transform 1 0 22908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1644511149
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_256
timestamp 1644511149
transform 1 0 24656 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_268
timestamp 1644511149
transform 1 0 25760 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_280
timestamp 1644511149
transform 1 0 26864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_453
timestamp 1644511149
transform 1 0 42780 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_459
timestamp 1644511149
transform 1 0 43332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_471
timestamp 1644511149
transform 1 0 44436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_483
timestamp 1644511149
transform 1 0 45540 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_487
timestamp 1644511149
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_86
timestamp 1644511149
transform 1 0 9016 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_92
timestamp 1644511149
transform 1 0 9568 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_96
timestamp 1644511149
transform 1 0 9936 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_104
timestamp 1644511149
transform 1 0 10672 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_118
timestamp 1644511149
transform 1 0 11960 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_144
timestamp 1644511149
transform 1 0 14352 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_152
timestamp 1644511149
transform 1 0 15088 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_176
timestamp 1644511149
transform 1 0 17296 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_204
timestamp 1644511149
transform 1 0 19872 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_211
timestamp 1644511149
transform 1 0 20516 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_218
timestamp 1644511149
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_233
timestamp 1644511149
transform 1 0 22540 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_241
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_287
timestamp 1644511149
transform 1 0 27508 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_291
timestamp 1644511149
transform 1 0 27876 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_298
timestamp 1644511149
transform 1 0 28520 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_310
timestamp 1644511149
transform 1 0 29624 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_318
timestamp 1644511149
transform 1 0 30360 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_324
timestamp 1644511149
transform 1 0 30912 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_412
timestamp 1644511149
transform 1 0 39008 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_437
timestamp 1644511149
transform 1 0 41308 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_445
timestamp 1644511149
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_13
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1644511149
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_106
timestamp 1644511149
transform 1 0 10856 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_117
timestamp 1644511149
transform 1 0 11868 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1644511149
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1644511149
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_162
timestamp 1644511149
transform 1 0 16008 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_171
timestamp 1644511149
transform 1 0 16836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_182
timestamp 1644511149
transform 1 0 17848 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1644511149
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_239
timestamp 1644511149
transform 1 0 23092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_273
timestamp 1644511149
transform 1 0 26220 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_285
timestamp 1644511149
transform 1 0 27324 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_297
timestamp 1644511149
transform 1 0 28428 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1644511149
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_330
timestamp 1644511149
transform 1 0 31464 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_342
timestamp 1644511149
transform 1 0 32568 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_354
timestamp 1644511149
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1644511149
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_101
timestamp 1644511149
transform 1 0 10396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_107
timestamp 1644511149
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_117
timestamp 1644511149
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_121
timestamp 1644511149
transform 1 0 12236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_131
timestamp 1644511149
transform 1 0 13156 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_135
timestamp 1644511149
transform 1 0 13524 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_143
timestamp 1644511149
transform 1 0 14260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_154
timestamp 1644511149
transform 1 0 15272 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1644511149
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_174
timestamp 1644511149
transform 1 0 17112 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_184
timestamp 1644511149
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_191
timestamp 1644511149
transform 1 0 18676 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_203
timestamp 1644511149
transform 1 0 19780 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_215
timestamp 1644511149
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_245
timestamp 1644511149
transform 1 0 23644 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_252
timestamp 1644511149
transform 1 0 24288 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_256
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_260
timestamp 1644511149
transform 1 0 25024 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_267
timestamp 1644511149
transform 1 0 25668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_289
timestamp 1644511149
transform 1 0 27692 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_299
timestamp 1644511149
transform 1 0 28612 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_306
timestamp 1644511149
transform 1 0 29256 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_324
timestamp 1644511149
transform 1 0 30912 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_328
timestamp 1644511149
transform 1 0 31280 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_494
timestamp 1644511149
transform 1 0 46552 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_502
timestamp 1644511149
transform 1 0 47288 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_112
timestamp 1644511149
transform 1 0 11408 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_124
timestamp 1644511149
transform 1 0 12512 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1644511149
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_149
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_172
timestamp 1644511149
transform 1 0 16928 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_184
timestamp 1644511149
transform 1 0 18032 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_210
timestamp 1644511149
transform 1 0 20424 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_214
timestamp 1644511149
transform 1 0 20792 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_222
timestamp 1644511149
transform 1 0 21528 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_234
timestamp 1644511149
transform 1 0 22632 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1644511149
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_263
timestamp 1644511149
transform 1 0 25300 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_272
timestamp 1644511149
transform 1 0 26128 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_280
timestamp 1644511149
transform 1 0 26864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_303
timestamp 1644511149
transform 1 0 28980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_316
timestamp 1644511149
transform 1 0 30176 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_324
timestamp 1644511149
transform 1 0 30912 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_507
timestamp 1644511149
transform 1 0 47748 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_515
timestamp 1644511149
transform 1 0 48484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_134
timestamp 1644511149
transform 1 0 13432 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_142
timestamp 1644511149
transform 1 0 14168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_146
timestamp 1644511149
transform 1 0 14536 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_153
timestamp 1644511149
transform 1 0 15180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_160
timestamp 1644511149
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_197
timestamp 1644511149
transform 1 0 19228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_201
timestamp 1644511149
transform 1 0 19596 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1644511149
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_233
timestamp 1644511149
transform 1 0 22540 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_245
timestamp 1644511149
transform 1 0 23644 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_253
timestamp 1644511149
transform 1 0 24380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_264
timestamp 1644511149
transform 1 0 25392 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_275
timestamp 1644511149
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_291
timestamp 1644511149
transform 1 0 27876 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_301
timestamp 1644511149
transform 1 0 28796 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_307
timestamp 1644511149
transform 1 0 29348 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_314
timestamp 1644511149
transform 1 0 29992 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_325
timestamp 1644511149
transform 1 0 31004 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_344
timestamp 1644511149
transform 1 0 32752 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_356
timestamp 1644511149
transform 1 0 33856 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_368
timestamp 1644511149
transform 1 0 34960 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_380
timestamp 1644511149
transform 1 0 36064 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_164
timestamp 1644511149
transform 1 0 16192 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_200
timestamp 1644511149
transform 1 0 19504 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_206
timestamp 1644511149
transform 1 0 20056 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_212
timestamp 1644511149
transform 1 0 20608 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_223
timestamp 1644511149
transform 1 0 21620 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_238
timestamp 1644511149
transform 1 0 23000 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_247
timestamp 1644511149
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_274
timestamp 1644511149
transform 1 0 26312 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_286
timestamp 1644511149
transform 1 0 27416 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_299
timestamp 1644511149
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_317
timestamp 1644511149
transform 1 0 30268 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_327
timestamp 1644511149
transform 1 0 31188 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_337
timestamp 1644511149
transform 1 0 32108 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_349
timestamp 1644511149
transform 1 0 33212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1644511149
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_191
timestamp 1644511149
transform 1 0 18676 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_199
timestamp 1644511149
transform 1 0 19412 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_208
timestamp 1644511149
transform 1 0 20240 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_230
timestamp 1644511149
transform 1 0 22264 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_240
timestamp 1644511149
transform 1 0 23184 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_255
timestamp 1644511149
transform 1 0 24564 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_269
timestamp 1644511149
transform 1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1644511149
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_310
timestamp 1644511149
transform 1 0 29624 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_318
timestamp 1644511149
transform 1 0 30360 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1644511149
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_500
timestamp 1644511149
transform 1 0 47104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_183
timestamp 1644511149
transform 1 0 17940 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_208
timestamp 1644511149
transform 1 0 20240 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_216
timestamp 1644511149
transform 1 0 20976 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_228
timestamp 1644511149
transform 1 0 22080 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_232
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_242
timestamp 1644511149
transform 1 0 23368 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1644511149
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_284
timestamp 1644511149
transform 1 0 27232 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_292
timestamp 1644511149
transform 1 0 27968 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_298
timestamp 1644511149
transform 1 0 28520 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1644511149
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_319
timestamp 1644511149
transform 1 0 30452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_331
timestamp 1644511149
transform 1 0 31556 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_343
timestamp 1644511149
transform 1 0 32660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_355
timestamp 1644511149
transform 1 0 33764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_189
timestamp 1644511149
transform 1 0 18492 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_196
timestamp 1644511149
transform 1 0 19136 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_206
timestamp 1644511149
transform 1 0 20056 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_210
timestamp 1644511149
transform 1 0 20424 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1644511149
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_233
timestamp 1644511149
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_254
timestamp 1644511149
transform 1 0 24472 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_265
timestamp 1644511149
transform 1 0 25484 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_285
timestamp 1644511149
transform 1 0 27324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_304
timestamp 1644511149
transform 1 0 29072 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_323
timestamp 1644511149
transform 1 0 30820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_340
timestamp 1644511149
transform 1 0 32384 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_352
timestamp 1644511149
transform 1 0 33488 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_364
timestamp 1644511149
transform 1 0 34592 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_376
timestamp 1644511149
transform 1 0 35696 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1644511149
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_186
timestamp 1644511149
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1644511149
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_204
timestamp 1644511149
transform 1 0 19872 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_217
timestamp 1644511149
transform 1 0 21068 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_229
timestamp 1644511149
transform 1 0 22172 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_241
timestamp 1644511149
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1644511149
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_264
timestamp 1644511149
transform 1 0 25392 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_272
timestamp 1644511149
transform 1 0 26128 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_280
timestamp 1644511149
transform 1 0 26864 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_302
timestamp 1644511149
transform 1 0 28888 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_315
timestamp 1644511149
transform 1 0 30084 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_339
timestamp 1644511149
transform 1 0 32292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_351
timestamp 1644511149
transform 1 0 33396 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_192
timestamp 1644511149
transform 1 0 18768 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_196
timestamp 1644511149
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_206
timestamp 1644511149
transform 1 0 20056 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_218
timestamp 1644511149
transform 1 0 21160 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_254
timestamp 1644511149
transform 1 0 24472 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_262
timestamp 1644511149
transform 1 0 25208 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_272
timestamp 1644511149
transform 1 0 26128 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_285
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_290
timestamp 1644511149
transform 1 0 27784 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_301
timestamp 1644511149
transform 1 0 28796 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_307
timestamp 1644511149
transform 1 0 29348 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_312
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_321
timestamp 1644511149
transform 1 0 30636 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_365
timestamp 1644511149
transform 1 0 34684 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_377
timestamp 1644511149
transform 1 0 35788 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_389
timestamp 1644511149
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1644511149
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_217
timestamp 1644511149
transform 1 0 21068 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_227
timestamp 1644511149
transform 1 0 21988 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_234
timestamp 1644511149
transform 1 0 22632 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1644511149
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_257
timestamp 1644511149
transform 1 0 24748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_266
timestamp 1644511149
transform 1 0 25576 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_274
timestamp 1644511149
transform 1 0 26312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_282
timestamp 1644511149
transform 1 0 27048 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_290
timestamp 1644511149
transform 1 0 27784 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_296
timestamp 1644511149
transform 1 0 28336 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1644511149
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_317
timestamp 1644511149
transform 1 0 30268 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_325
timestamp 1644511149
transform 1 0 31004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_337
timestamp 1644511149
transform 1 0 32108 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_349
timestamp 1644511149
transform 1 0 33212 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1644511149
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_495
timestamp 1644511149
transform 1 0 46644 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_509
timestamp 1644511149
transform 1 0 47932 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_515
timestamp 1644511149
transform 1 0 48484 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_37
timestamp 1644511149
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_49
timestamp 1644511149
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_64
timestamp 1644511149
transform 1 0 6992 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_76
timestamp 1644511149
transform 1 0 8096 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_88
timestamp 1644511149
transform 1 0 9200 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_100
timestamp 1644511149
transform 1 0 10304 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1644511149
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_177
timestamp 1644511149
transform 1 0 17388 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_184
timestamp 1644511149
transform 1 0 18032 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_192
timestamp 1644511149
transform 1 0 18768 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_203
timestamp 1644511149
transform 1 0 19780 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_211
timestamp 1644511149
transform 1 0 20516 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_245
timestamp 1644511149
transform 1 0 23644 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_253
timestamp 1644511149
transform 1 0 24380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_269
timestamp 1644511149
transform 1 0 25852 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_277
timestamp 1644511149
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_285
timestamp 1644511149
transform 1 0 27324 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_294
timestamp 1644511149
transform 1 0 28152 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_300
timestamp 1644511149
transform 1 0 28704 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_304
timestamp 1644511149
transform 1 0 29072 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_316
timestamp 1644511149
transform 1 0 30176 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_353
timestamp 1644511149
transform 1 0 33580 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_357
timestamp 1644511149
transform 1 0 33948 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_369
timestamp 1644511149
transform 1 0 35052 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_381
timestamp 1644511149
transform 1 0 36156 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1644511149
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_32
timestamp 1644511149
transform 1 0 4048 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_44
timestamp 1644511149
transform 1 0 5152 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_56
timestamp 1644511149
transform 1 0 6256 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_68
timestamp 1644511149
transform 1 0 7360 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_72
timestamp 1644511149
transform 1 0 7728 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_159
timestamp 1644511149
transform 1 0 15732 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_180
timestamp 1644511149
transform 1 0 17664 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_219
timestamp 1644511149
transform 1 0 21252 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_241
timestamp 1644511149
transform 1 0 23276 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1644511149
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_279
timestamp 1644511149
transform 1 0 26772 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1644511149
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_312
timestamp 1644511149
transform 1 0 29808 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_324
timestamp 1644511149
transform 1 0 30912 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_334
timestamp 1644511149
transform 1 0 31832 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1644511149
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_507
timestamp 1644511149
transform 1 0 47748 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_515
timestamp 1644511149
transform 1 0 48484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_32
timestamp 1644511149
transform 1 0 4048 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_44
timestamp 1644511149
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_176
timestamp 1644511149
transform 1 0 17296 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_180
timestamp 1644511149
transform 1 0 17664 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_191
timestamp 1644511149
transform 1 0 18676 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_202
timestamp 1644511149
transform 1 0 19688 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_232
timestamp 1644511149
transform 1 0 22448 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_240
timestamp 1644511149
transform 1 0 23184 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_264
timestamp 1644511149
transform 1 0 25392 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_289
timestamp 1644511149
transform 1 0 27692 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_297
timestamp 1644511149
transform 1 0 28428 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_304
timestamp 1644511149
transform 1 0 29072 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_312
timestamp 1644511149
transform 1 0 29808 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_322
timestamp 1644511149
transform 1 0 30728 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_342
timestamp 1644511149
transform 1 0 32568 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_356
timestamp 1644511149
transform 1 0 33856 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_368
timestamp 1644511149
transform 1 0 34960 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_380
timestamp 1644511149
transform 1 0 36064 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_512
timestamp 1644511149
transform 1 0 48208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_14
timestamp 1644511149
transform 1 0 2392 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1644511149
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_173
timestamp 1644511149
transform 1 0 17020 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_181
timestamp 1644511149
transform 1 0 17756 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_203
timestamp 1644511149
transform 1 0 19780 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_215
timestamp 1644511149
transform 1 0 20884 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_224
timestamp 1644511149
transform 1 0 21712 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_231
timestamp 1644511149
transform 1 0 22356 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_243
timestamp 1644511149
transform 1 0 23460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_257
timestamp 1644511149
transform 1 0 24748 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_268
timestamp 1644511149
transform 1 0 25760 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_275
timestamp 1644511149
transform 1 0 26404 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_283
timestamp 1644511149
transform 1 0 27140 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_292
timestamp 1644511149
transform 1 0 27968 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_296
timestamp 1644511149
transform 1 0 28336 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_312
timestamp 1644511149
transform 1 0 29808 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_324
timestamp 1644511149
transform 1 0 30912 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_346
timestamp 1644511149
transform 1 0 32936 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_358
timestamp 1644511149
transform 1 0 34040 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_173
timestamp 1644511149
transform 1 0 17020 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_180
timestamp 1644511149
transform 1 0 17664 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_192
timestamp 1644511149
transform 1 0 18768 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_207
timestamp 1644511149
transform 1 0 20148 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_219
timestamp 1644511149
transform 1 0 21252 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_230
timestamp 1644511149
transform 1 0 22264 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_238
timestamp 1644511149
transform 1 0 23000 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_250
timestamp 1644511149
transform 1 0 24104 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_255
timestamp 1644511149
transform 1 0 24564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_262
timestamp 1644511149
transform 1 0 25208 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_274
timestamp 1644511149
transform 1 0 26312 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_302
timestamp 1644511149
transform 1 0 28888 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_314
timestamp 1644511149
transform 1 0 29992 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_493
timestamp 1644511149
transform 1 0 46460 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_511
timestamp 1644511149
transform 1 0 48116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_515
timestamp 1644511149
transform 1 0 48484 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_179
timestamp 1644511149
transform 1 0 17572 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_191
timestamp 1644511149
transform 1 0 18676 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_206
timestamp 1644511149
transform 1 0 20056 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_214
timestamp 1644511149
transform 1 0 20792 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_224
timestamp 1644511149
transform 1 0 21712 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_234
timestamp 1644511149
transform 1 0 22632 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_242
timestamp 1644511149
transform 1 0 23368 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1644511149
transform 1 0 23828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_264
timestamp 1644511149
transform 1 0 25392 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_272
timestamp 1644511149
transform 1 0 26128 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1644511149
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_317
timestamp 1644511149
transform 1 0 30268 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_326
timestamp 1644511149
transform 1 0 31096 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_338
timestamp 1644511149
transform 1 0 32200 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_350
timestamp 1644511149
transform 1 0 33304 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1644511149
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_497
timestamp 1644511149
transform 1 0 46828 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_182
timestamp 1644511149
transform 1 0 17848 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_208
timestamp 1644511149
transform 1 0 20240 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_212
timestamp 1644511149
transform 1 0 20608 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_219
timestamp 1644511149
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_233
timestamp 1644511149
transform 1 0 22540 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_242
timestamp 1644511149
transform 1 0 23368 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_248
timestamp 1644511149
transform 1 0 23920 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_255
timestamp 1644511149
transform 1 0 24564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_259
timestamp 1644511149
transform 1 0 24932 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_268
timestamp 1644511149
transform 1 0 25760 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_296
timestamp 1644511149
transform 1 0 28336 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_303
timestamp 1644511149
transform 1 0 28980 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_314
timestamp 1644511149
transform 1 0 29992 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_326
timestamp 1644511149
transform 1 0 31096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1644511149
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_508
timestamp 1644511149
transform 1 0 47840 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_175
timestamp 1644511149
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_187
timestamp 1644511149
transform 1 0 18308 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_201
timestamp 1644511149
transform 1 0 19596 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1644511149
transform 1 0 20884 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_219
timestamp 1644511149
transform 1 0 21252 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_227
timestamp 1644511149
transform 1 0 21988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_239
timestamp 1644511149
transform 1 0 23092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_258
timestamp 1644511149
transform 1 0 24840 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_270
timestamp 1644511149
transform 1 0 25944 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_281
timestamp 1644511149
transform 1 0 26956 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_293
timestamp 1644511149
transform 1 0 28060 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_297
timestamp 1644511149
transform 1 0 28428 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_315
timestamp 1644511149
transform 1 0 30084 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_326
timestamp 1644511149
transform 1 0 31096 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_338
timestamp 1644511149
transform 1 0 32200 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_350
timestamp 1644511149
transform 1 0 33304 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1644511149
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_177
timestamp 1644511149
transform 1 0 17388 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_235
timestamp 1644511149
transform 1 0 22724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_247
timestamp 1644511149
transform 1 0 23828 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_257
timestamp 1644511149
transform 1 0 24748 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_265
timestamp 1644511149
transform 1 0 25484 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_289
timestamp 1644511149
transform 1 0 27692 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_298
timestamp 1644511149
transform 1 0 28520 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_311
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_332
timestamp 1644511149
transform 1 0 31648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_512
timestamp 1644511149
transform 1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1644511149
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_173
timestamp 1644511149
transform 1 0 17020 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_182
timestamp 1644511149
transform 1 0 17848 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_219
timestamp 1644511149
transform 1 0 21252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_226
timestamp 1644511149
transform 1 0 21896 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_230
timestamp 1644511149
transform 1 0 22264 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_235
timestamp 1644511149
transform 1 0 22724 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_243
timestamp 1644511149
transform 1 0 23460 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1644511149
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_261
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_268
timestamp 1644511149
transform 1 0 25760 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_276
timestamp 1644511149
transform 1 0 26496 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_288
timestamp 1644511149
transform 1 0 27600 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1644511149
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_314
timestamp 1644511149
transform 1 0 29992 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_326
timestamp 1644511149
transform 1 0 31096 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_338
timestamp 1644511149
transform 1 0 32200 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_350
timestamp 1644511149
transform 1 0 33304 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1644511149
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_28
timestamp 1644511149
transform 1 0 3680 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1644511149
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_190
timestamp 1644511149
transform 1 0 18584 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_198
timestamp 1644511149
transform 1 0 19320 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1644511149
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_265
timestamp 1644511149
transform 1 0 25484 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_269
timestamp 1644511149
transform 1 0 25852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_314
timestamp 1644511149
transform 1 0 29992 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_320
timestamp 1644511149
transform 1 0 30544 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_324
timestamp 1644511149
transform 1 0 30912 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1644511149
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_224
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_236
timestamp 1644511149
transform 1 0 22816 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_243
timestamp 1644511149
transform 1 0 23460 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_259
timestamp 1644511149
transform 1 0 24932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_267
timestamp 1644511149
transform 1 0 25668 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_290
timestamp 1644511149
transform 1 0 27784 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_314
timestamp 1644511149
transform 1 0 29992 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_326
timestamp 1644511149
transform 1 0 31096 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_338
timestamp 1644511149
transform 1 0 32200 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_350
timestamp 1644511149
transform 1 0 33304 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1644511149
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_187
timestamp 1644511149
transform 1 0 18308 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_199
timestamp 1644511149
transform 1 0 19412 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_231
timestamp 1644511149
transform 1 0 22356 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_252
timestamp 1644511149
transform 1 0 24288 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1644511149
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_284
timestamp 1644511149
transform 1 0 27232 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_291
timestamp 1644511149
transform 1 0 27876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_303
timestamp 1644511149
transform 1 0 28980 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_310
timestamp 1644511149
transform 1 0 29624 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_322
timestamp 1644511149
transform 1 0 30728 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 1644511149
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_412
timestamp 1644511149
transform 1 0 39008 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_427
timestamp 1644511149
transform 1 0 40388 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_439
timestamp 1644511149
transform 1 0 41492 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_493
timestamp 1644511149
transform 1 0 46460 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_499
timestamp 1644511149
transform 1 0 47012 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_200
timestamp 1644511149
transform 1 0 19504 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_212
timestamp 1644511149
transform 1 0 20608 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_216
timestamp 1644511149
transform 1 0 20976 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_220
timestamp 1644511149
transform 1 0 21344 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_224
timestamp 1644511149
transform 1 0 21712 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_236
timestamp 1644511149
transform 1 0 22816 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_240
timestamp 1644511149
transform 1 0 23184 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_256
timestamp 1644511149
transform 1 0 24656 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_268
timestamp 1644511149
transform 1 0 25760 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_280
timestamp 1644511149
transform 1 0 26864 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_292
timestamp 1644511149
transform 1 0 27968 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1644511149
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_416
timestamp 1644511149
transform 1 0 39376 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_201
timestamp 1644511149
transform 1 0 19596 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_208
timestamp 1644511149
transform 1 0 20240 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_220
timestamp 1644511149
transform 1 0 21344 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_245
timestamp 1644511149
transform 1 0 23644 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_256
timestamp 1644511149
transform 1 0 24656 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_268
timestamp 1644511149
transform 1 0 25760 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_412
timestamp 1644511149
transform 1 0 39008 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_425
timestamp 1644511149
transform 1 0 40204 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_437
timestamp 1644511149
transform 1 0 41308 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_445
timestamp 1644511149
transform 1 0 42044 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_237
timestamp 1644511149
transform 1 0 22908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_249
timestamp 1644511149
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_262
timestamp 1644511149
transform 1 0 25208 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_266
timestamp 1644511149
transform 1 0 25576 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_278
timestamp 1644511149
transform 1 0 26680 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_290
timestamp 1644511149
transform 1 0 27784 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_302
timestamp 1644511149
transform 1 0 28888 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_493
timestamp 1644511149
transform 1 0 46460 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_499
timestamp 1644511149
transform 1 0 47012 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1644511149
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_9
timestamp 1644511149
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_13
timestamp 1644511149
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_25
timestamp 1644511149
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_37
timestamp 1644511149
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1644511149
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1644511149
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1644511149
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1644511149
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_9
timestamp 1644511149
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_21
timestamp 1644511149
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_284
timestamp 1644511149
transform 1 0 27232 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_296
timestamp 1644511149
transform 1 0 28336 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_412
timestamp 1644511149
transform 1 0 39008 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_479
timestamp 1644511149
transform 1 0 45172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_486
timestamp 1644511149
transform 1 0 45816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_11
timestamp 1644511149
transform 1 0 2116 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_261
timestamp 1644511149
transform 1 0 25116 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_266
timestamp 1644511149
transform 1 0 25576 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_278
timestamp 1644511149
transform 1 0 26680 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_290
timestamp 1644511149
transform 1 0 27784 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_302
timestamp 1644511149
transform 1 0 28888 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_460
timestamp 1644511149
transform 1 0 43424 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_464
timestamp 1644511149
transform 1 0 43792 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_468
timestamp 1644511149
transform 1 0 44160 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_28
timestamp 1644511149
transform 1 0 3680 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_40
timestamp 1644511149
transform 1 0 4784 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1644511149
transform 1 0 5888 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_119
timestamp 1644511149
transform 1 0 12052 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_131
timestamp 1644511149
transform 1 0 13156 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_143
timestamp 1644511149
transform 1 0 14260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_155
timestamp 1644511149
transform 1 0 15364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_213
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_218
timestamp 1644511149
transform 1 0 21160 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_266
timestamp 1644511149
transform 1 0 25576 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1644511149
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_345
timestamp 1644511149
transform 1 0 32844 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_425
timestamp 1644511149
transform 1 0 40204 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_440
timestamp 1644511149
transform 1 0 41584 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_473
timestamp 1644511149
transform 1 0 44620 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_498
timestamp 1644511149
transform 1 0 46920 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_79_505
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_512
timestamp 1644511149
transform 1 0 48208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_7
timestamp 1644511149
transform 1 0 1748 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_11
timestamp 1644511149
transform 1 0 2116 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_23
timestamp 1644511149
transform 1 0 3220 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_38
timestamp 1644511149
transform 1 0 4600 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_42
timestamp 1644511149
transform 1 0 4968 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_46
timestamp 1644511149
transform 1 0 5336 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_58
timestamp 1644511149
transform 1 0 6440 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_70
timestamp 1644511149
transform 1 0 7544 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1644511149
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_125
timestamp 1644511149
transform 1 0 12604 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1644511149
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_206
timestamp 1644511149
transform 1 0 20056 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_235
timestamp 1644511149
transform 1 0 22724 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_247
timestamp 1644511149
transform 1 0 23828 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_258
timestamp 1644511149
transform 1 0 24840 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_283
timestamp 1644511149
transform 1 0 27140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_295
timestamp 1644511149
transform 1 0 28244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_342
timestamp 1644511149
transform 1 0 32568 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_354
timestamp 1644511149
transform 1 0 33672 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_362
timestamp 1644511149
transform 1 0 34408 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_406
timestamp 1644511149
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1644511149
transform 1 0 39560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_455
timestamp 1644511149
transform 1 0 42964 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_462
timestamp 1644511149
transform 1 0 43608 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_468
timestamp 1644511149
transform 1 0 44160 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_472
timestamp 1644511149
transform 1 0 44528 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_13
timestamp 1644511149
transform 1 0 2300 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_25
timestamp 1644511149
transform 1 0 3404 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1644511149
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1644511149
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_134
timestamp 1644511149
transform 1 0 13432 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_159
timestamp 1644511149
transform 1 0 15732 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_359
timestamp 1644511149
transform 1 0 34132 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_371
timestamp 1644511149
transform 1 0 35236 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_383
timestamp 1644511149
transform 1 0 36340 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_438
timestamp 1644511149
transform 1 0 41400 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_446
timestamp 1644511149
transform 1 0 42136 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1644511149
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_63
timestamp 1644511149
transform 1 0 6900 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_71
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_121
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_132
timestamp 1644511149
transform 1 0 13248 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_145
timestamp 1644511149
transform 1 0 14444 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_191
timestamp 1644511149
transform 1 0 18676 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_207
timestamp 1644511149
transform 1 0 20148 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_213
timestamp 1644511149
transform 1 0 20700 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_217
timestamp 1644511149
transform 1 0 21068 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_223
timestamp 1644511149
transform 1 0 21620 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_228
timestamp 1644511149
transform 1 0 22080 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_235
timestamp 1644511149
transform 1 0 22724 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_247
timestamp 1644511149
transform 1 0 23828 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1644511149
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_259
timestamp 1644511149
transform 1 0 24932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_271
timestamp 1644511149
transform 1 0 26036 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_279
timestamp 1644511149
transform 1 0 26772 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1644511149
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_332
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_406
timestamp 1644511149
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_418
timestamp 1644511149
transform 1 0 39560 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_440
timestamp 1644511149
transform 1 0 41584 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_453
timestamp 1644511149
transform 1 0 42780 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_461
timestamp 1644511149
transform 1 0 43516 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1644511149
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1644511149
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_511
timestamp 1644511149
transform 1 0 48116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_515
timestamp 1644511149
transform 1 0 48484 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24472 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0598_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29808 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0599_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0601_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0602_
timestamp 1644511149
transform 1 0 20792 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0603_
timestamp 1644511149
transform 1 0 21160 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0604_
timestamp 1644511149
transform 1 0 28520 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0605_
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0606_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0607_
timestamp 1644511149
transform 1 0 22080 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19780 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0609_
timestamp 1644511149
transform 1 0 23552 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0610_
timestamp 1644511149
transform 1 0 25668 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0611_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20976 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24472 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0613_
timestamp 1644511149
transform 1 0 24840 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1644511149
transform 1 0 26956 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23092 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0616_
timestamp 1644511149
transform 1 0 21160 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0618_
timestamp 1644511149
transform 1 0 16836 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0619_
timestamp 1644511149
transform 1 0 16008 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0620_
timestamp 1644511149
transform 1 0 22448 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0621_
timestamp 1644511149
transform 1 0 22080 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0622_
timestamp 1644511149
transform 1 0 22724 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0623_
timestamp 1644511149
transform 1 0 12420 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0624_
timestamp 1644511149
transform 1 0 16560 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0625_
timestamp 1644511149
transform 1 0 17204 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _0626_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20056 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0627_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0628_
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0629_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27600 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0631_
timestamp 1644511149
transform 1 0 28060 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0632_
timestamp 1644511149
transform 1 0 25668 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1644511149
transform 1 0 29900 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0634_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28796 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1644511149
transform 1 0 30268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0637_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0639_
timestamp 1644511149
transform 1 0 22816 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0640_
timestamp 1644511149
transform 1 0 22356 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0641_
timestamp 1644511149
transform 1 0 24288 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0642_
timestamp 1644511149
transform 1 0 20608 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1644511149
transform 1 0 22540 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0644_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1644511149
transform 1 0 23000 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0646_
timestamp 1644511149
transform 1 0 22080 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0647_
timestamp 1644511149
transform 1 0 23644 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1644511149
transform 1 0 20976 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0649_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1644511149
transform 1 0 20240 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0651_
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0652_
timestamp 1644511149
transform 1 0 16376 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0653_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0654_
timestamp 1644511149
transform 1 0 15824 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0655_
timestamp 1644511149
transform 1 0 18216 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0656_
timestamp 1644511149
transform 1 0 18400 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1644511149
transform 1 0 19504 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0658_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0661_
timestamp 1644511149
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1644511149
transform 1 0 15364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0663_
timestamp 1644511149
transform 1 0 16192 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1644511149
transform 1 0 14996 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0665_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0666_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13616 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0668_
timestamp 1644511149
transform 1 0 11224 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0669_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1644511149
transform 1 0 12512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0671_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0672_
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1644511149
transform 1 0 11960 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0674_
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0675_
timestamp 1644511149
transform 1 0 10396 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0676_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1644511149
transform 1 0 11960 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0678_
timestamp 1644511149
transform 1 0 10396 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1644511149
transform 1 0 12236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0680_
timestamp 1644511149
transform 1 0 16836 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0681_
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0682_
timestamp 1644511149
transform 1 0 12604 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1644511149
transform 1 0 13248 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0685_
timestamp 1644511149
transform 1 0 14076 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0686_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0688_
timestamp 1644511149
transform 1 0 13800 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0689_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0690_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14720 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0692_
timestamp 1644511149
transform 1 0 12420 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0693_
timestamp 1644511149
transform 1 0 17848 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0695_
timestamp 1644511149
transform 1 0 17940 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0696_
timestamp 1644511149
transform 1 0 17848 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0697_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1644511149
transform 1 0 19688 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0699_
timestamp 1644511149
transform 1 0 16744 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0700_
timestamp 1644511149
transform 1 0 18032 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1644511149
transform 1 0 18676 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0702_
timestamp 1644511149
transform 1 0 17940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0703_
timestamp 1644511149
transform 1 0 17848 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1644511149
transform 1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0705_
timestamp 1644511149
transform 1 0 17572 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1644511149
transform 1 0 24748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0708_
timestamp 1644511149
transform 1 0 23276 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0709_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0710_
timestamp 1644511149
transform 1 0 18952 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0711_
timestamp 1644511149
transform 1 0 22172 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0712_
timestamp 1644511149
transform 1 0 22816 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1644511149
transform 1 0 22816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0714_
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0715_
timestamp 1644511149
transform 1 0 21344 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1644511149
transform 1 0 24932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0717_
timestamp 1644511149
transform 1 0 23276 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1644511149
transform 1 0 22356 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0719_
timestamp 1644511149
transform 1 0 24472 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0720_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0721_
timestamp 1644511149
transform 1 0 20976 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1644511149
transform 1 0 22448 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0723_
timestamp 1644511149
transform 1 0 20608 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0725_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24932 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0726_
timestamp 1644511149
transform 1 0 24380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0727_
timestamp 1644511149
transform 1 0 25300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0728_
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0730_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0731_
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1644511149
transform 1 0 28704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0733_
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0734_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0735_
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0736_
timestamp 1644511149
transform 1 0 28244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0737_
timestamp 1644511149
transform 1 0 29256 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0738_
timestamp 1644511149
transform 1 0 26864 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1644511149
transform 1 0 26128 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0740_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20608 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0741_
timestamp 1644511149
transform 1 0 23368 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0742_
timestamp 1644511149
transform 1 0 24656 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1644511149
transform 1 0 28704 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0744_
timestamp 1644511149
transform 1 0 25944 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0745_
timestamp 1644511149
transform 1 0 25852 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0746_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24656 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0747_
timestamp 1644511149
transform 1 0 27324 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0748_
timestamp 1644511149
transform 1 0 22724 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0749_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24656 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0750_
timestamp 1644511149
transform 1 0 25484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0751_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0752_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0753_
timestamp 1644511149
transform 1 0 25760 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0754_
timestamp 1644511149
transform 1 0 25576 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0755_
timestamp 1644511149
transform 1 0 27324 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0756_
timestamp 1644511149
transform 1 0 22356 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0757_
timestamp 1644511149
transform 1 0 22632 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0758_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24840 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0759_
timestamp 1644511149
transform 1 0 25852 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0760_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0761_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _0762_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0763_
timestamp 1644511149
transform 1 0 27508 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0764_
timestamp 1644511149
transform 1 0 25116 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0765_
timestamp 1644511149
transform 1 0 25484 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0766_
timestamp 1644511149
transform 1 0 20884 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0767_
timestamp 1644511149
transform 1 0 20148 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0768_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0769_
timestamp 1644511149
transform 1 0 25116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0770_
timestamp 1644511149
transform 1 0 18308 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0771_
timestamp 1644511149
transform 1 0 19504 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0772_
timestamp 1644511149
transform 1 0 20424 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0773_
timestamp 1644511149
transform 1 0 20516 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0774_
timestamp 1644511149
transform 1 0 26680 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0775_
timestamp 1644511149
transform 1 0 24104 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0776_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0777_
timestamp 1644511149
transform 1 0 19780 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0778_
timestamp 1644511149
transform 1 0 19228 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0779_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0780_
timestamp 1644511149
transform 1 0 19320 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0781_
timestamp 1644511149
transform 1 0 19964 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0782_
timestamp 1644511149
transform 1 0 19504 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0783_
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0784_
timestamp 1644511149
transform 1 0 23460 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0785_
timestamp 1644511149
transform 1 0 21988 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0786_
timestamp 1644511149
transform 1 0 21068 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0787_
timestamp 1644511149
transform 1 0 20884 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0788_
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_2  _0789_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0790_
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0791_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0792_
timestamp 1644511149
transform 1 0 22632 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0793_
timestamp 1644511149
transform 1 0 26128 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0794_
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0795_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23552 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0796_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0797_
timestamp 1644511149
transform 1 0 23000 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1644511149
transform 1 0 25576 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0799_
timestamp 1644511149
transform 1 0 28704 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0800_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0801_
timestamp 1644511149
transform 1 0 24932 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26312 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0803_
timestamp 1644511149
transform 1 0 25668 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0804_
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0805_
timestamp 1644511149
transform 1 0 29440 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0806_
timestamp 1644511149
transform 1 0 26128 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0807_
timestamp 1644511149
transform 1 0 25760 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0808_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25024 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0809_
timestamp 1644511149
transform 1 0 25208 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0810_
timestamp 1644511149
transform 1 0 20516 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0811_
timestamp 1644511149
transform 1 0 28428 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0812_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0813_
timestamp 1644511149
transform 1 0 29348 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0814_
timestamp 1644511149
transform 1 0 30268 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0815_
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0816_
timestamp 1644511149
transform 1 0 28336 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0817_
timestamp 1644511149
transform 1 0 28152 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0818_
timestamp 1644511149
transform 1 0 28152 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0819_
timestamp 1644511149
transform 1 0 28888 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0820_
timestamp 1644511149
transform 1 0 27692 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0821_
timestamp 1644511149
transform 1 0 27508 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0822_
timestamp 1644511149
transform 1 0 27324 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0823_
timestamp 1644511149
transform 1 0 28796 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0824_
timestamp 1644511149
transform 1 0 27416 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0825_
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0826_
timestamp 1644511149
transform 1 0 18308 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0827_
timestamp 1644511149
transform 1 0 30728 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0828_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29900 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0829_
timestamp 1644511149
transform 1 0 18216 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0830_
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0831_
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0832_
timestamp 1644511149
transform 1 0 24472 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0833_
timestamp 1644511149
transform 1 0 24932 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0834_
timestamp 1644511149
transform 1 0 24288 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0835_
timestamp 1644511149
transform 1 0 21988 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0836_
timestamp 1644511149
transform 1 0 21988 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0837_
timestamp 1644511149
transform 1 0 21252 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _0838_
timestamp 1644511149
transform 1 0 17204 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0839_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0840_
timestamp 1644511149
transform 1 0 19044 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0841_
timestamp 1644511149
transform 1 0 18952 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0842_
timestamp 1644511149
transform 1 0 17204 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0843_
timestamp 1644511149
transform 1 0 18124 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0844_
timestamp 1644511149
transform 1 0 18216 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0845_
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 1644511149
transform 1 0 17388 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0847_
timestamp 1644511149
transform 1 0 17204 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0848_
timestamp 1644511149
transform 1 0 16652 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0849_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0851_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0852_
timestamp 1644511149
transform 1 0 20700 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0853_
timestamp 1644511149
transform 1 0 19504 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0854_
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0855_
timestamp 1644511149
transform 1 0 21344 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 1644511149
transform 1 0 22080 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0857_
timestamp 1644511149
transform 1 0 20700 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1644511149
transform 1 0 32936 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0859_
timestamp 1644511149
transform 1 0 30176 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0860_
timestamp 1644511149
transform 1 0 28796 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0861_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31280 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0862_
timestamp 1644511149
transform 1 0 32384 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0863_
timestamp 1644511149
transform 1 0 28612 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0864_
timestamp 1644511149
transform 1 0 28152 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0865_
timestamp 1644511149
transform 1 0 27416 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0866_
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0867_
timestamp 1644511149
transform 1 0 30084 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0868_
timestamp 1644511149
transform 1 0 30176 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0869_
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0870_
timestamp 1644511149
transform 1 0 30728 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0871_
timestamp 1644511149
transform 1 0 30452 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0872_
timestamp 1644511149
transform 1 0 31096 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1644511149
transform 1 0 29808 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0874_
timestamp 1644511149
transform 1 0 31556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0875_
timestamp 1644511149
transform 1 0 31004 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0876_
timestamp 1644511149
transform 1 0 32384 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0877_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0878_
timestamp 1644511149
transform 1 0 30360 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0879_
timestamp 1644511149
transform 1 0 29440 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0880_
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0881_
timestamp 1644511149
transform 1 0 29992 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0882_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0883_
timestamp 1644511149
transform 1 0 29808 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0884_
timestamp 1644511149
transform 1 0 30636 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0885_
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0886_
timestamp 1644511149
transform 1 0 26864 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0887_
timestamp 1644511149
transform 1 0 36800 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0888_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37628 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1644511149
transform 1 0 36708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 45540 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 46552 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 43792 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0894_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37536 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 46736 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform 1 0 42688 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 38732 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 25300 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0900_
timestamp 1644511149
transform 1 0 37536 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 20884 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 43332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 11776 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0906_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37536 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 45632 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1644511149
transform 1 0 2208 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 22172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0912_
timestamp 1644511149
transform 1 0 36432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1644511149
transform 1 0 31188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1644511149
transform 1 0 45080 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 35420 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0919_
timestamp 1644511149
transform 1 0 16376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1644511149
transform 1 0 15640 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1644511149
transform 1 0 15456 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 15548 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0925_
timestamp 1644511149
transform 1 0 16836 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 18124 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1644511149
transform 1 0 12604 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 14996 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 14260 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0931_
timestamp 1644511149
transform 1 0 36248 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 20332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 32292 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1644511149
transform 1 0 25392 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0937_
timestamp 1644511149
transform 1 0 36064 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 46736 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 24748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0943_
timestamp 1644511149
transform 1 0 38640 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0944_
timestamp 1644511149
transform 1 0 39376 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 7452 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0950_
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 43148 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0956_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38456 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 33488 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 46276 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 38732 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 32936 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0962_
timestamp 1644511149
transform 1 0 38548 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 5060 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0968_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39376 0 -1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 40296 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 15272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 14628 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 19780 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0974_
timestamp 1644511149
transform 1 0 41124 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0975_
timestamp 1644511149
transform 1 0 19872 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 17664 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 20884 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 8740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0981_
timestamp 1644511149
transform 1 0 25944 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 25300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform 1 0 27600 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1644511149
transform 1 0 28796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 28244 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 24104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0987_
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 46644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 47380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 43332 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0993_
timestamp 1644511149
transform 1 0 20240 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1644511149
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1644511149
transform 1 0 2024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 19780 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0999_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 35788 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1006_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1007_
timestamp 1644511149
transform 1 0 26128 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1644511149
transform 1 0 35604 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36984 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_2  _1012_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _1013_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1014_
timestamp 1644511149
transform 1 0 47656 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1644511149
transform 1 0 44896 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1016_
timestamp 1644511149
transform 1 0 45172 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1017_
timestamp 1644511149
transform 1 0 46644 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1644511149
transform 1 0 46000 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1019_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1644511149
transform 1 0 44252 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1021_
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1022_
timestamp 1644511149
transform 1 0 39836 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1644511149
transform 1 0 40756 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1024_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1025_
timestamp 1644511149
transform 1 0 40296 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1644511149
transform 1 0 40020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1027_
timestamp 1644511149
transform 1 0 40020 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1644511149
transform 1 0 39836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _1029_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21620 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _1030_
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1031_
timestamp 1644511149
transform 1 0 43056 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1032_
timestamp 1644511149
transform 1 0 46184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1033_
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1034_
timestamp 1644511149
transform 1 0 31096 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1035_
timestamp 1644511149
transform 1 0 31004 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1036_
timestamp 1644511149
transform 1 0 30360 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31004 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1038_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1039_
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1040_
timestamp 1644511149
transform 1 0 43884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1041_
timestamp 1644511149
transform 1 0 43700 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1042_
timestamp 1644511149
transform 1 0 43608 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1043_
timestamp 1644511149
transform 1 0 42688 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1044_
timestamp 1644511149
transform 1 0 43976 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1045_
timestamp 1644511149
transform 1 0 43332 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1046_
timestamp 1644511149
transform 1 0 42780 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1047_
timestamp 1644511149
transform 1 0 43056 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1048_
timestamp 1644511149
transform 1 0 42872 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1049_
timestamp 1644511149
transform 1 0 42688 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1050_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42780 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 1644511149
transform 1 0 43884 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1052_
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1053_
timestamp 1644511149
transform 1 0 44436 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1644511149
transform 1 0 45080 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43608 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1056_
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1644511149
transform 1 0 32936 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1058_
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1059_
timestamp 1644511149
transform 1 0 31832 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1060_
timestamp 1644511149
transform 1 0 32752 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 1644511149
transform 1 0 31924 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1062_
timestamp 1644511149
transform 1 0 33396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1063_
timestamp 1644511149
transform 1 0 32292 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1064_
timestamp 1644511149
transform 1 0 32568 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1065_
timestamp 1644511149
transform 1 0 33396 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1066_
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1067_
timestamp 1644511149
transform 1 0 39008 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1068_
timestamp 1644511149
transform 1 0 40020 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1069_
timestamp 1644511149
transform 1 0 32476 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1070_
timestamp 1644511149
transform 1 0 33396 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1071_
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1644511149
transform 1 0 26956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1073_
timestamp 1644511149
transform 1 0 1840 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1644511149
transform 1 0 2760 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1075_
timestamp 1644511149
transform 1 0 46184 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1644511149
transform 1 0 46736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1077_
timestamp 1644511149
transform -1 0 35236 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 1644511149
transform 1 0 34500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1079_
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1080_
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1081_
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1083_
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1084_
timestamp 1644511149
transform 1 0 37076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1085_
timestamp 1644511149
transform 1 0 11868 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1644511149
transform 1 0 28980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1644511149
transform 1 0 30636 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1089_
timestamp 1644511149
transform 1 0 27968 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1644511149
transform 1 0 33672 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1644511149
transform 1 0 33580 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1644511149
transform 1 0 28244 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 33672 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1095_
timestamp 1644511149
transform 1 0 20792 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1644511149
transform 1 0 21620 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1644511149
transform 1 0 19320 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1099_
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1644511149
transform 1 0 17480 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1101_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1644511149
transform 1 0 22080 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1644511149
transform 1 0 22356 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1644511149
transform 1 0 24932 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1105_
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1107_
timestamp 1644511149
transform 1 0 23276 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1644511149
transform 1 0 29348 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1644511149
transform 1 0 30636 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1111_
timestamp 1644511149
transform 1 0 27600 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1113_
timestamp 1644511149
transform 1 0 17940 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1644511149
transform 1 0 20700 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1644511149
transform 1 0 17664 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1644511149
transform 1 0 17940 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1119_
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1120_
timestamp 1644511149
transform 1 0 22816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1644511149
transform 1 0 24748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1123_
timestamp 1644511149
transform 1 0 25392 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27784 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1125_
timestamp 1644511149
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1126_
timestamp 1644511149
transform 1 0 23552 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1128_
timestamp 1644511149
transform 1 0 24748 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1129_
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1130_
timestamp 1644511149
transform 1 0 24104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1131_
timestamp 1644511149
transform 1 0 21620 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1132_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1133_
timestamp 1644511149
transform 1 0 17940 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1134_
timestamp 1644511149
transform 1 0 12144 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1135_
timestamp 1644511149
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1136_
timestamp 1644511149
transform 1 0 16928 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1137_
timestamp 1644511149
transform 1 0 14904 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1138_
timestamp 1644511149
transform 1 0 12604 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1139_
timestamp 1644511149
transform 1 0 12972 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1140_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1141_
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1142_
timestamp 1644511149
transform 1 0 10304 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1143_
timestamp 1644511149
transform 1 0 10672 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1644511149
transform 1 0 10672 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1145_
timestamp 1644511149
transform 1 0 10304 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1146_
timestamp 1644511149
transform 1 0 13248 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1644511149
transform 1 0 13248 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1148_
timestamp 1644511149
transform 1 0 14720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1149_
timestamp 1644511149
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1150_
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1151_
timestamp 1644511149
transform 1 0 17664 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1152_
timestamp 1644511149
transform 1 0 20148 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1153_
timestamp 1644511149
transform 1 0 20240 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1154_
timestamp 1644511149
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1155_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1156_
timestamp 1644511149
transform 1 0 24472 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1157_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1158_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1159_
timestamp 1644511149
transform 1 0 24932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1644511149
transform 1 0 27140 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27140 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1163_
timestamp 1644511149
transform 1 0 29624 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1164_
timestamp 1644511149
transform 1 0 31004 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1165_
timestamp 1644511149
transform 1 0 32844 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1166_
timestamp 1644511149
transform 1 0 31096 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1644511149
transform 1 0 30452 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1644511149
transform 1 0 27048 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1644511149
transform 1 0 32384 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1170_
timestamp 1644511149
transform 1 0 19504 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1644511149
transform 1 0 18400 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 1644511149
transform 1 0 15824 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1173_
timestamp 1644511149
transform 1 0 15732 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1175_
timestamp 1644511149
transform 1 0 19412 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 1644511149
transform 1 0 23552 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1178_
timestamp 1644511149
transform 1 0 27140 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1179_
timestamp 1644511149
transform 1 0 27232 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1180_
timestamp 1644511149
transform 1 0 28152 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1181_
timestamp 1644511149
transform 1 0 29808 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 1644511149
transform 1 0 24656 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 1644511149
transform 1 0 25944 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 1644511149
transform 1 0 22448 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 1644511149
transform 1 0 19504 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1187_
timestamp 1644511149
transform 1 0 16836 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1188_
timestamp 1644511149
transform 1 0 16928 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1189_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1644511149
transform 1 0 22632 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1644511149
transform 1 0 24380 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1194_
timestamp 1644511149
transform 1 0 27140 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27600 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1196_
timestamp 1644511149
transform 1 0 24104 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1197_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1199_
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1200_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1201_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1202_
timestamp 1644511149
transform 1 0 17572 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1203_
timestamp 1644511149
transform 1 0 17572 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1204_
timestamp 1644511149
transform 1 0 17480 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1205_
timestamp 1644511149
transform 1 0 14996 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1206_
timestamp 1644511149
transform 1 0 12420 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1644511149
transform 1 0 13064 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1208_
timestamp 1644511149
transform 1 0 11040 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 1644511149
transform 1 0 10396 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1210_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1211_
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1644511149
transform 1 0 10304 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 1644511149
transform 1 0 12512 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1214_
timestamp 1644511149
transform 1 0 14168 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1215_
timestamp 1644511149
transform 1 0 14352 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1216_
timestamp 1644511149
transform 1 0 18032 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1217_
timestamp 1644511149
transform 1 0 18032 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1218_
timestamp 1644511149
transform 1 0 19412 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1644511149
transform 1 0 21712 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1220_
timestamp 1644511149
transform 1 0 21528 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1221_
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1222_
timestamp 1644511149
transform 1 0 29440 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1223_
timestamp 1644511149
transform 1 0 27692 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1224_
timestamp 1644511149
transform 1 0 25576 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1225_
timestamp 1644511149
transform 1 0 27508 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1226_
timestamp 1644511149
transform 1 0 22724 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1227__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1228__82
timestamp 1644511149
transform 1 0 32292 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1229__83
timestamp 1644511149
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1230__84
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1231__85
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1232__86
timestamp 1644511149
transform 1 0 20792 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1233__87
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1234__88
timestamp 1644511149
transform 1 0 24656 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1235__89
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1236__90
timestamp 1644511149
transform 1 0 25300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1237__91
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1238__92
timestamp 1644511149
transform 1 0 1840 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1239__93
timestamp 1644511149
transform 1 0 33672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1240__94
timestamp 1644511149
transform 1 0 4324 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1241__95
timestamp 1644511149
transform 1 0 1472 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1242__96
timestamp 1644511149
transform 1 0 43976 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1243__97
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1244__98
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1245__99
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1246__100
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1247__101
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1248__102
timestamp 1644511149
transform 1 0 7268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1249__103
timestamp 1644511149
transform 1 0 41124 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1250__104
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1251__105
timestamp 1644511149
transform 1 0 47472 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1252__106
timestamp 1644511149
transform 1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1253__107
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1254__108
timestamp 1644511149
transform 1 0 45908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1255__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1256__110
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1257__111
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1258__112
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1259__113
timestamp 1644511149
transform 1 0 41308 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1260__114
timestamp 1644511149
transform 1 0 45264 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1261__115
timestamp 1644511149
transform 1 0 25392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1262__116
timestamp 1644511149
transform 1 0 42504 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1263__117
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1264__118
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1265__119
timestamp 1644511149
transform 1 0 6716 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1266__120
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1267__121
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1268__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1269__123
timestamp 1644511149
transform 1 0 47472 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1270__124
timestamp 1644511149
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1271__125
timestamp 1644511149
transform 1 0 44896 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1272__126
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1273__127
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1274__128
timestamp 1644511149
transform 1 0 47472 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1275__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1276__130
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1277__131
timestamp 1644511149
transform 1 0 1840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1278__132
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1279__133
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1280__134
timestamp 1644511149
transform 1 0 47472 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1281__135
timestamp 1644511149
transform 1 0 43884 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34868 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1283_
timestamp 1644511149
transform 1 0 33304 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1284_
timestamp 1644511149
transform 1 0 43700 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1285_
timestamp 1644511149
transform 1 0 44712 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1286_
timestamp 1644511149
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1644511149
transform 1 0 42596 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1644511149
transform 1 0 45172 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1644511149
transform 1 0 39376 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1644511149
transform 1 0 38640 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1644511149
transform 1 0 32200 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1644511149
transform 1 0 19320 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1644511149
transform 1 0 20792 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1644511149
transform 1 0 25208 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1644511149
transform 1 0 1748 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1644511149
transform 1 0 32936 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1644511149
transform 1 0 3956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1309_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1310_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1311_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1312_
timestamp 1644511149
transform 1 0 7176 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1313_
timestamp 1644511149
transform 1 0 41032 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1314_
timestamp 1644511149
transform 1 0 37352 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1315_
timestamp 1644511149
transform 1 0 36156 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1316_
timestamp 1644511149
transform 1 0 22080 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1317_
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1318_
timestamp 1644511149
transform 1 0 15272 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1319_
timestamp 1644511149
transform 1 0 30360 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1320_
timestamp 1644511149
transform 1 0 14996 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1321_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1322_
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1323_
timestamp 1644511149
transform 1 0 19688 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1324_
timestamp 1644511149
transform 1 0 18124 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1325_
timestamp 1644511149
transform 1 0 15548 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1326_
timestamp 1644511149
transform 1 0 13340 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1327_
timestamp 1644511149
transform 1 0 15732 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1328_
timestamp 1644511149
transform 1 0 13524 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1329_
timestamp 1644511149
transform 1 0 8464 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1330_
timestamp 1644511149
transform 1 0 14260 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1331_
timestamp 1644511149
transform 1 0 16560 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1332_
timestamp 1644511149
transform 1 0 8372 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1333_
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1334_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1335_
timestamp 1644511149
transform 1 0 17572 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1336_
timestamp 1644511149
transform 1 0 20240 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1337_
timestamp 1644511149
transform 1 0 14996 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1338_
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1339_
timestamp 1644511149
transform 1 0 25208 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1340_
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1341_
timestamp 1644511149
transform 1 0 27140 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1342_
timestamp 1644511149
transform 1 0 32200 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1343_
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1344_
timestamp 1644511149
transform 1 0 25300 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1345_
timestamp 1644511149
transform 1 0 27508 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1346_
timestamp 1644511149
transform 1 0 9108 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1347_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1348_
timestamp 1644511149
transform 1 0 23184 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1349_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1350_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1351_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1352_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1353_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1354_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1355_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1356_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1357_
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1358_
timestamp 1644511149
transform 1 0 42688 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1359_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1360_
timestamp 1644511149
transform 1 0 13800 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1361_
timestamp 1644511149
transform 1 0 6532 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1362_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1363_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1364_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1365_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1366_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1367_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1368_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1369_
timestamp 1644511149
transform 1 0 13616 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1370_
timestamp 1644511149
transform 1 0 45172 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1371_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1372_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1373_
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1374_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1375_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1376_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1377_
timestamp 1644511149
transform 1 0 44988 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 24932 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 22816 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 22908 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 22632 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 27416 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 28428 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 47840 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 47932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1644511149
transform 1 0 19596 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1644511149
transform 1 0 47288 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 47932 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 45632 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 41584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 39192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1644511149
transform 1 0 46736 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 47656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1644511149
transform 1 0 47748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 47656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1644511149
transform 1 0 9292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1644511149
transform 1 0 12328 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 22448 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 14812 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1644511149
transform 1 0 46552 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 30728 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 43148 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1644511149
transform 1 0 11684 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 46184 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform 1 0 26128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 45632 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 47840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40480 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 41032 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 39192 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 39928 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 41124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 39744 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 40388 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 13248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 14720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 14168 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 15824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 15364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 17296 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 17940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  instrumented_adder.tristate_ext_inputs\[0\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33304 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[1\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2116 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 46920 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 34500 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37076 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 31280 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2576 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45356 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35144 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 46736 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42504 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37536 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 35420 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 34684 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 45816 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 45356 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 40020 0 1 22848
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
