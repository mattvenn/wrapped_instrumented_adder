magic
tech sky130A
magscale 1 2
timestamp 1654258224
<< viali >>
rect 13369 47209 13403 47243
rect 9597 47141 9631 47175
rect 29929 47141 29963 47175
rect 48145 47141 48179 47175
rect 2053 47073 2087 47107
rect 6653 47073 6687 47107
rect 20085 47073 20119 47107
rect 47041 47073 47075 47107
rect 1777 47005 1811 47039
rect 3801 47005 3835 47039
rect 4721 47005 4755 47039
rect 6377 47005 6411 47039
rect 7297 47005 7331 47039
rect 9413 47005 9447 47039
rect 11621 47005 11655 47039
rect 12357 47005 12391 47039
rect 13093 47005 13127 47039
rect 16681 47005 16715 47039
rect 16957 47005 16991 47039
rect 18337 47005 18371 47039
rect 20361 47005 20395 47039
rect 24869 47005 24903 47039
rect 25513 47005 25547 47039
rect 28549 47005 28583 47039
rect 29745 47005 29779 47039
rect 31125 47005 31159 47039
rect 38393 47005 38427 47039
rect 42717 47005 42751 47039
rect 43177 47005 43211 47039
rect 44005 47005 44039 47039
rect 45201 47005 45235 47039
rect 47961 47005 47995 47039
rect 2789 46937 2823 46971
rect 3157 46937 3191 46971
rect 4077 46937 4111 46971
rect 4997 46937 5031 46971
rect 11805 46937 11839 46971
rect 12541 46937 12575 46971
rect 14565 46937 14599 46971
rect 14749 46937 14783 46971
rect 18705 46937 18739 46971
rect 28733 46937 28767 46971
rect 31309 46937 31343 46971
rect 40325 46937 40359 46971
rect 40509 46937 40543 46971
rect 44189 46937 44223 46971
rect 45385 46937 45419 46971
rect 7481 46869 7515 46903
rect 43361 46869 43395 46903
rect 1869 46597 1903 46631
rect 44557 46597 44591 46631
rect 47041 46597 47075 46631
rect 24593 46529 24627 46563
rect 38209 46529 38243 46563
rect 42717 46529 42751 46563
rect 47961 46529 47995 46563
rect 3433 46461 3467 46495
rect 3617 46461 3651 46495
rect 4169 46461 4203 46495
rect 13093 46461 13127 46495
rect 13553 46461 13587 46495
rect 13737 46461 13771 46495
rect 14289 46461 14323 46495
rect 19441 46461 19475 46495
rect 19625 46461 19659 46495
rect 20637 46461 20671 46495
rect 24777 46461 24811 46495
rect 25145 46461 25179 46495
rect 32413 46461 32447 46495
rect 32597 46461 32631 46495
rect 33425 46461 33459 46495
rect 38393 46461 38427 46495
rect 38669 46461 38703 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 2145 46325 2179 46359
rect 2881 46325 2915 46359
rect 10793 46325 10827 46359
rect 22017 46325 22051 46359
rect 41613 46325 41647 46359
rect 48053 46325 48087 46359
rect 3893 46121 3927 46155
rect 4629 46121 4663 46155
rect 14197 46121 14231 46155
rect 20361 46121 20395 46155
rect 24685 46121 24719 46155
rect 32689 46121 32723 46155
rect 38393 46121 38427 46155
rect 43821 46121 43855 46155
rect 10517 45985 10551 46019
rect 11069 45985 11103 46019
rect 20821 45985 20855 46019
rect 21281 45985 21315 46019
rect 25237 45985 25271 46019
rect 26617 45985 26651 46019
rect 41429 45985 41463 46019
rect 42533 45985 42567 46019
rect 46305 45985 46339 46019
rect 48145 45985 48179 46019
rect 2881 45917 2915 45951
rect 3801 45917 3835 45951
rect 14105 45917 14139 45951
rect 24593 45917 24627 45951
rect 38301 45917 38335 45951
rect 43729 45917 43763 45951
rect 45661 45917 45695 45951
rect 10701 45849 10735 45883
rect 21005 45849 21039 45883
rect 25421 45849 25455 45883
rect 41613 45849 41647 45883
rect 46489 45849 46523 45883
rect 2973 45781 3007 45815
rect 45753 45781 45787 45815
rect 10701 45577 10735 45611
rect 20361 45577 20395 45611
rect 21005 45577 21039 45611
rect 25421 45577 25455 45611
rect 2237 45509 2271 45543
rect 33333 45509 33367 45543
rect 41061 45509 41095 45543
rect 43913 45509 43947 45543
rect 44649 45509 44683 45543
rect 46857 45509 46891 45543
rect 10609 45441 10643 45475
rect 20269 45441 20303 45475
rect 20913 45441 20947 45475
rect 25329 45441 25363 45475
rect 33241 45441 33275 45475
rect 40969 45441 41003 45475
rect 43821 45441 43855 45475
rect 47593 45441 47627 45475
rect 2053 45373 2087 45407
rect 2973 45373 3007 45407
rect 38669 45373 38703 45407
rect 38853 45373 38887 45407
rect 39865 45373 39899 45407
rect 44465 45373 44499 45407
rect 45845 45373 45879 45407
rect 47685 45305 47719 45339
rect 41797 45237 41831 45271
rect 46949 45237 46983 45271
rect 38853 45033 38887 45067
rect 44465 45033 44499 45067
rect 45109 45033 45143 45067
rect 41429 44897 41463 44931
rect 42901 44897 42935 44931
rect 48145 44897 48179 44931
rect 28733 44829 28767 44863
rect 38761 44829 38795 44863
rect 45017 44829 45051 44863
rect 45661 44829 45695 44863
rect 46305 44829 46339 44863
rect 41613 44761 41647 44795
rect 45753 44761 45787 44795
rect 46489 44761 46523 44795
rect 28825 44693 28859 44727
rect 41613 44489 41647 44523
rect 46949 44489 46983 44523
rect 41521 44353 41555 44387
rect 45661 44353 45695 44387
rect 46397 44353 46431 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 47685 44149 47719 44183
rect 45845 43945 45879 43979
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 46305 43741 46339 43775
rect 1409 43265 1443 43299
rect 47041 43265 47075 43299
rect 1593 43197 1627 43231
rect 47777 43197 47811 43231
rect 46305 42653 46339 42687
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 47685 42313 47719 42347
rect 47041 42177 47075 42211
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 48145 41565 48179 41599
rect 1593 41497 1627 41531
rect 46489 41497 46523 41531
rect 2237 41225 2271 41259
rect 46949 41225 46983 41259
rect 2145 41089 2179 41123
rect 46857 41089 46891 41123
rect 47961 41089 47995 41123
rect 48053 40885 48087 40919
rect 47685 40681 47719 40715
rect 1409 40477 1443 40511
rect 1593 40341 1627 40375
rect 47777 39797 47811 39831
rect 40233 39457 40267 39491
rect 46305 39457 46339 39491
rect 48145 39457 48179 39491
rect 39957 39389 39991 39423
rect 46489 39321 46523 39355
rect 46949 39049 46983 39083
rect 40141 38913 40175 38947
rect 46857 38913 46891 38947
rect 47685 38913 47719 38947
rect 40417 38845 40451 38879
rect 47869 38845 47903 38879
rect 41981 38369 42015 38403
rect 39037 38301 39071 38335
rect 46305 38301 46339 38335
rect 40233 38233 40267 38267
rect 46489 38233 46523 38267
rect 48145 38233 48179 38267
rect 39221 38165 39255 38199
rect 47685 37961 47719 37995
rect 40141 37825 40175 37859
rect 47593 37825 47627 37859
rect 40417 37757 40451 37791
rect 47685 37417 47719 37451
rect 2237 37213 2271 37247
rect 25697 37213 25731 37247
rect 40141 37213 40175 37247
rect 25881 37145 25915 37179
rect 40509 37145 40543 37179
rect 26065 37077 26099 37111
rect 27353 36873 27387 36907
rect 1961 36737 1995 36771
rect 23213 36737 23247 36771
rect 26065 36737 26099 36771
rect 2145 36669 2179 36703
rect 2973 36669 3007 36703
rect 26157 36669 26191 36703
rect 26433 36669 26467 36703
rect 27445 36669 27479 36703
rect 27537 36669 27571 36703
rect 26985 36601 27019 36635
rect 23029 36533 23063 36567
rect 2881 36329 2915 36363
rect 22109 36193 22143 36227
rect 2789 36125 2823 36159
rect 24409 36125 24443 36159
rect 28549 36125 28583 36159
rect 33425 36125 33459 36159
rect 22385 36057 22419 36091
rect 24685 36057 24719 36091
rect 23857 35989 23891 36023
rect 26157 35989 26191 36023
rect 28641 35989 28675 36023
rect 33241 35989 33275 36023
rect 22661 35785 22695 35819
rect 25605 35785 25639 35819
rect 33333 35785 33367 35819
rect 33701 35785 33735 35819
rect 29653 35717 29687 35751
rect 1593 35649 1627 35683
rect 22569 35649 22603 35683
rect 24409 35649 24443 35683
rect 25973 35649 26007 35683
rect 25789 35581 25823 35615
rect 25881 35581 25915 35615
rect 26065 35581 26099 35615
rect 27169 35581 27203 35615
rect 27445 35581 27479 35615
rect 29377 35581 29411 35615
rect 33793 35581 33827 35615
rect 33885 35581 33919 35615
rect 1409 35445 1443 35479
rect 24593 35445 24627 35479
rect 28917 35445 28951 35479
rect 31125 35445 31159 35479
rect 24777 35241 24811 35275
rect 26065 35241 26099 35275
rect 26433 35241 26467 35275
rect 27169 35241 27203 35275
rect 28089 35241 28123 35275
rect 30481 35241 30515 35275
rect 33517 35241 33551 35275
rect 27353 35173 27387 35207
rect 25605 35105 25639 35139
rect 33057 35105 33091 35139
rect 20545 35037 20579 35071
rect 24685 35037 24719 35071
rect 25329 35037 25363 35071
rect 25421 35037 25455 35071
rect 26249 35037 26283 35071
rect 26525 35037 26559 35071
rect 30389 35037 30423 35071
rect 31033 35037 31067 35071
rect 33149 35037 33183 35071
rect 48145 35037 48179 35071
rect 26985 34969 27019 35003
rect 27997 34969 28031 35003
rect 20729 34901 20763 34935
rect 25329 34901 25363 34935
rect 27185 34901 27219 34935
rect 31125 34901 31159 34935
rect 47961 34901 47995 34935
rect 29009 34697 29043 34731
rect 29285 34697 29319 34731
rect 29469 34697 29503 34731
rect 31125 34697 31159 34731
rect 30757 34629 30791 34663
rect 30973 34629 31007 34663
rect 33333 34629 33367 34663
rect 22109 34561 22143 34595
rect 25697 34561 25731 34595
rect 25973 34561 26007 34595
rect 29466 34561 29500 34595
rect 29837 34561 29871 34595
rect 29929 34561 29963 34595
rect 48145 34561 48179 34595
rect 22201 34493 22235 34527
rect 23489 34493 23523 34527
rect 23765 34493 23799 34527
rect 25237 34493 25271 34527
rect 25789 34493 25823 34527
rect 33057 34493 33091 34527
rect 34805 34493 34839 34527
rect 25973 34357 26007 34391
rect 26157 34357 26191 34391
rect 30941 34357 30975 34391
rect 47961 34357 47995 34391
rect 24685 34153 24719 34187
rect 26065 34153 26099 34187
rect 29929 34153 29963 34187
rect 34805 34153 34839 34187
rect 26249 34085 26283 34119
rect 21373 34017 21407 34051
rect 25973 34017 26007 34051
rect 28457 34017 28491 34051
rect 30481 34017 30515 34051
rect 20545 33949 20579 33983
rect 24593 33949 24627 33983
rect 25881 33949 25915 33983
rect 28181 33949 28215 33983
rect 28273 33949 28307 33983
rect 29837 33949 29871 33983
rect 30021 33949 30055 33983
rect 34713 33949 34747 33983
rect 47869 33949 47903 33983
rect 21649 33881 21683 33915
rect 28457 33881 28491 33915
rect 30757 33881 30791 33915
rect 20637 33813 20671 33847
rect 23121 33813 23155 33847
rect 32229 33813 32263 33847
rect 48053 33813 48087 33847
rect 22569 33609 22603 33643
rect 24961 33609 24995 33643
rect 28457 33609 28491 33643
rect 29285 33609 29319 33643
rect 32597 33609 32631 33643
rect 15853 33541 15887 33575
rect 25605 33541 25639 33575
rect 29837 33541 29871 33575
rect 30757 33541 30791 33575
rect 32137 33541 32171 33575
rect 1961 33473 1995 33507
rect 19533 33473 19567 33507
rect 21833 33473 21867 33507
rect 22017 33473 22051 33507
rect 22109 33473 22143 33507
rect 22385 33473 22419 33507
rect 24777 33473 24811 33507
rect 25789 33473 25823 33507
rect 27721 33473 27755 33507
rect 27905 33473 27939 33507
rect 28273 33473 28307 33507
rect 29561 33473 29595 33507
rect 30389 33473 30423 33507
rect 30573 33473 30607 33507
rect 32413 33473 32447 33507
rect 33057 33473 33091 33507
rect 35357 33473 35391 33507
rect 47041 33473 47075 33507
rect 47593 33473 47627 33507
rect 2145 33405 2179 33439
rect 3801 33405 3835 33439
rect 14013 33405 14047 33439
rect 14197 33405 14231 33439
rect 19809 33405 19843 33439
rect 22201 33405 22235 33439
rect 24317 33405 24351 33439
rect 24685 33405 24719 33439
rect 27997 33405 28031 33439
rect 28089 33405 28123 33439
rect 29469 33405 29503 33439
rect 29929 33405 29963 33439
rect 32321 33405 32355 33439
rect 33333 33405 33367 33439
rect 48053 33405 48087 33439
rect 21281 33269 21315 33303
rect 25973 33269 26007 33303
rect 32137 33269 32171 33303
rect 33149 33269 33183 33303
rect 33241 33269 33275 33303
rect 35449 33269 35483 33303
rect 46857 33269 46891 33303
rect 47869 33269 47903 33303
rect 2789 33065 2823 33099
rect 3801 33065 3835 33099
rect 22661 33065 22695 33099
rect 25053 33065 25087 33099
rect 25881 33065 25915 33099
rect 28365 33065 28399 33099
rect 28825 33065 28859 33099
rect 31033 33065 31067 33099
rect 32505 33065 32539 33099
rect 21465 32997 21499 33031
rect 26157 32997 26191 33031
rect 27261 32997 27295 33031
rect 32873 32997 32907 33031
rect 1409 32929 1443 32963
rect 3157 32929 3191 32963
rect 14105 32929 14139 32963
rect 15945 32929 15979 32963
rect 21189 32929 21223 32963
rect 22201 32929 22235 32963
rect 22293 32929 22327 32963
rect 25789 32929 25823 32963
rect 26801 32929 26835 32963
rect 30573 32929 30607 32963
rect 47133 32929 47167 32963
rect 47409 32929 47443 32963
rect 1685 32861 1719 32895
rect 2697 32861 2731 32895
rect 3985 32861 4019 32895
rect 13369 32861 13403 32895
rect 21097 32861 21131 32895
rect 21925 32861 21959 32895
rect 22109 32861 22143 32895
rect 22477 32861 22511 32895
rect 24869 32861 24903 32895
rect 25145 32861 25179 32895
rect 25973 32861 26007 32895
rect 26893 32861 26927 32895
rect 27997 32861 28031 32895
rect 28181 32861 28215 32895
rect 28825 32861 28859 32895
rect 29009 32861 29043 32895
rect 29101 32861 29135 32895
rect 30297 32861 30331 32895
rect 30481 32861 30515 32895
rect 30665 32861 30699 32895
rect 30849 32861 30883 32895
rect 32505 32861 32539 32895
rect 32689 32861 32723 32895
rect 34713 32861 34747 32895
rect 46581 32861 46615 32895
rect 13461 32793 13495 32827
rect 14289 32793 14323 32827
rect 25697 32793 25731 32827
rect 30021 32793 30055 32827
rect 33793 32793 33827 32827
rect 33977 32793 34011 32827
rect 34989 32793 35023 32827
rect 47225 32793 47259 32827
rect 24685 32725 24719 32759
rect 29285 32725 29319 32759
rect 34161 32725 34195 32759
rect 36461 32725 36495 32759
rect 2789 32453 2823 32487
rect 14105 32453 14139 32487
rect 20913 32453 20947 32487
rect 21281 32453 21315 32487
rect 22017 32453 22051 32487
rect 22201 32453 22235 32487
rect 25145 32453 25179 32487
rect 27169 32453 27203 32487
rect 29929 32453 29963 32487
rect 35173 32453 35207 32487
rect 14013 32385 14047 32419
rect 21097 32385 21131 32419
rect 21833 32385 21867 32419
rect 25421 32385 25455 32419
rect 26985 32385 27019 32419
rect 28365 32385 28399 32419
rect 29009 32385 29043 32419
rect 30113 32385 30147 32419
rect 30205 32385 30239 32419
rect 30389 32385 30423 32419
rect 30481 32385 30515 32419
rect 31033 32385 31067 32419
rect 32321 32385 32355 32419
rect 33333 32385 33367 32419
rect 33517 32385 33551 32419
rect 34437 32385 34471 32419
rect 34621 32385 34655 32419
rect 34989 32385 35023 32419
rect 46489 32385 46523 32419
rect 47593 32385 47627 32419
rect 2605 32317 2639 32351
rect 4445 32317 4479 32351
rect 9137 32317 9171 32351
rect 9321 32317 9355 32351
rect 10517 32317 10551 32351
rect 11529 32317 11563 32351
rect 11805 32317 11839 32351
rect 13277 32317 13311 32351
rect 25329 32317 25363 32351
rect 28549 32317 28583 32351
rect 32229 32317 32263 32351
rect 33425 32317 33459 32351
rect 34713 32317 34747 32351
rect 34805 32317 34839 32351
rect 46213 32317 46247 32351
rect 25605 32249 25639 32283
rect 27353 32249 27387 32283
rect 2145 32181 2179 32215
rect 25421 32181 25455 32215
rect 29193 32181 29227 32215
rect 31217 32181 31251 32215
rect 32689 32181 32723 32215
rect 47685 32181 47719 32215
rect 1409 31977 1443 32011
rect 9781 31977 9815 32011
rect 10793 31977 10827 32011
rect 11805 31977 11839 32011
rect 12633 31977 12667 32011
rect 15117 31977 15151 32011
rect 21465 31977 21499 32011
rect 22753 31977 22787 32011
rect 22937 31977 22971 32011
rect 26893 31977 26927 32011
rect 27629 31977 27663 32011
rect 28549 31977 28583 32011
rect 31861 31909 31895 31943
rect 32781 31909 32815 31943
rect 11621 31841 11655 31875
rect 13277 31841 13311 31875
rect 14565 31841 14599 31875
rect 31401 31841 31435 31875
rect 46305 31841 46339 31875
rect 46489 31841 46523 31875
rect 48145 31841 48179 31875
rect 1593 31773 1627 31807
rect 2881 31773 2915 31807
rect 9689 31773 9723 31807
rect 10701 31773 10735 31807
rect 11529 31773 11563 31807
rect 12541 31773 12575 31807
rect 13185 31773 13219 31807
rect 13369 31773 13403 31807
rect 14289 31773 14323 31807
rect 14473 31773 14507 31807
rect 15025 31773 15059 31807
rect 19993 31773 20027 31807
rect 20085 31773 20119 31807
rect 21281 31773 21315 31807
rect 21373 31773 21407 31807
rect 22385 31773 22419 31807
rect 22753 31773 22787 31807
rect 24685 31773 24719 31807
rect 24961 31773 24995 31807
rect 25697 31773 25731 31807
rect 26065 31773 26099 31807
rect 26801 31773 26835 31807
rect 28733 31773 28767 31807
rect 31309 31773 31343 31807
rect 31493 31773 31527 31807
rect 32137 31773 32171 31807
rect 32285 31773 32319 31807
rect 32413 31773 32447 31807
rect 32505 31773 32539 31807
rect 32643 31773 32677 31807
rect 34713 31773 34747 31807
rect 34805 31773 34839 31807
rect 24869 31705 24903 31739
rect 25881 31705 25915 31739
rect 25973 31705 26007 31739
rect 27537 31705 27571 31739
rect 2973 31637 3007 31671
rect 14105 31637 14139 31671
rect 21649 31637 21683 31671
rect 24501 31637 24535 31671
rect 26249 31637 26283 31671
rect 15485 31433 15519 31467
rect 20637 31433 20671 31467
rect 23581 31433 23615 31467
rect 34713 31433 34747 31467
rect 2237 31365 2271 31399
rect 14013 31365 14047 31399
rect 46121 31365 46155 31399
rect 2053 31297 2087 31331
rect 10885 31297 10919 31331
rect 12265 31297 12299 31331
rect 15945 31297 15979 31331
rect 16681 31297 16715 31331
rect 21097 31297 21131 31331
rect 21925 31297 21959 31331
rect 23397 31297 23431 31331
rect 23673 31297 23707 31331
rect 24133 31297 24167 31331
rect 32965 31297 32999 31331
rect 2789 31229 2823 31263
rect 13737 31229 13771 31263
rect 16037 31229 16071 31263
rect 18889 31229 18923 31263
rect 19165 31229 19199 31263
rect 22201 31229 22235 31263
rect 24409 31229 24443 31263
rect 33241 31229 33275 31263
rect 46029 31229 46063 31263
rect 46857 31229 46891 31263
rect 10885 31093 10919 31127
rect 12357 31093 12391 31127
rect 16773 31093 16807 31127
rect 21189 31093 21223 31127
rect 23213 31093 23247 31127
rect 25881 31093 25915 31127
rect 21005 30889 21039 30923
rect 22293 30889 22327 30923
rect 22937 30889 22971 30923
rect 25697 30889 25731 30923
rect 26341 30889 26375 30923
rect 28549 30889 28583 30923
rect 29561 30889 29595 30923
rect 30021 30889 30055 30923
rect 13001 30821 13035 30855
rect 23305 30821 23339 30855
rect 10793 30753 10827 30787
rect 14657 30753 14691 30787
rect 17417 30753 17451 30787
rect 19257 30753 19291 30787
rect 25513 30753 25547 30787
rect 29653 30753 29687 30787
rect 35265 30753 35299 30787
rect 13277 30685 13311 30719
rect 14749 30685 14783 30719
rect 15669 30685 15703 30719
rect 21925 30685 21959 30719
rect 22293 30685 22327 30719
rect 23121 30685 23155 30719
rect 23397 30685 23431 30719
rect 25421 30685 25455 30719
rect 26249 30685 26283 30719
rect 28181 30685 28215 30719
rect 29837 30685 29871 30719
rect 30573 30685 30607 30719
rect 30757 30685 30791 30719
rect 32137 30685 32171 30719
rect 33793 30685 33827 30719
rect 34161 30685 34195 30719
rect 34897 30685 34931 30719
rect 35081 30685 35115 30719
rect 35173 30685 35207 30719
rect 35449 30685 35483 30719
rect 11069 30617 11103 30651
rect 13369 30617 13403 30651
rect 15945 30617 15979 30651
rect 19533 30617 19567 30651
rect 24593 30617 24627 30651
rect 28365 30617 28399 30651
rect 29561 30617 29595 30651
rect 31493 30617 31527 30651
rect 33977 30617 34011 30651
rect 12541 30549 12575 30583
rect 13185 30549 13219 30583
rect 13553 30549 13587 30583
rect 15117 30549 15151 30583
rect 22477 30549 22511 30583
rect 24685 30549 24719 30583
rect 30665 30549 30699 30583
rect 31585 30549 31619 30583
rect 32229 30549 32263 30583
rect 35633 30549 35667 30583
rect 11713 30345 11747 30379
rect 14289 30345 14323 30379
rect 15761 30345 15795 30379
rect 24317 30345 24351 30379
rect 34529 30345 34563 30379
rect 12265 30277 12299 30311
rect 12541 30277 12575 30311
rect 21189 30277 21223 30311
rect 26249 30277 26283 30311
rect 33149 30277 33183 30311
rect 35265 30277 35299 30311
rect 10609 30209 10643 30243
rect 10701 30209 10735 30243
rect 10977 30209 11011 30243
rect 11621 30209 11655 30243
rect 11805 30209 11839 30243
rect 12449 30209 12483 30243
rect 12633 30209 12667 30243
rect 14105 30209 14139 30243
rect 14289 30209 14323 30243
rect 15577 30209 15611 30243
rect 20913 30209 20947 30243
rect 21005 30209 21039 30243
rect 21925 30209 21959 30243
rect 22109 30209 22143 30243
rect 22201 30209 22235 30243
rect 22477 30209 22511 30243
rect 24258 30209 24292 30243
rect 24685 30209 24719 30243
rect 25421 30209 25455 30243
rect 26065 30209 26099 30243
rect 27537 30209 27571 30243
rect 28549 30209 28583 30243
rect 29837 30209 29871 30243
rect 33333 30209 33367 30243
rect 34161 30209 34195 30243
rect 10793 30141 10827 30175
rect 12817 30141 12851 30175
rect 20545 30141 20579 30175
rect 22293 30141 22327 30175
rect 24777 30141 24811 30175
rect 27445 30141 27479 30175
rect 28825 30141 28859 30175
rect 30113 30141 30147 30175
rect 34069 30141 34103 30175
rect 34989 30141 35023 30175
rect 10977 30073 11011 30107
rect 22661 30073 22695 30107
rect 24133 30073 24167 30107
rect 26433 30073 26467 30107
rect 23765 30005 23799 30039
rect 25513 30005 25547 30039
rect 27905 30005 27939 30039
rect 31585 30005 31619 30039
rect 33517 30005 33551 30039
rect 36737 30005 36771 30039
rect 21281 29801 21315 29835
rect 21833 29801 21867 29835
rect 24961 29801 24995 29835
rect 29009 29801 29043 29835
rect 30573 29801 30607 29835
rect 31033 29801 31067 29835
rect 32137 29801 32171 29835
rect 34713 29801 34747 29835
rect 35173 29801 35207 29835
rect 35909 29801 35943 29835
rect 31493 29733 31527 29767
rect 9321 29665 9355 29699
rect 21925 29665 21959 29699
rect 27261 29665 27295 29699
rect 30113 29665 30147 29699
rect 31217 29665 31251 29699
rect 33333 29665 33367 29699
rect 34897 29665 34931 29699
rect 47593 29665 47627 29699
rect 15393 29597 15427 29631
rect 15669 29597 15703 29631
rect 16129 29597 16163 29631
rect 21462 29597 21496 29631
rect 24777 29597 24811 29631
rect 25145 29597 25179 29631
rect 25789 29597 25823 29631
rect 25973 29597 26007 29631
rect 26157 29597 26191 29631
rect 26249 29597 26283 29631
rect 29837 29597 29871 29631
rect 30021 29597 30055 29631
rect 30205 29597 30239 29631
rect 30389 29597 30423 29631
rect 31309 29597 31343 29631
rect 32045 29597 32079 29631
rect 32413 29597 32447 29631
rect 33057 29597 33091 29631
rect 33241 29597 33275 29631
rect 33425 29597 33459 29631
rect 33609 29597 33643 29631
rect 34989 29597 35023 29631
rect 35817 29597 35851 29631
rect 47317 29597 47351 29631
rect 9505 29529 9539 29563
rect 11161 29529 11195 29563
rect 16405 29529 16439 29563
rect 27537 29529 27571 29563
rect 31033 29529 31067 29563
rect 34713 29529 34747 29563
rect 17877 29461 17911 29495
rect 21465 29461 21499 29495
rect 25329 29461 25363 29495
rect 32597 29461 32631 29495
rect 33793 29461 33827 29495
rect 9689 29257 9723 29291
rect 16957 29257 16991 29291
rect 29193 29257 29227 29291
rect 32321 29257 32355 29291
rect 33149 29257 33183 29291
rect 36001 29257 36035 29291
rect 13461 29189 13495 29223
rect 21833 29189 21867 29223
rect 32229 29189 32263 29223
rect 34529 29189 34563 29223
rect 9597 29121 9631 29155
rect 14105 29121 14139 29155
rect 15393 29121 15427 29155
rect 16865 29121 16899 29155
rect 22017 29121 22051 29155
rect 24317 29121 24351 29155
rect 27905 29121 27939 29155
rect 30665 29121 30699 29155
rect 30849 29121 30883 29155
rect 33333 29121 33367 29155
rect 34253 29121 34287 29155
rect 15485 29053 15519 29087
rect 15761 29053 15795 29087
rect 33517 29053 33551 29087
rect 33609 29053 33643 29087
rect 13645 28985 13679 29019
rect 14289 28985 14323 29019
rect 26065 28985 26099 29019
rect 31033 28985 31067 29019
rect 22201 28917 22235 28951
rect 24580 28917 24614 28951
rect 30665 28917 30699 28951
rect 14473 28713 14507 28747
rect 25881 28713 25915 28747
rect 27997 28713 28031 28747
rect 28733 28713 28767 28747
rect 30113 28713 30147 28747
rect 30757 28713 30791 28747
rect 32321 28713 32355 28747
rect 33517 28713 33551 28747
rect 34897 28713 34931 28747
rect 35541 28713 35575 28747
rect 28917 28645 28951 28679
rect 30665 28645 30699 28679
rect 10241 28577 10275 28611
rect 10517 28577 10551 28611
rect 11253 28577 11287 28611
rect 13001 28577 13035 28611
rect 16037 28577 16071 28611
rect 19533 28577 19567 28611
rect 24777 28577 24811 28611
rect 28641 28577 28675 28611
rect 30849 28577 30883 28611
rect 10149 28509 10183 28543
rect 10977 28509 11011 28543
rect 14105 28509 14139 28543
rect 14289 28509 14323 28543
rect 15117 28509 15151 28543
rect 15301 28509 15335 28543
rect 15485 28509 15519 28543
rect 18245 28509 18279 28543
rect 19257 28509 19291 28543
rect 21465 28509 21499 28543
rect 21833 28509 21867 28543
rect 22661 28509 22695 28543
rect 22937 28509 22971 28543
rect 24409 28509 24443 28543
rect 24593 28509 24627 28543
rect 24685 28509 24719 28543
rect 24961 28509 24995 28543
rect 25697 28509 25731 28543
rect 27353 28509 27387 28543
rect 27501 28509 27535 28543
rect 27721 28509 27755 28543
rect 27818 28509 27852 28543
rect 28549 28509 28583 28543
rect 29929 28509 29963 28543
rect 30573 28509 30607 28543
rect 31585 28509 31619 28543
rect 31677 28509 31711 28543
rect 32321 28509 32355 28543
rect 32505 28509 32539 28543
rect 34713 28509 34747 28543
rect 35449 28509 35483 28543
rect 47685 28509 47719 28543
rect 14933 28441 14967 28475
rect 16313 28441 16347 28475
rect 21649 28441 21683 28475
rect 21741 28441 21775 28475
rect 25145 28441 25179 28475
rect 27629 28441 27663 28475
rect 29745 28441 29779 28475
rect 33425 28441 33459 28475
rect 15209 28373 15243 28407
rect 17785 28373 17819 28407
rect 18337 28373 18371 28407
rect 21005 28373 21039 28407
rect 22017 28373 22051 28407
rect 22477 28373 22511 28407
rect 22845 28373 22879 28407
rect 31861 28373 31895 28407
rect 14657 28169 14691 28203
rect 16957 28169 16991 28203
rect 20545 28169 20579 28203
rect 21189 28169 21223 28203
rect 22201 28169 22235 28203
rect 24869 28169 24903 28203
rect 25605 28169 25639 28203
rect 26341 28169 26375 28203
rect 27169 28169 27203 28203
rect 27905 28169 27939 28203
rect 11805 28101 11839 28135
rect 14933 28101 14967 28135
rect 17049 28101 17083 28135
rect 18245 28101 18279 28135
rect 21833 28101 21867 28135
rect 29193 28101 29227 28135
rect 30389 28101 30423 28135
rect 35265 28101 35299 28135
rect 9137 28033 9171 28067
rect 11529 28033 11563 28067
rect 13553 28033 13587 28067
rect 14565 28033 14599 28067
rect 14749 28033 14783 28067
rect 15577 28033 15611 28067
rect 15761 28033 15795 28067
rect 15853 28033 15887 28067
rect 17141 28033 17175 28067
rect 18061 28033 18095 28067
rect 20453 28033 20487 28067
rect 21097 28033 21131 28067
rect 21281 28033 21315 28067
rect 22063 28033 22097 28067
rect 22293 28033 22327 28067
rect 22937 28033 22971 28067
rect 24685 28033 24719 28067
rect 25513 28033 25547 28067
rect 26249 28033 26283 28067
rect 26433 28033 26467 28067
rect 27077 28033 27111 28067
rect 27721 28033 27755 28067
rect 28457 28033 28491 28067
rect 29101 28033 29135 28067
rect 31217 28033 31251 28067
rect 31401 28033 31435 28067
rect 31493 28033 31527 28067
rect 35173 28033 35207 28067
rect 47593 28033 47627 28067
rect 9321 27965 9355 27999
rect 9781 27965 9815 27999
rect 15393 27965 15427 27999
rect 16681 27965 16715 27999
rect 19901 27965 19935 27999
rect 28549 27965 28583 27999
rect 32965 27965 32999 27999
rect 33241 27965 33275 27999
rect 34713 27965 34747 27999
rect 14381 27897 14415 27931
rect 30573 27897 30607 27931
rect 13645 27829 13679 27863
rect 23121 27829 23155 27863
rect 31033 27829 31067 27863
rect 47685 27829 47719 27863
rect 21557 27625 21591 27659
rect 23213 27625 23247 27659
rect 9689 27557 9723 27591
rect 12081 27557 12115 27591
rect 20545 27557 20579 27591
rect 23581 27557 23615 27591
rect 27077 27557 27111 27591
rect 30757 27557 30791 27591
rect 32137 27557 32171 27591
rect 14565 27489 14599 27523
rect 16681 27489 16715 27523
rect 20821 27489 20855 27523
rect 21465 27489 21499 27523
rect 22753 27489 22787 27523
rect 23305 27489 23339 27523
rect 46305 27489 46339 27523
rect 46489 27489 46523 27523
rect 48145 27489 48179 27523
rect 9597 27421 9631 27455
rect 10885 27421 10919 27455
rect 11069 27421 11103 27455
rect 11989 27421 12023 27455
rect 13369 27421 13403 27455
rect 14105 27421 14139 27455
rect 16405 27421 16439 27455
rect 17877 27421 17911 27455
rect 20453 27421 20487 27455
rect 20729 27421 20763 27455
rect 21649 27421 21683 27455
rect 22385 27421 22419 27455
rect 23213 27421 23247 27455
rect 24869 27421 24903 27455
rect 26157 27421 26191 27455
rect 27905 27421 27939 27455
rect 28089 27421 28123 27455
rect 29561 27421 29595 27455
rect 29745 27421 29779 27455
rect 30113 27421 30147 27455
rect 30573 27421 30607 27455
rect 31493 27421 31527 27455
rect 31641 27421 31675 27455
rect 31958 27421 31992 27455
rect 13461 27353 13495 27387
rect 14289 27353 14323 27387
rect 21373 27353 21407 27387
rect 22569 27353 22603 27387
rect 25053 27353 25087 27387
rect 26893 27353 26927 27387
rect 27721 27353 27755 27387
rect 28181 27353 28215 27387
rect 28733 27353 28767 27387
rect 28917 27353 28951 27387
rect 31769 27353 31803 27387
rect 31861 27353 31895 27387
rect 10977 27285 11011 27319
rect 17969 27285 18003 27319
rect 20913 27285 20947 27319
rect 21833 27285 21867 27319
rect 26249 27285 26283 27319
rect 30021 27285 30055 27319
rect 15301 27081 15335 27115
rect 17233 27081 17267 27115
rect 27829 27081 27863 27115
rect 28641 27081 28675 27115
rect 29285 27081 29319 27115
rect 30849 27081 30883 27115
rect 18061 27013 18095 27047
rect 27629 27013 27663 27047
rect 10701 26945 10735 26979
rect 11621 26945 11655 26979
rect 13921 26945 13955 26979
rect 15117 26945 15151 26979
rect 15393 26945 15427 26979
rect 15853 26945 15887 26979
rect 17141 26945 17175 26979
rect 17877 26945 17911 26979
rect 20729 26945 20763 26979
rect 21833 26945 21867 26979
rect 22017 26945 22051 26979
rect 22109 26945 22143 26979
rect 22385 26945 22419 26979
rect 24041 26945 24075 26979
rect 24317 26945 24351 26979
rect 25697 26945 25731 26979
rect 28549 26945 28583 26979
rect 29193 26945 29227 26979
rect 30846 26945 30880 26979
rect 32321 26945 32355 26979
rect 32413 26945 32447 26979
rect 32597 26945 32631 26979
rect 32689 26945 32723 26979
rect 33425 26945 33459 26979
rect 33609 26945 33643 26979
rect 33977 26945 34011 26979
rect 19717 26877 19751 26911
rect 22201 26877 22235 26911
rect 31309 26877 31343 26911
rect 33701 26877 33735 26911
rect 33793 26877 33827 26911
rect 24133 26809 24167 26843
rect 24225 26809 24259 26843
rect 10701 26741 10735 26775
rect 11713 26741 11747 26775
rect 14105 26741 14139 26775
rect 15117 26741 15151 26775
rect 15853 26741 15887 26775
rect 20821 26741 20855 26775
rect 22569 26741 22603 26775
rect 23857 26741 23891 26775
rect 25881 26741 25915 26775
rect 27813 26741 27847 26775
rect 27997 26741 28031 26775
rect 30665 26741 30699 26775
rect 31217 26741 31251 26775
rect 32137 26741 32171 26775
rect 34161 26741 34195 26775
rect 47777 26741 47811 26775
rect 12357 26537 12391 26571
rect 14565 26537 14599 26571
rect 16865 26537 16899 26571
rect 19796 26537 19830 26571
rect 24777 26537 24811 26571
rect 27077 26537 27111 26571
rect 27261 26537 27295 26571
rect 28273 26537 28307 26571
rect 28733 26537 28767 26571
rect 32413 26537 32447 26571
rect 30113 26469 30147 26503
rect 10609 26401 10643 26435
rect 10885 26401 10919 26435
rect 15117 26401 15151 26435
rect 19533 26401 19567 26435
rect 21281 26401 21315 26435
rect 21833 26401 21867 26435
rect 23857 26401 23891 26435
rect 30665 26401 30699 26435
rect 33701 26401 33735 26435
rect 46305 26401 46339 26435
rect 14197 26333 14231 26367
rect 14381 26333 14415 26367
rect 21741 26333 21775 26367
rect 23489 26333 23523 26367
rect 24685 26333 24719 26367
rect 24869 26333 24903 26367
rect 26709 26333 26743 26367
rect 27077 26333 27111 26367
rect 28181 26333 28215 26367
rect 28457 26333 28491 26367
rect 29837 26333 29871 26367
rect 29929 26333 29963 26367
rect 30187 26333 30221 26367
rect 33333 26333 33367 26367
rect 33517 26333 33551 26367
rect 33609 26333 33643 26367
rect 33885 26333 33919 26367
rect 15393 26265 15427 26299
rect 23673 26265 23707 26299
rect 24409 26265 24443 26299
rect 29653 26265 29687 26299
rect 30941 26265 30975 26299
rect 46489 26265 46523 26299
rect 48145 26265 48179 26299
rect 25053 26197 25087 26231
rect 34069 26197 34103 26231
rect 13277 25993 13311 26027
rect 15117 25993 15151 26027
rect 15301 25993 15335 26027
rect 16037 25993 16071 26027
rect 17417 25993 17451 26027
rect 23857 25993 23891 26027
rect 28825 25993 28859 26027
rect 30481 25993 30515 26027
rect 31309 25993 31343 26027
rect 32597 25993 32631 26027
rect 35633 25993 35667 26027
rect 46121 25993 46155 26027
rect 11713 25925 11747 25959
rect 12909 25925 12943 25959
rect 13125 25925 13159 25959
rect 14933 25925 14967 25959
rect 18061 25925 18095 25959
rect 30941 25925 30975 25959
rect 34161 25925 34195 25959
rect 9965 25857 9999 25891
rect 11529 25857 11563 25891
rect 11805 25857 11839 25891
rect 14197 25857 14231 25891
rect 15209 25857 15243 25891
rect 15945 25857 15979 25891
rect 17233 25857 17267 25891
rect 18245 25857 18279 25891
rect 20821 25857 20855 25891
rect 21005 25857 21039 25891
rect 21281 25857 21315 25891
rect 22937 25857 22971 25891
rect 23765 25857 23799 25891
rect 24593 25857 24627 25891
rect 24685 25857 24719 25891
rect 26985 25857 27019 25891
rect 28641 25857 28675 25891
rect 30297 25857 30331 25891
rect 31125 25857 31159 25891
rect 32505 25857 32539 25891
rect 46305 25857 46339 25891
rect 46765 25857 46799 25891
rect 15485 25789 15519 25823
rect 20913 25789 20947 25823
rect 24041 25789 24075 25823
rect 24869 25789 24903 25823
rect 30113 25789 30147 25823
rect 33885 25789 33919 25823
rect 11529 25721 11563 25755
rect 21097 25721 21131 25755
rect 23397 25721 23431 25755
rect 47777 25721 47811 25755
rect 10057 25653 10091 25687
rect 13093 25653 13127 25687
rect 14381 25653 14415 25687
rect 20545 25653 20579 25687
rect 22753 25653 22787 25687
rect 24777 25653 24811 25687
rect 27169 25653 27203 25687
rect 46857 25653 46891 25687
rect 14289 25449 14323 25483
rect 15117 25449 15151 25483
rect 15669 25449 15703 25483
rect 28825 25449 28859 25483
rect 31585 25449 31619 25483
rect 12081 25381 12115 25415
rect 23857 25381 23891 25415
rect 24409 25381 24443 25415
rect 26709 25381 26743 25415
rect 34069 25381 34103 25415
rect 9689 25313 9723 25347
rect 22385 25313 22419 25347
rect 27169 25313 27203 25347
rect 27353 25313 27387 25347
rect 30941 25313 30975 25347
rect 31493 25313 31527 25347
rect 34713 25313 34747 25347
rect 46489 25313 46523 25347
rect 48145 25313 48179 25347
rect 1869 25245 1903 25279
rect 11897 25245 11931 25279
rect 12633 25245 12667 25279
rect 13369 25245 13403 25279
rect 14933 25245 14967 25279
rect 15669 25245 15703 25279
rect 15853 25245 15887 25279
rect 16497 25245 16531 25279
rect 17693 25245 17727 25279
rect 22109 25245 22143 25279
rect 24593 25245 24627 25279
rect 24685 25245 24719 25279
rect 25605 25245 25639 25279
rect 25881 25245 25915 25279
rect 27077 25245 27111 25279
rect 28641 25245 28675 25279
rect 29829 25223 29863 25257
rect 29929 25245 29963 25279
rect 30072 25245 30106 25279
rect 30195 25245 30229 25279
rect 31677 25245 31711 25279
rect 33977 25245 34011 25279
rect 45477 25245 45511 25279
rect 46305 25245 46339 25279
rect 9965 25177 9999 25211
rect 12725 25177 12759 25211
rect 14105 25177 14139 25211
rect 14321 25177 14355 25211
rect 24409 25177 24443 25211
rect 30757 25177 30791 25211
rect 31401 25177 31435 25211
rect 34989 25177 35023 25211
rect 1961 25109 1995 25143
rect 11437 25109 11471 25143
rect 13461 25109 13495 25143
rect 14473 25109 14507 25143
rect 16681 25109 16715 25143
rect 17785 25109 17819 25143
rect 25421 25109 25455 25143
rect 25789 25109 25823 25143
rect 29653 25109 29687 25143
rect 31861 25109 31895 25143
rect 36461 25109 36495 25143
rect 45569 25109 45603 25143
rect 24869 24905 24903 24939
rect 11529 24837 11563 24871
rect 11729 24837 11763 24871
rect 13645 24837 13679 24871
rect 21281 24837 21315 24871
rect 26065 24837 26099 24871
rect 26157 24837 26191 24871
rect 29469 24837 29503 24871
rect 31217 24837 31251 24871
rect 35725 24837 35759 24871
rect 12449 24769 12483 24803
rect 23029 24769 23063 24803
rect 23121 24769 23155 24803
rect 24685 24769 24719 24803
rect 24961 24769 24995 24803
rect 25881 24769 25915 24803
rect 26249 24769 26283 24803
rect 26985 24769 27019 24803
rect 27997 24769 28031 24803
rect 28181 24769 28215 24803
rect 29285 24769 29319 24803
rect 30297 24769 30331 24803
rect 31033 24769 31067 24803
rect 34713 24769 34747 24803
rect 34805 24769 34839 24803
rect 36093 24769 36127 24803
rect 43453 24769 43487 24803
rect 43637 24769 43671 24803
rect 44649 24769 44683 24803
rect 45293 24769 45327 24803
rect 47593 24769 47627 24803
rect 8401 24701 8435 24735
rect 8585 24701 8619 24735
rect 8861 24701 8895 24735
rect 13461 24701 13495 24735
rect 14565 24701 14599 24735
rect 17233 24701 17267 24735
rect 17509 24701 17543 24735
rect 18981 24701 19015 24735
rect 19441 24701 19475 24735
rect 19625 24701 19659 24735
rect 28457 24701 28491 24735
rect 30573 24701 30607 24735
rect 40049 24701 40083 24735
rect 40233 24701 40267 24735
rect 40509 24701 40543 24735
rect 47685 24701 47719 24735
rect 11897 24633 11931 24667
rect 27169 24633 27203 24667
rect 11713 24565 11747 24599
rect 12541 24565 12575 24599
rect 24501 24565 24535 24599
rect 26433 24565 26467 24599
rect 28365 24565 28399 24599
rect 30113 24565 30147 24599
rect 30481 24565 30515 24599
rect 31401 24565 31435 24599
rect 36369 24565 36403 24599
rect 43545 24565 43579 24599
rect 44741 24565 44775 24599
rect 46581 24565 46615 24599
rect 10333 24361 10367 24395
rect 12541 24361 12575 24395
rect 17049 24361 17083 24395
rect 18521 24361 18555 24395
rect 19441 24361 19475 24395
rect 28181 24361 28215 24395
rect 28641 24361 28675 24395
rect 30205 24361 30239 24395
rect 33241 24361 33275 24395
rect 12725 24293 12759 24327
rect 18705 24293 18739 24327
rect 27261 24293 27295 24327
rect 41521 24293 41555 24327
rect 10885 24225 10919 24259
rect 10977 24225 11011 24259
rect 14841 24225 14875 24259
rect 15117 24225 15151 24259
rect 19993 24225 20027 24259
rect 26985 24225 27019 24259
rect 29653 24225 29687 24259
rect 31769 24225 31803 24259
rect 37105 24225 37139 24259
rect 41061 24225 41095 24259
rect 46397 24225 46431 24259
rect 46673 24225 46707 24259
rect 10514 24157 10548 24191
rect 11621 24157 11655 24191
rect 11897 24157 11931 24191
rect 13185 24157 13219 24191
rect 14749 24157 14783 24191
rect 15761 24157 15795 24191
rect 16957 24157 16991 24191
rect 17785 24157 17819 24191
rect 17877 24157 17911 24191
rect 19349 24157 19383 24191
rect 23397 24157 23431 24191
rect 25973 24157 26007 24191
rect 26157 24157 26191 24191
rect 26249 24157 26283 24191
rect 26893 24157 26927 24191
rect 28181 24157 28215 24191
rect 28365 24157 28399 24191
rect 28457 24157 28491 24191
rect 29561 24157 29595 24191
rect 29745 24157 29779 24191
rect 30205 24157 30239 24191
rect 30481 24157 30515 24191
rect 31493 24157 31527 24191
rect 35541 24157 35575 24191
rect 36369 24157 36403 24191
rect 40233 24157 40267 24191
rect 40325 24157 40359 24191
rect 41231 24157 41265 24191
rect 43361 24157 43395 24191
rect 43545 24157 43579 24191
rect 44005 24157 44039 24191
rect 45293 24157 45327 24191
rect 46213 24157 46247 24191
rect 12357 24089 12391 24123
rect 12573 24089 12607 24123
rect 17601 24089 17635 24123
rect 18337 24089 18371 24123
rect 20177 24089 20211 24123
rect 21833 24089 21867 24123
rect 30389 24089 30423 24123
rect 44281 24089 44315 24123
rect 45569 24089 45603 24123
rect 10517 24021 10551 24055
rect 11437 24021 11471 24055
rect 11805 24021 11839 24055
rect 13369 24021 13403 24055
rect 15761 24021 15795 24055
rect 17699 24021 17733 24055
rect 18547 24021 18581 24055
rect 23489 24021 23523 24055
rect 25789 24021 25823 24055
rect 35633 24021 35667 24055
rect 43453 24021 43487 24055
rect 8769 23817 8803 23851
rect 18061 23817 18095 23851
rect 18981 23817 19015 23851
rect 19073 23817 19107 23851
rect 20085 23817 20119 23851
rect 30757 23817 30791 23851
rect 31401 23817 31435 23851
rect 32873 23817 32907 23851
rect 33609 23817 33643 23851
rect 40969 23817 41003 23851
rect 42533 23817 42567 23851
rect 43177 23817 43211 23851
rect 11529 23749 11563 23783
rect 18705 23749 18739 23783
rect 23029 23749 23063 23783
rect 27997 23749 28031 23783
rect 36277 23749 36311 23783
rect 38117 23749 38151 23783
rect 47777 23749 47811 23783
rect 1409 23681 1443 23715
rect 8677 23681 8711 23715
rect 10977 23681 11011 23715
rect 13645 23681 13679 23715
rect 16681 23681 16715 23715
rect 17969 23681 18003 23715
rect 18153 23681 18187 23715
rect 18889 23681 18923 23715
rect 19993 23681 20027 23715
rect 21925 23681 21959 23715
rect 22753 23681 22787 23715
rect 28181 23681 28215 23715
rect 29745 23681 29779 23715
rect 29929 23681 29963 23715
rect 30389 23681 30423 23715
rect 30573 23681 30607 23715
rect 31217 23681 31251 23715
rect 31493 23681 31527 23715
rect 32781 23681 32815 23715
rect 33425 23681 33459 23715
rect 35541 23681 35575 23715
rect 37289 23681 37323 23715
rect 40601 23681 40635 23715
rect 42993 23681 43027 23715
rect 43729 23681 43763 23715
rect 43913 23681 43947 23715
rect 44741 23681 44775 23715
rect 45201 23681 45235 23715
rect 47593 23681 47627 23715
rect 11989 23613 12023 23647
rect 13829 23613 13863 23647
rect 14105 23613 14139 23647
rect 24501 23613 24535 23647
rect 28365 23613 28399 23647
rect 29837 23613 29871 23647
rect 40693 23613 40727 23647
rect 42901 23613 42935 23647
rect 45385 23613 45419 23647
rect 45661 23613 45695 23647
rect 1593 23545 1627 23579
rect 11805 23545 11839 23579
rect 10793 23477 10827 23511
rect 16773 23477 16807 23511
rect 19257 23477 19291 23511
rect 22017 23477 22051 23511
rect 31217 23477 31251 23511
rect 47961 23477 47995 23511
rect 13185 23273 13219 23307
rect 14197 23273 14231 23307
rect 16865 23273 16899 23307
rect 26985 23273 27019 23307
rect 33885 23273 33919 23307
rect 43729 23273 43763 23307
rect 44281 23273 44315 23307
rect 28181 23205 28215 23239
rect 11713 23137 11747 23171
rect 25513 23137 25547 23171
rect 32137 23137 32171 23171
rect 36185 23137 36219 23171
rect 37841 23137 37875 23171
rect 40877 23137 40911 23171
rect 42073 23137 42107 23171
rect 46305 23137 46339 23171
rect 48145 23137 48179 23171
rect 11437 23069 11471 23103
rect 14105 23069 14139 23103
rect 15117 23069 15151 23103
rect 17417 23069 17451 23103
rect 19441 23069 19475 23103
rect 19625 23069 19659 23103
rect 20913 23069 20947 23103
rect 25237 23069 25271 23103
rect 28181 23069 28215 23103
rect 28457 23069 28491 23103
rect 30389 23069 30423 23103
rect 30665 23069 30699 23103
rect 30757 23069 30791 23103
rect 31677 23069 31711 23103
rect 36001 23069 36035 23103
rect 40417 23069 40451 23103
rect 43361 23069 43395 23103
rect 44465 23069 44499 23103
rect 45201 23069 45235 23103
rect 15393 23001 15427 23035
rect 21189 23001 21223 23035
rect 30573 23001 30607 23035
rect 32413 23001 32447 23035
rect 41061 23001 41095 23035
rect 43545 23001 43579 23035
rect 45569 23001 45603 23035
rect 46489 23001 46523 23035
rect 17509 22933 17543 22967
rect 19809 22933 19843 22967
rect 22661 22933 22695 22967
rect 28365 22933 28399 22967
rect 30941 22933 30975 22967
rect 31493 22933 31527 22967
rect 40233 22933 40267 22967
rect 12449 22729 12483 22763
rect 18429 22729 18463 22763
rect 19165 22729 19199 22763
rect 21189 22729 21223 22763
rect 27077 22729 27111 22763
rect 28273 22729 28307 22763
rect 31585 22729 31619 22763
rect 33333 22729 33367 22763
rect 40785 22729 40819 22763
rect 46949 22729 46983 22763
rect 48145 22729 48179 22763
rect 29101 22661 29135 22695
rect 29193 22661 29227 22695
rect 31217 22661 31251 22695
rect 31401 22661 31435 22695
rect 45477 22661 45511 22695
rect 46305 22661 46339 22695
rect 8953 22593 8987 22627
rect 9781 22593 9815 22627
rect 10609 22593 10643 22627
rect 11529 22593 11563 22627
rect 12357 22593 12391 22627
rect 13921 22593 13955 22627
rect 18981 22593 19015 22627
rect 19257 22593 19291 22627
rect 20453 22593 20487 22627
rect 21097 22593 21131 22627
rect 21925 22593 21959 22627
rect 26985 22593 27019 22627
rect 28089 22593 28123 22627
rect 28273 22593 28307 22627
rect 28917 22593 28951 22627
rect 29285 22593 29319 22627
rect 30205 22593 30239 22627
rect 33241 22593 33275 22627
rect 36093 22593 36127 22627
rect 40325 22593 40359 22627
rect 44833 22593 44867 22627
rect 45017 22593 45051 22627
rect 46857 22593 46891 22627
rect 47593 22593 47627 22627
rect 9873 22525 9907 22559
rect 16681 22525 16715 22559
rect 16957 22525 16991 22559
rect 22937 22525 22971 22559
rect 23121 22525 23155 22559
rect 23489 22525 23523 22559
rect 29929 22525 29963 22559
rect 36645 22525 36679 22559
rect 43361 22525 43395 22559
rect 47869 22525 47903 22559
rect 43637 22457 43671 22491
rect 9045 22389 9079 22423
rect 10149 22389 10183 22423
rect 10701 22389 10735 22423
rect 11621 22389 11655 22423
rect 14105 22389 14139 22423
rect 18981 22389 19015 22423
rect 20545 22389 20579 22423
rect 22017 22389 22051 22423
rect 29469 22389 29503 22423
rect 40049 22389 40083 22423
rect 40509 22389 40543 22423
rect 43821 22389 43855 22423
rect 44925 22389 44959 22423
rect 47685 22389 47719 22423
rect 10314 22185 10348 22219
rect 17969 22185 18003 22219
rect 23213 22185 23247 22219
rect 25408 22185 25442 22219
rect 10057 22049 10091 22083
rect 11805 22049 11839 22083
rect 14105 22049 14139 22083
rect 17693 22049 17727 22083
rect 21005 22049 21039 22083
rect 26893 22049 26927 22083
rect 29009 22049 29043 22083
rect 42809 22049 42843 22083
rect 43913 22049 43947 22083
rect 47593 22049 47627 22083
rect 8953 21981 8987 22015
rect 12357 21981 12391 22015
rect 13369 21981 13403 22015
rect 16405 21981 16439 22015
rect 17601 21981 17635 22015
rect 18429 21981 18463 22015
rect 18613 21981 18647 22015
rect 20821 21981 20855 22015
rect 23121 21981 23155 22015
rect 25145 21981 25179 22015
rect 27353 21981 27387 22015
rect 28181 21981 28215 22015
rect 28825 21981 28859 22015
rect 34897 21981 34931 22015
rect 40325 21981 40359 22015
rect 40509 21981 40543 22015
rect 42717 21981 42751 22015
rect 42901 21981 42935 22015
rect 43361 21981 43395 22015
rect 43545 21981 43579 22015
rect 45569 21981 45603 22015
rect 46029 21981 46063 22015
rect 46305 21981 46339 22015
rect 47317 21981 47351 22015
rect 14289 21913 14323 21947
rect 15945 21913 15979 21947
rect 22661 21913 22695 21947
rect 27445 21913 27479 21947
rect 28641 21913 28675 21947
rect 40601 21913 40635 21947
rect 9045 21845 9079 21879
rect 12541 21845 12575 21879
rect 13461 21845 13495 21879
rect 16589 21845 16623 21879
rect 18521 21845 18555 21879
rect 27997 21845 28031 21879
rect 34713 21845 34747 21879
rect 43545 21845 43579 21879
rect 45385 21845 45419 21879
rect 33333 21641 33367 21675
rect 34161 21641 34195 21675
rect 43085 21641 43119 21675
rect 47777 21641 47811 21675
rect 47961 21641 47995 21675
rect 8769 21573 8803 21607
rect 13645 21573 13679 21607
rect 14381 21573 14415 21607
rect 18153 21573 18187 21607
rect 22017 21573 22051 21607
rect 27721 21573 27755 21607
rect 34805 21573 34839 21607
rect 47869 21573 47903 21607
rect 11529 21505 11563 21539
rect 13553 21505 13587 21539
rect 16037 21505 16071 21539
rect 16865 21505 16899 21539
rect 20821 21505 20855 21539
rect 21833 21505 21867 21539
rect 27445 21505 27479 21539
rect 32321 21505 32355 21539
rect 33701 21505 33735 21539
rect 42901 21505 42935 21539
rect 43085 21505 43119 21539
rect 43729 21505 43763 21539
rect 44741 21505 44775 21539
rect 47593 21505 47627 21539
rect 8585 21437 8619 21471
rect 9045 21437 9079 21471
rect 14197 21437 14231 21471
rect 17877 21437 17911 21471
rect 19625 21437 19659 21471
rect 22293 21437 22327 21471
rect 29193 21437 29227 21471
rect 34713 21437 34747 21471
rect 43821 21437 43855 21471
rect 45201 21437 45235 21471
rect 45385 21437 45419 21471
rect 46857 21437 46891 21471
rect 11529 21369 11563 21403
rect 16681 21369 16715 21403
rect 35265 21369 35299 21403
rect 44097 21369 44131 21403
rect 44557 21369 44591 21403
rect 20913 21301 20947 21335
rect 32137 21301 32171 21335
rect 33793 21301 33827 21335
rect 48145 21301 48179 21335
rect 17233 21097 17267 21131
rect 19349 21097 19383 21131
rect 23857 21097 23891 21131
rect 26893 21097 26927 21131
rect 27813 21097 27847 21131
rect 30205 20961 30239 20995
rect 31217 20961 31251 20995
rect 31769 20961 31803 20995
rect 32137 20961 32171 20995
rect 35265 20961 35299 20995
rect 43085 20961 43119 20995
rect 45201 20961 45235 20995
rect 46305 20961 46339 20995
rect 48145 20961 48179 20995
rect 8953 20893 8987 20927
rect 17141 20893 17175 20927
rect 19257 20893 19291 20927
rect 21373 20893 21407 20927
rect 21649 20893 21683 20927
rect 22109 20893 22143 20927
rect 26709 20893 26743 20927
rect 27721 20893 27755 20927
rect 35909 20893 35943 20927
rect 43269 20893 43303 20927
rect 43453 20893 43487 20927
rect 43913 20893 43947 20927
rect 44097 20893 44131 20927
rect 45661 20893 45695 20927
rect 9137 20825 9171 20859
rect 10793 20825 10827 20859
rect 22385 20825 22419 20859
rect 30297 20825 30331 20859
rect 31861 20825 31895 20859
rect 35357 20825 35391 20859
rect 45753 20825 45787 20859
rect 46489 20825 46523 20859
rect 44005 20757 44039 20791
rect 13277 20553 13311 20587
rect 13921 20553 13955 20587
rect 14289 20553 14323 20587
rect 20101 20553 20135 20587
rect 21097 20553 21131 20587
rect 23305 20553 23339 20587
rect 32597 20553 32631 20587
rect 42533 20553 42567 20587
rect 44189 20553 44223 20587
rect 48053 20553 48087 20587
rect 13737 20485 13771 20519
rect 19901 20485 19935 20519
rect 20913 20485 20947 20519
rect 28365 20485 28399 20519
rect 29101 20485 29135 20519
rect 10885 20417 10919 20451
rect 14013 20417 14047 20451
rect 14105 20417 14139 20451
rect 15117 20417 15151 20451
rect 15945 20417 15979 20451
rect 17049 20417 17083 20451
rect 18061 20417 18095 20451
rect 21005 20417 21039 20451
rect 22385 20417 22419 20451
rect 23213 20417 23247 20451
rect 24869 20417 24903 20451
rect 25789 20417 25823 20451
rect 26249 20417 26283 20451
rect 26985 20417 27019 20451
rect 28273 20417 28307 20451
rect 31217 20417 31251 20451
rect 32137 20417 32171 20451
rect 42441 20417 42475 20451
rect 42625 20417 42659 20451
rect 43453 20417 43487 20451
rect 44649 20417 44683 20451
rect 47593 20417 47627 20451
rect 10977 20349 11011 20383
rect 11529 20349 11563 20383
rect 11805 20349 11839 20383
rect 21281 20349 21315 20383
rect 22293 20349 22327 20383
rect 22753 20349 22787 20383
rect 28917 20349 28951 20383
rect 30021 20349 30055 20383
rect 43545 20349 43579 20383
rect 44833 20349 44867 20383
rect 46029 20349 46063 20383
rect 17233 20281 17267 20315
rect 20729 20281 20763 20315
rect 15301 20213 15335 20247
rect 16037 20213 16071 20247
rect 18153 20213 18187 20247
rect 20085 20213 20119 20247
rect 20269 20213 20303 20247
rect 25053 20213 25087 20247
rect 25605 20213 25639 20247
rect 26341 20213 26375 20247
rect 27077 20213 27111 20247
rect 31309 20213 31343 20247
rect 32321 20213 32355 20247
rect 47685 20213 47719 20247
rect 45201 20009 45235 20043
rect 11529 19941 11563 19975
rect 12817 19941 12851 19975
rect 21741 19941 21775 19975
rect 43821 19941 43855 19975
rect 16865 19873 16899 19907
rect 17141 19873 17175 19907
rect 25237 19873 25271 19907
rect 25513 19873 25547 19907
rect 30205 19873 30239 19907
rect 31677 19873 31711 19907
rect 43361 19873 43395 19907
rect 43913 19873 43947 19907
rect 46213 19873 46247 19907
rect 46397 19873 46431 19907
rect 46949 19873 46983 19907
rect 11713 19805 11747 19839
rect 11989 19805 12023 19839
rect 12173 19805 12207 19839
rect 12725 19805 12759 19839
rect 13369 19805 13403 19839
rect 13461 19805 13495 19839
rect 14473 19805 14507 19839
rect 19993 19805 20027 19839
rect 24501 19805 24535 19839
rect 30021 19805 30055 19839
rect 43085 19805 43119 19839
rect 43637 19805 43671 19839
rect 45109 19805 45143 19839
rect 14749 19737 14783 19771
rect 20269 19737 20303 19771
rect 24777 19737 24811 19771
rect 16221 19669 16255 19703
rect 18613 19669 18647 19703
rect 26985 19669 27019 19703
rect 23949 19465 23983 19499
rect 27997 19465 28031 19499
rect 28917 19465 28951 19499
rect 29929 19465 29963 19499
rect 43545 19465 43579 19499
rect 47777 19465 47811 19499
rect 48145 19465 48179 19499
rect 2237 19397 2271 19431
rect 13829 19397 13863 19431
rect 14013 19397 14047 19431
rect 14105 19397 14139 19431
rect 14841 19397 14875 19431
rect 15041 19397 15075 19431
rect 15761 19397 15795 19431
rect 17049 19397 17083 19431
rect 19533 19397 19567 19431
rect 21925 19397 21959 19431
rect 47869 19397 47903 19431
rect 11897 19329 11931 19363
rect 13001 19329 13035 19363
rect 14197 19329 14231 19363
rect 15669 19329 15703 19363
rect 16773 19329 16807 19363
rect 17969 19329 18003 19363
rect 19441 19329 19475 19363
rect 20177 19329 20211 19363
rect 21005 19329 21039 19363
rect 21189 19329 21223 19363
rect 21281 19329 21315 19363
rect 21833 19329 21867 19363
rect 22477 19329 22511 19363
rect 23765 19329 23799 19363
rect 24593 19329 24627 19363
rect 25427 19329 25461 19363
rect 25605 19329 25639 19363
rect 28273 19329 28307 19363
rect 28457 19329 28491 19363
rect 29285 19329 29319 19363
rect 29469 19329 29503 19363
rect 30113 19329 30147 19363
rect 43361 19329 43395 19363
rect 43545 19329 43579 19363
rect 45937 19329 45971 19363
rect 46489 19329 46523 19363
rect 46673 19329 46707 19363
rect 46857 19329 46891 19363
rect 47961 19329 47995 19363
rect 2053 19261 2087 19295
rect 2789 19261 2823 19295
rect 13093 19261 13127 19295
rect 18061 19261 18095 19295
rect 18337 19261 18371 19295
rect 20269 19261 20303 19295
rect 20545 19261 20579 19295
rect 23581 19261 23615 19295
rect 24685 19261 24719 19295
rect 28641 19261 28675 19295
rect 29101 19261 29135 19295
rect 15209 19193 15243 19227
rect 47593 19193 47627 19227
rect 11897 19125 11931 19159
rect 13369 19125 13403 19159
rect 14381 19125 14415 19159
rect 15025 19125 15059 19159
rect 21005 19125 21039 19159
rect 22569 19125 22603 19159
rect 24869 19125 24903 19159
rect 25513 19125 25547 19159
rect 45477 19125 45511 19159
rect 46213 19125 46247 19159
rect 2329 18921 2363 18955
rect 3065 18921 3099 18955
rect 13553 18921 13587 18955
rect 14105 18921 14139 18955
rect 14749 18853 14783 18887
rect 24777 18853 24811 18887
rect 27169 18853 27203 18887
rect 28917 18853 28951 18887
rect 45661 18853 45695 18887
rect 11805 18785 11839 18819
rect 12081 18785 12115 18819
rect 25697 18785 25731 18819
rect 27905 18785 27939 18819
rect 30297 18785 30331 18819
rect 46305 18785 46339 18819
rect 48145 18785 48179 18819
rect 2973 18717 3007 18751
rect 14105 18717 14139 18751
rect 14289 18717 14323 18751
rect 14749 18717 14783 18751
rect 15025 18717 15059 18751
rect 17141 18717 17175 18751
rect 20177 18717 20211 18751
rect 20361 18717 20395 18751
rect 20821 18717 20855 18751
rect 24409 18717 24443 18751
rect 24593 18717 24627 18751
rect 25421 18717 25455 18751
rect 27997 18717 28031 18751
rect 28825 18717 28859 18751
rect 29009 18717 29043 18751
rect 43729 18717 43763 18751
rect 43913 18717 43947 18751
rect 45017 18717 45051 18751
rect 45201 18717 45235 18751
rect 45845 18717 45879 18751
rect 20269 18649 20303 18683
rect 21097 18649 21131 18683
rect 30481 18649 30515 18683
rect 32137 18649 32171 18683
rect 46489 18649 46523 18683
rect 14933 18581 14967 18615
rect 17325 18581 17359 18615
rect 22569 18581 22603 18615
rect 28365 18581 28399 18615
rect 43821 18581 43855 18615
rect 45109 18581 45143 18615
rect 13185 18377 13219 18411
rect 20913 18377 20947 18411
rect 47685 18377 47719 18411
rect 42717 18309 42751 18343
rect 45385 18309 45419 18343
rect 1409 18241 1443 18275
rect 13093 18241 13127 18275
rect 16957 18241 16991 18275
rect 20913 18241 20947 18275
rect 23305 18241 23339 18275
rect 24777 18241 24811 18275
rect 27537 18241 27571 18275
rect 28181 18241 28215 18275
rect 30665 18241 30699 18275
rect 31125 18241 31159 18275
rect 40785 18241 40819 18275
rect 40969 18241 41003 18275
rect 41429 18241 41463 18275
rect 41613 18241 41647 18275
rect 42441 18241 42475 18275
rect 43545 18241 43579 18275
rect 43821 18241 43855 18275
rect 47593 18241 47627 18275
rect 17141 18173 17175 18207
rect 18797 18173 18831 18207
rect 23581 18173 23615 18207
rect 28365 18173 28399 18207
rect 28641 18173 28675 18207
rect 31585 18173 31619 18207
rect 41521 18173 41555 18207
rect 42717 18173 42751 18207
rect 44557 18173 44591 18207
rect 45201 18173 45235 18207
rect 46857 18173 46891 18207
rect 27629 18105 27663 18139
rect 1593 18037 1627 18071
rect 24593 18037 24627 18071
rect 30481 18037 30515 18071
rect 31401 18037 31435 18071
rect 40785 18037 40819 18071
rect 42533 18037 42567 18071
rect 17233 17833 17267 17867
rect 21741 17833 21775 17867
rect 45385 17833 45419 17867
rect 28917 17765 28951 17799
rect 41337 17765 41371 17799
rect 42441 17765 42475 17799
rect 14657 17697 14691 17731
rect 24685 17697 24719 17731
rect 24777 17697 24811 17731
rect 30205 17697 30239 17731
rect 30389 17697 30423 17731
rect 32045 17697 32079 17731
rect 40969 17697 41003 17731
rect 1685 17629 1719 17663
rect 2145 17629 2179 17663
rect 14841 17629 14875 17663
rect 17141 17629 17175 17663
rect 18521 17629 18555 17663
rect 19257 17629 19291 17663
rect 21557 17629 21591 17663
rect 23581 17629 23615 17663
rect 23673 17629 23707 17663
rect 24593 17629 24627 17663
rect 24869 17629 24903 17663
rect 25421 17629 25455 17663
rect 27813 17629 27847 17663
rect 28181 17629 28215 17663
rect 28457 17629 28491 17663
rect 28641 17629 28675 17663
rect 41889 17629 41923 17663
rect 42165 17629 42199 17663
rect 42349 17629 42383 17663
rect 43361 17629 43395 17663
rect 43453 17629 43487 17663
rect 43637 17629 43671 17663
rect 45017 17629 45051 17663
rect 46305 17629 46339 17663
rect 18613 17561 18647 17595
rect 19441 17561 19475 17595
rect 21097 17561 21131 17595
rect 23305 17561 23339 17595
rect 42717 17561 42751 17595
rect 44005 17561 44039 17595
rect 45201 17561 45235 17595
rect 46489 17561 46523 17595
rect 48145 17561 48179 17595
rect 2237 17493 2271 17527
rect 15025 17493 15059 17527
rect 23489 17493 23523 17527
rect 23857 17493 23891 17527
rect 24409 17493 24443 17527
rect 25605 17493 25639 17527
rect 41429 17493 41463 17527
rect 47685 17289 47719 17323
rect 1961 17221 1995 17255
rect 22385 17221 22419 17255
rect 22753 17221 22787 17255
rect 23581 17221 23615 17255
rect 24777 17221 24811 17255
rect 27813 17221 27847 17255
rect 43729 17221 43763 17255
rect 1777 17153 1811 17187
rect 14841 17153 14875 17187
rect 15393 17153 15427 17187
rect 17969 17153 18003 17187
rect 20269 17153 20303 17187
rect 22477 17153 22511 17187
rect 22569 17153 22603 17187
rect 23489 17153 23523 17187
rect 23673 17153 23707 17187
rect 27077 17153 27111 17187
rect 42625 17153 42659 17187
rect 46397 17153 46431 17187
rect 46857 17153 46891 17187
rect 47593 17153 47627 17187
rect 2789 17085 2823 17119
rect 24501 17085 24535 17119
rect 26249 17085 26283 17119
rect 29285 17085 29319 17119
rect 29469 17085 29503 17119
rect 31125 17085 31159 17119
rect 42533 17085 42567 17119
rect 43545 17085 43579 17119
rect 44189 17085 44223 17119
rect 20453 17017 20487 17051
rect 22201 17017 22235 17051
rect 23305 17017 23339 17051
rect 42993 17017 43027 17051
rect 14657 16949 14691 16983
rect 15485 16949 15519 16983
rect 18061 16949 18095 16983
rect 23857 16949 23891 16983
rect 46949 16949 46983 16983
rect 23029 16745 23063 16779
rect 27261 16745 27295 16779
rect 29653 16745 29687 16779
rect 23213 16677 23247 16711
rect 24685 16677 24719 16711
rect 14381 16609 14415 16643
rect 17601 16609 17635 16643
rect 18061 16609 18095 16643
rect 24409 16609 24443 16643
rect 26893 16609 26927 16643
rect 46305 16609 46339 16643
rect 16865 16541 16899 16575
rect 17693 16541 17727 16575
rect 19625 16541 19659 16575
rect 21833 16541 21867 16575
rect 25421 16541 25455 16575
rect 25513 16541 25547 16575
rect 27077 16541 27111 16575
rect 29561 16541 29595 16575
rect 45017 16541 45051 16575
rect 14657 16473 14691 16507
rect 16405 16473 16439 16507
rect 22845 16473 22879 16507
rect 23061 16473 23095 16507
rect 46489 16473 46523 16507
rect 48145 16473 48179 16507
rect 16957 16405 16991 16439
rect 19717 16405 19751 16439
rect 21925 16405 21959 16439
rect 24869 16405 24903 16439
rect 45109 16405 45143 16439
rect 17509 16201 17543 16235
rect 24593 16201 24627 16235
rect 17141 16133 17175 16167
rect 17357 16133 17391 16167
rect 18245 16133 18279 16167
rect 13921 16065 13955 16099
rect 14933 16065 14967 16099
rect 15669 16065 15703 16099
rect 15945 16065 15979 16099
rect 16129 16065 16163 16099
rect 17969 16065 18003 16099
rect 20453 16065 20487 16099
rect 22385 16065 22419 16099
rect 22569 16065 22603 16099
rect 22661 16065 22695 16099
rect 23121 16065 23155 16099
rect 23305 16065 23339 16099
rect 23765 16065 23799 16099
rect 24409 16065 24443 16099
rect 43913 16065 43947 16099
rect 47777 16065 47811 16099
rect 14013 15997 14047 16031
rect 14289 15997 14323 16031
rect 44097 15997 44131 16031
rect 45477 15997 45511 16031
rect 22385 15929 22419 15963
rect 14933 15861 14967 15895
rect 15485 15861 15519 15895
rect 17325 15861 17359 15895
rect 19717 15861 19751 15895
rect 20637 15861 20671 15895
rect 23121 15861 23155 15895
rect 23857 15861 23891 15895
rect 17601 15657 17635 15691
rect 17785 15657 17819 15691
rect 44097 15657 44131 15691
rect 14933 15521 14967 15555
rect 15209 15521 15243 15555
rect 20913 15521 20947 15555
rect 21189 15521 21223 15555
rect 23581 15521 23615 15555
rect 23857 15521 23891 15555
rect 24685 15521 24719 15555
rect 45017 15521 45051 15555
rect 45201 15521 45235 15555
rect 46673 15521 46707 15555
rect 2053 15453 2087 15487
rect 18429 15453 18463 15487
rect 18613 15453 18647 15487
rect 19441 15453 19475 15487
rect 19993 15453 20027 15487
rect 23489 15453 23523 15487
rect 24409 15453 24443 15487
rect 44005 15453 44039 15487
rect 17417 15385 17451 15419
rect 16681 15317 16715 15351
rect 17627 15317 17661 15351
rect 18521 15317 18555 15351
rect 19441 15317 19475 15351
rect 20085 15317 20119 15351
rect 22661 15317 22695 15351
rect 26157 15317 26191 15351
rect 18429 15113 18463 15147
rect 25329 15113 25363 15147
rect 19165 15045 19199 15079
rect 1777 14977 1811 15011
rect 16681 14977 16715 15011
rect 18061 14977 18095 15011
rect 25237 14977 25271 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 18153 14909 18187 14943
rect 18889 14909 18923 14943
rect 22109 14909 22143 14943
rect 22293 14909 22327 14943
rect 23949 14909 23983 14943
rect 16773 14773 16807 14807
rect 20637 14773 20671 14807
rect 2237 14569 2271 14603
rect 20821 14501 20855 14535
rect 15945 14433 15979 14467
rect 16129 14433 16163 14467
rect 16405 14433 16439 14467
rect 23581 14433 23615 14467
rect 2145 14365 2179 14399
rect 20729 14365 20763 14399
rect 21373 14365 21407 14399
rect 22017 14365 22051 14399
rect 22201 14297 22235 14331
rect 21465 14229 21499 14263
rect 18245 13957 18279 13991
rect 18981 13957 19015 13991
rect 22017 13957 22051 13991
rect 16773 13889 16807 13923
rect 17417 13889 17451 13923
rect 18153 13889 18187 13923
rect 18797 13889 18831 13923
rect 21833 13889 21867 13923
rect 46765 13889 46799 13923
rect 20637 13821 20671 13855
rect 22845 13821 22879 13855
rect 16865 13685 16899 13719
rect 17509 13685 17543 13719
rect 46857 13685 46891 13719
rect 22477 13481 22511 13515
rect 16773 13345 16807 13379
rect 17049 13345 17083 13379
rect 46489 13345 46523 13379
rect 16589 13277 16623 13311
rect 22385 13277 22419 13311
rect 46305 13277 46339 13311
rect 48145 13209 48179 13243
rect 16957 12869 16991 12903
rect 1409 12801 1443 12835
rect 16773 12801 16807 12835
rect 47777 12801 47811 12835
rect 18613 12733 18647 12767
rect 1593 12597 1627 12631
rect 47777 11509 47811 11543
rect 46305 11169 46339 11203
rect 46489 11033 46523 11067
rect 48145 11033 48179 11067
rect 46857 10761 46891 10795
rect 46765 10625 46799 10659
rect 47593 10625 47627 10659
rect 46305 10421 46339 10455
rect 47685 10421 47719 10455
rect 46305 10081 46339 10115
rect 46489 10081 46523 10115
rect 48145 10081 48179 10115
rect 47869 9537 47903 9571
rect 48053 9401 48087 9435
rect 47777 8857 47811 8891
rect 47869 8789 47903 8823
rect 44925 8449 44959 8483
rect 46029 8449 46063 8483
rect 44557 8381 44591 8415
rect 45385 8381 45419 8415
rect 45017 8245 45051 8279
rect 45845 8245 45879 8279
rect 45569 7905 45603 7939
rect 47593 7905 47627 7939
rect 47317 7837 47351 7871
rect 45293 7769 45327 7803
rect 45385 7769 45419 7803
rect 45753 7429 45787 7463
rect 46673 7429 46707 7463
rect 48145 7361 48179 7395
rect 45661 7293 45695 7327
rect 47961 7225 47995 7259
rect 48053 6409 48087 6443
rect 47961 6273 47995 6307
rect 40141 5661 40175 5695
rect 40233 5525 40267 5559
rect 39681 5321 39715 5355
rect 43821 5321 43855 5355
rect 37473 5253 37507 5287
rect 42625 5253 42659 5287
rect 18337 5185 18371 5219
rect 21833 5185 21867 5219
rect 22477 5185 22511 5219
rect 38669 5185 38703 5219
rect 39589 5185 39623 5219
rect 40417 5185 40451 5219
rect 40877 5185 40911 5219
rect 47869 5185 47903 5219
rect 37381 5117 37415 5151
rect 38393 5117 38427 5151
rect 42533 5117 42567 5151
rect 43545 5117 43579 5151
rect 48053 5049 48087 5083
rect 18429 4981 18463 5015
rect 21925 4981 21959 5015
rect 22569 4981 22603 5015
rect 40233 4981 40267 5015
rect 40877 4981 40911 5015
rect 39221 4777 39255 4811
rect 42533 4777 42567 4811
rect 22201 4709 22235 4743
rect 22845 4641 22879 4675
rect 38485 4641 38519 4675
rect 40233 4641 40267 4675
rect 40417 4641 40451 4675
rect 47593 4641 47627 4675
rect 9505 4573 9539 4607
rect 18061 4573 18095 4607
rect 19257 4573 19291 4607
rect 20085 4573 20119 4607
rect 20177 4573 20211 4607
rect 20821 4573 20855 4607
rect 21465 4573 21499 4607
rect 22109 4573 22143 4607
rect 22753 4573 22787 4607
rect 23581 4573 23615 4607
rect 25789 4573 25823 4607
rect 39129 4573 39163 4607
rect 42717 4573 42751 4607
rect 46673 4573 46707 4607
rect 47317 4573 47351 4607
rect 21557 4505 21591 4539
rect 37473 4505 37507 4539
rect 37565 4505 37599 4539
rect 42073 4505 42107 4539
rect 18153 4437 18187 4471
rect 19349 4437 19383 4471
rect 20913 4437 20947 4471
rect 23397 4437 23431 4471
rect 46765 4437 46799 4471
rect 21005 4233 21039 4267
rect 21925 4233 21959 4267
rect 37289 4233 37323 4267
rect 40877 4233 40911 4267
rect 25237 4165 25271 4199
rect 40049 4165 40083 4199
rect 40509 4165 40543 4199
rect 42901 4165 42935 4199
rect 43821 4165 43855 4199
rect 47777 4165 47811 4199
rect 2145 4097 2179 4131
rect 2881 4097 2915 4131
rect 8861 4097 8895 4131
rect 10057 4097 10091 4131
rect 13737 4097 13771 4131
rect 17325 4097 17359 4131
rect 17969 4097 18003 4131
rect 18981 4097 19015 4131
rect 19625 4097 19659 4131
rect 20269 4097 20303 4131
rect 20913 4097 20947 4131
rect 21833 4097 21867 4131
rect 22477 4097 22511 4131
rect 23121 4097 23155 4131
rect 23213 4097 23247 4131
rect 23765 4097 23799 4131
rect 37473 4097 37507 4131
rect 39589 4097 39623 4131
rect 40693 4097 40727 4131
rect 46765 4097 46799 4131
rect 17417 4029 17451 4063
rect 23857 4029 23891 4063
rect 25145 4029 25179 4063
rect 26065 4029 26099 4063
rect 39405 4029 39439 4063
rect 42809 4029 42843 4063
rect 48053 4029 48087 4063
rect 19717 3961 19751 3995
rect 46949 3961 46983 3995
rect 1685 3893 1719 3927
rect 2237 3893 2271 3927
rect 2973 3893 3007 3927
rect 6561 3893 6595 3927
rect 7205 3893 7239 3927
rect 8953 3893 8987 3927
rect 10149 3893 10183 3927
rect 11713 3893 11747 3927
rect 13829 3893 13863 3927
rect 18061 3893 18095 3927
rect 19073 3893 19107 3927
rect 20361 3893 20395 3927
rect 22569 3893 22603 3927
rect 46305 3893 46339 3927
rect 17141 3689 17175 3723
rect 20913 3689 20947 3723
rect 21557 3689 21591 3723
rect 23765 3689 23799 3723
rect 24501 3689 24535 3723
rect 40141 3689 40175 3723
rect 1409 3553 1443 3587
rect 1593 3553 1627 3587
rect 2329 3553 2363 3587
rect 5917 3553 5951 3587
rect 6469 3553 6503 3587
rect 9229 3553 9263 3587
rect 9689 3553 9723 3587
rect 26893 3553 26927 3587
rect 46305 3553 46339 3587
rect 46489 3553 46523 3587
rect 3985 3485 4019 3519
rect 5273 3485 5307 3519
rect 8401 3485 8435 3519
rect 11989 3485 12023 3519
rect 14289 3485 14323 3519
rect 17049 3485 17083 3519
rect 17693 3485 17727 3519
rect 18337 3485 18371 3519
rect 19533 3485 19567 3519
rect 20361 3485 20395 3519
rect 20821 3485 20855 3519
rect 21465 3485 21499 3519
rect 22569 3485 22603 3519
rect 23029 3485 23063 3519
rect 23673 3485 23707 3519
rect 24409 3485 24443 3519
rect 25513 3485 25547 3519
rect 33057 3485 33091 3519
rect 33885 3485 33919 3519
rect 40049 3485 40083 3519
rect 40785 3485 40819 3519
rect 43085 3485 43119 3519
rect 43913 3485 43947 3519
rect 45201 3485 45235 3519
rect 45661 3485 45695 3519
rect 5365 3417 5399 3451
rect 6101 3417 6135 3451
rect 9413 3417 9447 3451
rect 18429 3417 18463 3451
rect 23121 3417 23155 3451
rect 25697 3417 25731 3451
rect 40969 3417 41003 3451
rect 42625 3417 42659 3451
rect 48145 3417 48179 3451
rect 12081 3349 12115 3383
rect 17785 3349 17819 3383
rect 19625 3349 19659 3383
rect 33149 3349 33183 3383
rect 43177 3349 43211 3383
rect 45753 3349 45787 3383
rect 37749 3145 37783 3179
rect 39681 3145 39715 3179
rect 40969 3145 41003 3179
rect 47869 3145 47903 3179
rect 2237 3077 2271 3111
rect 8125 3077 8159 3111
rect 11713 3077 11747 3111
rect 14013 3077 14047 3111
rect 17785 3077 17819 3111
rect 18889 3077 18923 3111
rect 19625 3077 19659 3111
rect 22477 3077 22511 3111
rect 25145 3077 25179 3111
rect 25237 3077 25271 3111
rect 26157 3077 26191 3111
rect 33149 3077 33183 3111
rect 43085 3077 43119 3111
rect 45385 3077 45419 3111
rect 2053 3009 2087 3043
rect 6653 3009 6687 3043
rect 7941 3009 7975 3043
rect 11529 3009 11563 3043
rect 13829 3009 13863 3043
rect 16865 3009 16899 3043
rect 17693 3009 17727 3043
rect 18797 3009 18831 3043
rect 22293 3009 22327 3043
rect 27169 3009 27203 3043
rect 32965 3009 32999 3043
rect 37289 3009 37323 3043
rect 39221 3009 39255 3043
rect 39865 3009 39899 3043
rect 41613 3009 41647 3043
rect 45201 3009 45235 3043
rect 47777 3009 47811 3043
rect 2973 2941 3007 2975
rect 8401 2941 8435 2975
rect 11989 2941 12023 2975
rect 14289 2941 14323 2975
rect 16773 2941 16807 2975
rect 17233 2941 17267 2975
rect 19441 2941 19475 2975
rect 20453 2941 20487 2975
rect 22753 2941 22787 2975
rect 33517 2941 33551 2975
rect 40325 2941 40359 2975
rect 40509 2941 40543 2975
rect 42901 2941 42935 2975
rect 44005 2941 44039 2975
rect 47041 2941 47075 2975
rect 39037 2873 39071 2907
rect 41429 2873 41463 2907
rect 6745 2805 6779 2839
rect 26985 2805 27019 2839
rect 37381 2805 37415 2839
rect 9137 2601 9171 2635
rect 17509 2601 17543 2635
rect 18153 2601 18187 2635
rect 24685 2601 24719 2635
rect 25513 2601 25547 2635
rect 26341 2601 26375 2635
rect 28641 2601 28675 2635
rect 29745 2601 29779 2635
rect 36369 2601 36403 2635
rect 40417 2601 40451 2635
rect 40601 2601 40635 2635
rect 42533 2601 42567 2635
rect 42901 2601 42935 2635
rect 16865 2533 16899 2567
rect 20545 2533 20579 2567
rect 25697 2533 25731 2567
rect 27629 2533 27663 2567
rect 41337 2533 41371 2567
rect 5273 2465 5307 2499
rect 6561 2465 6595 2499
rect 6745 2465 6779 2499
rect 7113 2465 7147 2499
rect 38393 2465 38427 2499
rect 39313 2465 39347 2499
rect 46489 2465 46523 2499
rect 47869 2465 47903 2499
rect 4997 2397 5031 2431
rect 8953 2397 8987 2431
rect 16681 2397 16715 2431
rect 17417 2397 17451 2431
rect 18061 2397 18095 2431
rect 21281 2397 21315 2431
rect 22109 2397 22143 2431
rect 22937 2397 22971 2431
rect 23305 2397 23339 2431
rect 25237 2397 25271 2431
rect 26157 2397 26191 2431
rect 29929 2397 29963 2431
rect 35725 2397 35759 2431
rect 40049 2397 40083 2431
rect 40417 2397 40451 2431
rect 41153 2397 41187 2431
rect 42441 2397 42475 2431
rect 43637 2397 43671 2431
rect 43913 2397 43947 2431
rect 46213 2397 46247 2431
rect 47685 2397 47719 2431
rect 1869 2329 1903 2363
rect 2789 2329 2823 2363
rect 3157 2329 3191 2363
rect 15669 2329 15703 2363
rect 20361 2329 20395 2363
rect 21097 2329 21131 2363
rect 24593 2329 24627 2363
rect 27445 2329 27479 2363
rect 28549 2329 28583 2363
rect 36277 2329 36311 2363
rect 38209 2329 38243 2363
rect 39129 2329 39163 2363
rect 45385 2329 45419 2363
rect 2145 2261 2179 2295
rect 15761 2261 15795 2295
rect 35541 2261 35575 2295
rect 45477 2261 45511 2295
<< metal1 >>
rect 13354 47540 13360 47592
rect 13412 47580 13418 47592
rect 20530 47580 20536 47592
rect 13412 47552 20536 47580
rect 13412 47540 13418 47552
rect 20530 47540 20536 47552
rect 20588 47540 20594 47592
rect 6638 47472 6644 47524
rect 6696 47512 6702 47524
rect 37366 47512 37372 47524
rect 6696 47484 37372 47512
rect 6696 47472 6702 47484
rect 37366 47472 37372 47484
rect 37424 47472 37430 47524
rect 2038 47404 2044 47456
rect 2096 47444 2102 47456
rect 38194 47444 38200 47456
rect 2096 47416 38200 47444
rect 2096 47404 2102 47416
rect 38194 47404 38200 47416
rect 38252 47404 38258 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 13354 47240 13360 47252
rect 13315 47212 13360 47240
rect 13354 47200 13360 47212
rect 13412 47200 13418 47252
rect 38194 47200 38200 47252
rect 38252 47240 38258 47252
rect 40494 47240 40500 47252
rect 38252 47212 40500 47240
rect 38252 47200 38258 47212
rect 40494 47200 40500 47212
rect 40552 47200 40558 47252
rect 9585 47175 9643 47181
rect 9585 47141 9597 47175
rect 9631 47172 9643 47175
rect 28994 47172 29000 47184
rect 9631 47144 29000 47172
rect 9631 47141 9643 47144
rect 9585 47135 9643 47141
rect 28994 47132 29000 47144
rect 29052 47132 29058 47184
rect 29822 47132 29828 47184
rect 29880 47172 29886 47184
rect 29917 47175 29975 47181
rect 29917 47172 29929 47175
rect 29880 47144 29929 47172
rect 29880 47132 29886 47144
rect 29917 47141 29929 47144
rect 29963 47141 29975 47175
rect 29917 47135 29975 47141
rect 33686 47132 33692 47184
rect 33744 47172 33750 47184
rect 48133 47175 48191 47181
rect 48133 47172 48145 47175
rect 33744 47144 48145 47172
rect 33744 47132 33750 47144
rect 48133 47141 48145 47144
rect 48179 47141 48191 47175
rect 48133 47135 48191 47141
rect 2038 47104 2044 47116
rect 1999 47076 2044 47104
rect 2038 47064 2044 47076
rect 2096 47064 2102 47116
rect 6638 47104 6644 47116
rect 6599 47076 6644 47104
rect 6638 47064 6644 47076
rect 6696 47064 6702 47116
rect 18690 47104 18696 47116
rect 6886 47076 18276 47104
rect 1765 47039 1823 47045
rect 1765 47005 1777 47039
rect 1811 47036 1823 47039
rect 1946 47036 1952 47048
rect 1811 47008 1952 47036
rect 1811 47005 1823 47008
rect 1765 46999 1823 47005
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4706 47036 4712 47048
rect 4667 47008 4712 47036
rect 3789 46999 3847 47005
rect 4706 46996 4712 47008
rect 4764 46996 4770 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6365 47039 6423 47045
rect 6365 47036 6377 47039
rect 5868 47008 6377 47036
rect 5868 46996 5874 47008
rect 6365 47005 6377 47008
rect 6411 47005 6423 47039
rect 6365 46999 6423 47005
rect 2777 46971 2835 46977
rect 2777 46937 2789 46971
rect 2823 46937 2835 46971
rect 2777 46931 2835 46937
rect 2590 46860 2596 46912
rect 2648 46900 2654 46912
rect 2792 46900 2820 46931
rect 3050 46928 3056 46980
rect 3108 46968 3114 46980
rect 3145 46971 3203 46977
rect 3145 46968 3157 46971
rect 3108 46940 3157 46968
rect 3108 46928 3114 46940
rect 3145 46937 3157 46940
rect 3191 46937 3203 46971
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 3145 46931 3203 46937
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 4985 46971 5043 46977
rect 4985 46937 4997 46971
rect 5031 46968 5043 46971
rect 6886 46968 6914 47076
rect 7282 47036 7288 47048
rect 7243 47008 7288 47036
rect 7282 46996 7288 47008
rect 7340 46996 7346 47048
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 9088 47008 9413 47036
rect 9088 46996 9094 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 11606 47036 11612 47048
rect 11567 47008 11612 47036
rect 9401 46999 9459 47005
rect 11606 46996 11612 47008
rect 11664 46996 11670 47048
rect 12250 46996 12256 47048
rect 12308 47036 12314 47048
rect 12345 47039 12403 47045
rect 12345 47036 12357 47039
rect 12308 47008 12357 47036
rect 12308 46996 12314 47008
rect 12345 47005 12357 47008
rect 12391 47005 12403 47039
rect 12345 46999 12403 47005
rect 12894 46996 12900 47048
rect 12952 47036 12958 47048
rect 13081 47039 13139 47045
rect 13081 47036 13093 47039
rect 12952 47008 13093 47036
rect 12952 46996 12958 47008
rect 13081 47005 13093 47008
rect 13127 47005 13139 47039
rect 13081 46999 13139 47005
rect 16482 46996 16488 47048
rect 16540 47036 16546 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16540 47008 16681 47036
rect 16540 46996 16546 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16942 47036 16948 47048
rect 16903 47008 16948 47036
rect 16669 46999 16727 47005
rect 16942 46996 16948 47008
rect 17000 46996 17006 47048
rect 5031 46940 6914 46968
rect 5031 46937 5043 46940
rect 4985 46931 5043 46937
rect 11698 46928 11704 46980
rect 11756 46968 11762 46980
rect 11793 46971 11851 46977
rect 11793 46968 11805 46971
rect 11756 46940 11805 46968
rect 11756 46928 11762 46940
rect 11793 46937 11805 46940
rect 11839 46937 11851 46971
rect 11793 46931 11851 46937
rect 12434 46928 12440 46980
rect 12492 46968 12498 46980
rect 12529 46971 12587 46977
rect 12529 46968 12541 46971
rect 12492 46940 12541 46968
rect 12492 46928 12498 46940
rect 12529 46937 12541 46940
rect 12575 46937 12587 46971
rect 12529 46931 12587 46937
rect 14553 46971 14611 46977
rect 14553 46937 14565 46971
rect 14599 46937 14611 46971
rect 14734 46968 14740 46980
rect 14695 46940 14740 46968
rect 14553 46931 14611 46937
rect 7466 46900 7472 46912
rect 2648 46872 2820 46900
rect 7427 46872 7472 46900
rect 2648 46860 2654 46872
rect 7466 46860 7472 46872
rect 7524 46860 7530 46912
rect 13538 46860 13544 46912
rect 13596 46900 13602 46912
rect 14568 46900 14596 46931
rect 14734 46928 14740 46940
rect 14792 46928 14798 46980
rect 18248 46968 18276 47076
rect 18340 47076 18696 47104
rect 18340 47045 18368 47076
rect 18690 47064 18696 47076
rect 18748 47064 18754 47116
rect 19978 47064 19984 47116
rect 20036 47104 20042 47116
rect 20073 47107 20131 47113
rect 20073 47104 20085 47107
rect 20036 47076 20085 47104
rect 20036 47064 20042 47076
rect 20073 47073 20085 47076
rect 20119 47073 20131 47107
rect 28902 47104 28908 47116
rect 20073 47067 20131 47073
rect 26206 47076 28908 47104
rect 18325 47039 18383 47045
rect 18325 47005 18337 47039
rect 18371 47005 18383 47039
rect 20346 47036 20352 47048
rect 18325 46999 18383 47005
rect 18432 47008 18828 47036
rect 20307 47008 20352 47036
rect 18432 46968 18460 47008
rect 18690 46968 18696 46980
rect 18248 46940 18460 46968
rect 18651 46940 18696 46968
rect 18690 46928 18696 46940
rect 18748 46928 18754 46980
rect 18800 46968 18828 47008
rect 20346 46996 20352 47008
rect 20404 46996 20410 47048
rect 24854 47036 24860 47048
rect 24815 47008 24860 47036
rect 24854 46996 24860 47008
rect 24912 46996 24918 47048
rect 25498 47036 25504 47048
rect 25459 47008 25504 47036
rect 25498 46996 25504 47008
rect 25556 46996 25562 47048
rect 26206 46968 26234 47076
rect 28902 47064 28908 47076
rect 28960 47064 28966 47116
rect 44450 47104 44456 47116
rect 43180 47076 44456 47104
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28537 47039 28595 47045
rect 28537 47036 28549 47039
rect 28408 47008 28549 47036
rect 28408 46996 28414 47008
rect 28537 47005 28549 47008
rect 28583 47005 28595 47039
rect 28537 46999 28595 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 30926 46996 30932 47048
rect 30984 47036 30990 47048
rect 31113 47039 31171 47045
rect 31113 47036 31125 47039
rect 30984 47008 31125 47036
rect 30984 46996 30990 47008
rect 31113 47005 31125 47008
rect 31159 47005 31171 47039
rect 31113 46999 31171 47005
rect 38194 46996 38200 47048
rect 38252 47036 38258 47048
rect 38381 47039 38439 47045
rect 38381 47036 38393 47039
rect 38252 47008 38393 47036
rect 38252 46996 38258 47008
rect 38381 47005 38393 47008
rect 38427 47005 38439 47039
rect 42702 47036 42708 47048
rect 42663 47008 42708 47036
rect 38381 46999 38439 47005
rect 42702 46996 42708 47008
rect 42760 46996 42766 47048
rect 43180 47045 43208 47076
rect 44450 47064 44456 47076
rect 44508 47064 44514 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 43165 47039 43223 47045
rect 43165 47005 43177 47039
rect 43211 47005 43223 47039
rect 43165 46999 43223 47005
rect 43806 46996 43812 47048
rect 43864 47036 43870 47048
rect 43993 47039 44051 47045
rect 43993 47036 44005 47039
rect 43864 47008 44005 47036
rect 43864 46996 43870 47008
rect 43993 47005 44005 47008
rect 44039 47005 44051 47039
rect 45186 47036 45192 47048
rect 45147 47008 45192 47036
rect 43993 46999 44051 47005
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47949 47039 48007 47045
rect 47949 47036 47961 47039
rect 47728 47008 47961 47036
rect 47728 46996 47734 47008
rect 47949 47005 47961 47008
rect 47995 47005 48007 47039
rect 47949 46999 48007 47005
rect 28718 46968 28724 46980
rect 18800 46940 26234 46968
rect 28679 46940 28724 46968
rect 28718 46928 28724 46940
rect 28776 46928 28782 46980
rect 31297 46971 31355 46977
rect 31297 46937 31309 46971
rect 31343 46968 31355 46971
rect 31386 46968 31392 46980
rect 31343 46940 31392 46968
rect 31343 46937 31355 46940
rect 31297 46931 31355 46937
rect 31386 46928 31392 46940
rect 31444 46928 31450 46980
rect 40313 46971 40371 46977
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 40313 46931 40371 46937
rect 13596 46872 14596 46900
rect 13596 46860 13602 46872
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 40402 46928 40408 46980
rect 40460 46968 40466 46980
rect 40497 46971 40555 46977
rect 40497 46968 40509 46971
rect 40460 46940 40509 46968
rect 40460 46928 40466 46940
rect 40497 46937 40509 46940
rect 40543 46937 40555 46971
rect 40497 46931 40555 46937
rect 44177 46971 44235 46977
rect 44177 46937 44189 46971
rect 44223 46968 44235 46971
rect 44358 46968 44364 46980
rect 44223 46940 44364 46968
rect 44223 46937 44235 46940
rect 44177 46931 44235 46937
rect 44358 46928 44364 46940
rect 44416 46928 44422 46980
rect 45373 46971 45431 46977
rect 45373 46937 45385 46971
rect 45419 46968 45431 46971
rect 45462 46968 45468 46980
rect 45419 46940 45468 46968
rect 45419 46937 45431 46940
rect 45373 46931 45431 46937
rect 45462 46928 45468 46940
rect 45520 46928 45526 46980
rect 39356 46872 40356 46900
rect 39356 46860 39362 46872
rect 41874 46860 41880 46912
rect 41932 46900 41938 46912
rect 42886 46900 42892 46912
rect 41932 46872 42892 46900
rect 41932 46860 41938 46872
rect 42886 46860 42892 46872
rect 42944 46860 42950 46912
rect 43346 46900 43352 46912
rect 43307 46872 43352 46900
rect 43346 46860 43352 46872
rect 43404 46860 43410 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 1854 46628 1860 46640
rect 1815 46600 1860 46628
rect 1854 46588 1860 46600
rect 1912 46588 1918 46640
rect 24854 46628 24860 46640
rect 24596 46600 24860 46628
rect 24596 46569 24624 46600
rect 24854 46588 24860 46600
rect 24912 46588 24918 46640
rect 43162 46588 43168 46640
rect 43220 46628 43226 46640
rect 44545 46631 44603 46637
rect 44545 46628 44557 46631
rect 43220 46600 44557 46628
rect 43220 46588 43226 46600
rect 44545 46597 44557 46600
rect 44591 46597 44603 46631
rect 47026 46628 47032 46640
rect 46987 46600 47032 46628
rect 44545 46591 44603 46597
rect 47026 46588 47032 46600
rect 47084 46588 47090 46640
rect 24581 46563 24639 46569
rect 24581 46529 24593 46563
rect 24627 46529 24639 46563
rect 38194 46560 38200 46572
rect 38155 46532 38200 46560
rect 24581 46523 24639 46529
rect 38194 46520 38200 46532
rect 38252 46520 38258 46572
rect 42702 46560 42708 46572
rect 42663 46532 42708 46560
rect 42702 46520 42708 46532
rect 42760 46520 42766 46572
rect 47946 46560 47952 46572
rect 47907 46532 47952 46560
rect 47946 46520 47952 46532
rect 48004 46520 48010 46572
rect 3421 46495 3479 46501
rect 3421 46461 3433 46495
rect 3467 46461 3479 46495
rect 3421 46455 3479 46461
rect 3605 46495 3663 46501
rect 3605 46461 3617 46495
rect 3651 46492 3663 46495
rect 3878 46492 3884 46504
rect 3651 46464 3884 46492
rect 3651 46461 3663 46464
rect 3605 46455 3663 46461
rect 3436 46424 3464 46455
rect 3878 46452 3884 46464
rect 3936 46452 3942 46504
rect 3970 46452 3976 46504
rect 4028 46492 4034 46504
rect 4157 46495 4215 46501
rect 4157 46492 4169 46495
rect 4028 46464 4169 46492
rect 4028 46452 4034 46464
rect 4157 46461 4169 46464
rect 4203 46461 4215 46495
rect 4157 46455 4215 46461
rect 13081 46495 13139 46501
rect 13081 46461 13093 46495
rect 13127 46492 13139 46495
rect 13541 46495 13599 46501
rect 13541 46492 13553 46495
rect 13127 46464 13553 46492
rect 13127 46461 13139 46464
rect 13081 46455 13139 46461
rect 13541 46461 13553 46464
rect 13587 46461 13599 46495
rect 13541 46455 13599 46461
rect 13725 46495 13783 46501
rect 13725 46461 13737 46495
rect 13771 46492 13783 46495
rect 14182 46492 14188 46504
rect 13771 46464 14188 46492
rect 13771 46461 13783 46464
rect 13725 46455 13783 46461
rect 14182 46452 14188 46464
rect 14240 46452 14246 46504
rect 14274 46452 14280 46504
rect 14332 46492 14338 46504
rect 19426 46492 19432 46504
rect 14332 46464 14377 46492
rect 19387 46464 19432 46492
rect 14332 46452 14338 46464
rect 19426 46452 19432 46464
rect 19484 46452 19490 46504
rect 19613 46495 19671 46501
rect 19613 46461 19625 46495
rect 19659 46492 19671 46495
rect 20254 46492 20260 46504
rect 19659 46464 20260 46492
rect 19659 46461 19671 46464
rect 19613 46455 19671 46461
rect 20254 46452 20260 46464
rect 20312 46452 20318 46504
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 24762 46492 24768 46504
rect 24723 46464 24768 46492
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 25130 46492 25136 46504
rect 25091 46464 25136 46492
rect 25130 46452 25136 46464
rect 25188 46452 25194 46504
rect 32398 46492 32404 46504
rect 32359 46464 32404 46492
rect 32398 46452 32404 46464
rect 32456 46452 32462 46504
rect 32585 46495 32643 46501
rect 32585 46461 32597 46495
rect 32631 46492 32643 46495
rect 33318 46492 33324 46504
rect 32631 46464 33324 46492
rect 32631 46461 32643 46464
rect 32585 46455 32643 46461
rect 33318 46452 33324 46464
rect 33376 46452 33382 46504
rect 33413 46495 33471 46501
rect 33413 46461 33425 46495
rect 33459 46461 33471 46495
rect 38378 46492 38384 46504
rect 38339 46464 38384 46492
rect 33413 46455 33471 46461
rect 4614 46424 4620 46436
rect 3436 46396 4620 46424
rect 4614 46384 4620 46396
rect 4672 46384 4678 46436
rect 32214 46384 32220 46436
rect 32272 46424 32278 46436
rect 33428 46424 33456 46455
rect 38378 46452 38384 46464
rect 38436 46452 38442 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46492 42947 46495
rect 43806 46492 43812 46504
rect 42935 46464 43812 46492
rect 42935 46461 42947 46464
rect 42889 46455 42947 46461
rect 43806 46452 43812 46464
rect 43864 46452 43870 46504
rect 45189 46495 45247 46501
rect 45189 46461 45201 46495
rect 45235 46461 45247 46495
rect 45370 46492 45376 46504
rect 45331 46464 45376 46492
rect 45189 46455 45247 46461
rect 32272 46396 33456 46424
rect 45204 46424 45232 46455
rect 45370 46452 45376 46464
rect 45428 46452 45434 46504
rect 45554 46424 45560 46436
rect 45204 46396 45560 46424
rect 32272 46384 32278 46396
rect 45554 46384 45560 46396
rect 45612 46384 45618 46436
rect 2133 46359 2191 46365
rect 2133 46325 2145 46359
rect 2179 46356 2191 46359
rect 2314 46356 2320 46368
rect 2179 46328 2320 46356
rect 2179 46325 2191 46328
rect 2133 46319 2191 46325
rect 2314 46316 2320 46328
rect 2372 46316 2378 46368
rect 2866 46356 2872 46368
rect 2827 46328 2872 46356
rect 2866 46316 2872 46328
rect 2924 46316 2930 46368
rect 10502 46316 10508 46368
rect 10560 46356 10566 46368
rect 10781 46359 10839 46365
rect 10781 46356 10793 46359
rect 10560 46328 10793 46356
rect 10560 46316 10566 46328
rect 10781 46325 10793 46328
rect 10827 46325 10839 46359
rect 10781 46319 10839 46325
rect 20806 46316 20812 46368
rect 20864 46356 20870 46368
rect 22005 46359 22063 46365
rect 22005 46356 22017 46359
rect 20864 46328 22017 46356
rect 20864 46316 20870 46328
rect 22005 46325 22017 46328
rect 22051 46325 22063 46359
rect 22005 46319 22063 46325
rect 41414 46316 41420 46368
rect 41472 46356 41478 46368
rect 41601 46359 41659 46365
rect 41601 46356 41613 46359
rect 41472 46328 41613 46356
rect 41472 46316 41478 46328
rect 41601 46325 41613 46328
rect 41647 46325 41659 46359
rect 41601 46319 41659 46325
rect 47854 46316 47860 46368
rect 47912 46356 47918 46368
rect 48041 46359 48099 46365
rect 48041 46356 48053 46359
rect 47912 46328 48053 46356
rect 47912 46316 47918 46328
rect 48041 46325 48053 46328
rect 48087 46325 48099 46359
rect 48041 46319 48099 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 3878 46152 3884 46164
rect 3839 46124 3884 46152
rect 3878 46112 3884 46124
rect 3936 46112 3942 46164
rect 4614 46152 4620 46164
rect 4575 46124 4620 46152
rect 4614 46112 4620 46124
rect 4672 46112 4678 46164
rect 14182 46152 14188 46164
rect 14143 46124 14188 46152
rect 14182 46112 14188 46124
rect 14240 46112 14246 46164
rect 19426 46112 19432 46164
rect 19484 46152 19490 46164
rect 20349 46155 20407 46161
rect 20349 46152 20361 46155
rect 19484 46124 20361 46152
rect 19484 46112 19490 46124
rect 20349 46121 20361 46124
rect 20395 46121 20407 46155
rect 20349 46115 20407 46121
rect 24673 46155 24731 46161
rect 24673 46121 24685 46155
rect 24719 46152 24731 46155
rect 24762 46152 24768 46164
rect 24719 46124 24768 46152
rect 24719 46121 24731 46124
rect 24673 46115 24731 46121
rect 24762 46112 24768 46124
rect 24820 46112 24826 46164
rect 32398 46112 32404 46164
rect 32456 46152 32462 46164
rect 32677 46155 32735 46161
rect 32677 46152 32689 46155
rect 32456 46124 32689 46152
rect 32456 46112 32462 46124
rect 32677 46121 32689 46124
rect 32723 46121 32735 46155
rect 38378 46152 38384 46164
rect 38339 46124 38384 46152
rect 32677 46115 32735 46121
rect 38378 46112 38384 46124
rect 38436 46112 38442 46164
rect 43806 46152 43812 46164
rect 43767 46124 43812 46152
rect 43806 46112 43812 46124
rect 43864 46112 43870 46164
rect 16546 46056 43760 46084
rect 10502 46016 10508 46028
rect 10463 45988 10508 46016
rect 10502 45976 10508 45988
rect 10560 45976 10566 46028
rect 10962 45976 10968 46028
rect 11020 46016 11026 46028
rect 11057 46019 11115 46025
rect 11057 46016 11069 46019
rect 11020 45988 11069 46016
rect 11020 45976 11026 45988
rect 11057 45985 11069 45988
rect 11103 45985 11115 46019
rect 11057 45979 11115 45985
rect 2869 45951 2927 45957
rect 2869 45917 2881 45951
rect 2915 45917 2927 45951
rect 2869 45911 2927 45917
rect 2884 45880 2912 45911
rect 3142 45908 3148 45960
rect 3200 45948 3206 45960
rect 3789 45951 3847 45957
rect 3789 45948 3801 45951
rect 3200 45920 3801 45948
rect 3200 45908 3206 45920
rect 3789 45917 3801 45920
rect 3835 45917 3847 45951
rect 3789 45911 3847 45917
rect 14093 45951 14151 45957
rect 14093 45917 14105 45951
rect 14139 45948 14151 45951
rect 16546 45948 16574 46056
rect 20806 46016 20812 46028
rect 20767 45988 20812 46016
rect 20806 45976 20812 45988
rect 20864 45976 20870 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 25225 46019 25283 46025
rect 25225 45985 25237 46019
rect 25271 46016 25283 46019
rect 25498 46016 25504 46028
rect 25271 45988 25504 46016
rect 25271 45985 25283 45988
rect 25225 45979 25283 45985
rect 25498 45976 25504 45988
rect 25556 45976 25562 46028
rect 26605 46019 26663 46025
rect 26605 45985 26617 46019
rect 26651 45985 26663 46019
rect 41414 46016 41420 46028
rect 41375 45988 41420 46016
rect 26605 45979 26663 45985
rect 14139 45920 16574 45948
rect 24581 45951 24639 45957
rect 14139 45917 14151 45920
rect 14093 45911 14151 45917
rect 24581 45917 24593 45951
rect 24627 45948 24639 45951
rect 24854 45948 24860 45960
rect 24627 45920 24860 45948
rect 24627 45917 24639 45920
rect 24581 45911 24639 45917
rect 24854 45908 24860 45920
rect 24912 45908 24918 45960
rect 10686 45880 10692 45892
rect 2884 45852 6914 45880
rect 10647 45852 10692 45880
rect 2958 45812 2964 45824
rect 2919 45784 2964 45812
rect 2958 45772 2964 45784
rect 3016 45772 3022 45824
rect 6886 45812 6914 45852
rect 10686 45840 10692 45852
rect 10744 45840 10750 45892
rect 20990 45880 20996 45892
rect 20951 45852 20996 45880
rect 20990 45840 20996 45852
rect 21048 45840 21054 45892
rect 25406 45880 25412 45892
rect 25367 45852 25412 45880
rect 25406 45840 25412 45852
rect 25464 45840 25470 45892
rect 10594 45812 10600 45824
rect 6886 45784 10600 45812
rect 10594 45772 10600 45784
rect 10652 45772 10658 45824
rect 25774 45772 25780 45824
rect 25832 45812 25838 45824
rect 26620 45812 26648 45979
rect 41414 45976 41420 45988
rect 41472 45976 41478 46028
rect 42518 46016 42524 46028
rect 42479 45988 42524 46016
rect 42518 45976 42524 45988
rect 42576 45976 42582 46028
rect 43732 46016 43760 46056
rect 45830 46016 45836 46028
rect 43732 45988 45836 46016
rect 38289 45951 38347 45957
rect 38289 45917 38301 45951
rect 38335 45948 38347 45951
rect 40310 45948 40316 45960
rect 38335 45920 40316 45948
rect 38335 45917 38347 45920
rect 38289 45911 38347 45917
rect 40310 45908 40316 45920
rect 40368 45908 40374 45960
rect 43732 45957 43760 45988
rect 45830 45976 45836 45988
rect 45888 45976 45894 46028
rect 46293 46019 46351 46025
rect 46293 45985 46305 46019
rect 46339 46016 46351 46019
rect 46750 46016 46756 46028
rect 46339 45988 46756 46016
rect 46339 45985 46351 45988
rect 46293 45979 46351 45985
rect 46750 45976 46756 45988
rect 46808 45976 46814 46028
rect 48130 46016 48136 46028
rect 48091 45988 48136 46016
rect 48130 45976 48136 45988
rect 48188 45976 48194 46028
rect 43717 45951 43775 45957
rect 43717 45917 43729 45951
rect 43763 45917 43775 45951
rect 43717 45911 43775 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45948 45707 45951
rect 45738 45948 45744 45960
rect 45695 45920 45744 45948
rect 45695 45917 45707 45920
rect 45649 45911 45707 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 41598 45880 41604 45892
rect 41559 45852 41604 45880
rect 41598 45840 41604 45852
rect 41656 45840 41662 45892
rect 46477 45883 46535 45889
rect 46477 45849 46489 45883
rect 46523 45880 46535 45883
rect 46934 45880 46940 45892
rect 46523 45852 46940 45880
rect 46523 45849 46535 45852
rect 46477 45843 46535 45849
rect 46934 45840 46940 45852
rect 46992 45840 46998 45892
rect 25832 45784 26648 45812
rect 25832 45772 25838 45784
rect 27338 45772 27344 45824
rect 27396 45812 27402 45824
rect 45741 45815 45799 45821
rect 45741 45812 45753 45815
rect 27396 45784 45753 45812
rect 27396 45772 27402 45784
rect 45741 45781 45753 45784
rect 45787 45781 45799 45815
rect 45741 45775 45799 45781
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 10686 45608 10692 45620
rect 10647 45580 10692 45608
rect 10686 45568 10692 45580
rect 10744 45568 10750 45620
rect 15930 45568 15936 45620
rect 15988 45608 15994 45620
rect 17402 45608 17408 45620
rect 15988 45580 17408 45608
rect 15988 45568 15994 45580
rect 17402 45568 17408 45580
rect 17460 45568 17466 45620
rect 20254 45568 20260 45620
rect 20312 45608 20318 45620
rect 20349 45611 20407 45617
rect 20349 45608 20361 45611
rect 20312 45580 20361 45608
rect 20312 45568 20318 45580
rect 20349 45577 20361 45580
rect 20395 45577 20407 45611
rect 20990 45608 20996 45620
rect 20951 45580 20996 45608
rect 20349 45571 20407 45577
rect 20990 45568 20996 45580
rect 21048 45568 21054 45620
rect 25406 45608 25412 45620
rect 25367 45580 25412 45608
rect 25406 45568 25412 45580
rect 25464 45568 25470 45620
rect 45094 45568 45100 45620
rect 45152 45608 45158 45620
rect 45152 45580 45784 45608
rect 45152 45568 45158 45580
rect 2225 45543 2283 45549
rect 2225 45509 2237 45543
rect 2271 45540 2283 45543
rect 2958 45540 2964 45552
rect 2271 45512 2964 45540
rect 2271 45509 2283 45512
rect 2225 45503 2283 45509
rect 2958 45500 2964 45512
rect 3016 45500 3022 45552
rect 33318 45540 33324 45552
rect 16546 45512 24900 45540
rect 33279 45512 33324 45540
rect 10594 45472 10600 45484
rect 10507 45444 10600 45472
rect 10594 45432 10600 45444
rect 10652 45472 10658 45484
rect 16546 45472 16574 45512
rect 24872 45484 24900 45512
rect 33318 45500 33324 45512
rect 33376 45500 33382 45552
rect 41049 45543 41107 45549
rect 41049 45509 41061 45543
rect 41095 45540 41107 45543
rect 41598 45540 41604 45552
rect 41095 45512 41604 45540
rect 41095 45509 41107 45512
rect 41049 45503 41107 45509
rect 41598 45500 41604 45512
rect 41656 45500 41662 45552
rect 43901 45543 43959 45549
rect 43901 45509 43913 45543
rect 43947 45540 43959 45543
rect 44637 45543 44695 45549
rect 44637 45540 44649 45543
rect 43947 45512 44649 45540
rect 43947 45509 43959 45512
rect 43901 45503 43959 45509
rect 44637 45509 44649 45512
rect 44683 45509 44695 45543
rect 45756 45540 45784 45580
rect 46842 45540 46848 45552
rect 45756 45512 45876 45540
rect 46803 45512 46848 45540
rect 44637 45503 44695 45509
rect 10652 45444 16574 45472
rect 20257 45475 20315 45481
rect 10652 45432 10658 45444
rect 20257 45441 20269 45475
rect 20303 45441 20315 45475
rect 20257 45435 20315 45441
rect 2041 45407 2099 45413
rect 2041 45373 2053 45407
rect 2087 45404 2099 45407
rect 2866 45404 2872 45416
rect 2087 45376 2872 45404
rect 2087 45373 2099 45376
rect 2041 45367 2099 45373
rect 2866 45364 2872 45376
rect 2924 45364 2930 45416
rect 2961 45407 3019 45413
rect 2961 45373 2973 45407
rect 3007 45373 3019 45407
rect 20272 45404 20300 45435
rect 20806 45432 20812 45484
rect 20864 45472 20870 45484
rect 20901 45475 20959 45481
rect 20901 45472 20913 45475
rect 20864 45444 20913 45472
rect 20864 45432 20870 45444
rect 20901 45441 20913 45444
rect 20947 45441 20959 45475
rect 20901 45435 20959 45441
rect 24854 45432 24860 45484
rect 24912 45472 24918 45484
rect 25314 45472 25320 45484
rect 24912 45444 25320 45472
rect 24912 45432 24918 45444
rect 25314 45432 25320 45444
rect 25372 45432 25378 45484
rect 33229 45475 33287 45481
rect 33229 45441 33241 45475
rect 33275 45472 33287 45475
rect 40954 45472 40960 45484
rect 33275 45444 35894 45472
rect 40915 45444 40960 45472
rect 33275 45441 33287 45444
rect 33229 45435 33287 45441
rect 20272 45376 26234 45404
rect 2961 45367 3019 45373
rect 2774 45296 2780 45348
rect 2832 45336 2838 45348
rect 2976 45336 3004 45367
rect 2832 45308 3004 45336
rect 2832 45296 2838 45308
rect 26206 45268 26234 45376
rect 35866 45336 35894 45444
rect 40954 45432 40960 45444
rect 41012 45432 41018 45484
rect 43806 45472 43812 45484
rect 43767 45444 43812 45472
rect 43806 45432 43812 45444
rect 43864 45432 43870 45484
rect 38654 45404 38660 45416
rect 38615 45376 38660 45404
rect 38654 45364 38660 45376
rect 38712 45364 38718 45416
rect 38838 45404 38844 45416
rect 38799 45376 38844 45404
rect 38838 45364 38844 45376
rect 38896 45364 38902 45416
rect 39850 45404 39856 45416
rect 39811 45376 39856 45404
rect 39850 45364 39856 45376
rect 39908 45364 39914 45416
rect 44450 45404 44456 45416
rect 44411 45376 44456 45404
rect 44450 45364 44456 45376
rect 44508 45364 44514 45416
rect 45848 45413 45876 45512
rect 46842 45500 46848 45512
rect 46900 45500 46906 45552
rect 47486 45432 47492 45484
rect 47544 45472 47550 45484
rect 47581 45475 47639 45481
rect 47581 45472 47593 45475
rect 47544 45444 47593 45472
rect 47544 45432 47550 45444
rect 47581 45441 47593 45444
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 45833 45407 45891 45413
rect 45833 45373 45845 45407
rect 45879 45373 45891 45407
rect 45833 45367 45891 45373
rect 38746 45336 38752 45348
rect 35866 45308 38752 45336
rect 38746 45296 38752 45308
rect 38804 45296 38810 45348
rect 45462 45296 45468 45348
rect 45520 45336 45526 45348
rect 47673 45339 47731 45345
rect 47673 45336 47685 45339
rect 45520 45308 47685 45336
rect 45520 45296 45526 45308
rect 47673 45305 47685 45308
rect 47719 45305 47731 45339
rect 47673 45299 47731 45305
rect 36262 45268 36268 45280
rect 26206 45240 36268 45268
rect 36262 45228 36268 45240
rect 36320 45228 36326 45280
rect 41414 45228 41420 45280
rect 41472 45268 41478 45280
rect 41785 45271 41843 45277
rect 41785 45268 41797 45271
rect 41472 45240 41797 45268
rect 41472 45228 41478 45240
rect 41785 45237 41797 45240
rect 41831 45237 41843 45271
rect 41785 45231 41843 45237
rect 43438 45228 43444 45280
rect 43496 45268 43502 45280
rect 46937 45271 46995 45277
rect 46937 45268 46949 45271
rect 43496 45240 46949 45268
rect 43496 45228 43502 45240
rect 46937 45237 46949 45240
rect 46983 45237 46995 45271
rect 46937 45231 46995 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 38838 45064 38844 45076
rect 38799 45036 38844 45064
rect 38838 45024 38844 45036
rect 38896 45024 38902 45076
rect 44450 45064 44456 45076
rect 44411 45036 44456 45064
rect 44450 45024 44456 45036
rect 44508 45024 44514 45076
rect 45097 45067 45155 45073
rect 45097 45033 45109 45067
rect 45143 45064 45155 45067
rect 45370 45064 45376 45076
rect 45143 45036 45376 45064
rect 45143 45033 45155 45036
rect 45097 45027 45155 45033
rect 45370 45024 45376 45036
rect 45428 45024 45434 45076
rect 41414 44928 41420 44940
rect 41375 44900 41420 44928
rect 41414 44888 41420 44900
rect 41472 44888 41478 44940
rect 42886 44928 42892 44940
rect 42847 44900 42892 44928
rect 42886 44888 42892 44900
rect 42944 44888 42950 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 28074 44820 28080 44872
rect 28132 44860 28138 44872
rect 28721 44863 28779 44869
rect 28721 44860 28733 44863
rect 28132 44832 28733 44860
rect 28132 44820 28138 44832
rect 28721 44829 28733 44832
rect 28767 44829 28779 44863
rect 38746 44860 38752 44872
rect 38707 44832 38752 44860
rect 28721 44823 28779 44829
rect 38746 44820 38752 44832
rect 38804 44820 38810 44872
rect 45002 44860 45008 44872
rect 44963 44832 45008 44860
rect 45002 44820 45008 44832
rect 45060 44820 45066 44872
rect 45649 44863 45707 44869
rect 45649 44829 45661 44863
rect 45695 44860 45707 44863
rect 45830 44860 45836 44872
rect 45695 44832 45836 44860
rect 45695 44829 45707 44832
rect 45649 44823 45707 44829
rect 45830 44820 45836 44832
rect 45888 44820 45894 44872
rect 46290 44860 46296 44872
rect 46251 44832 46296 44860
rect 46290 44820 46296 44832
rect 46348 44820 46354 44872
rect 41598 44792 41604 44804
rect 41559 44764 41604 44792
rect 41598 44752 41604 44764
rect 41656 44752 41662 44804
rect 45741 44795 45799 44801
rect 45741 44761 45753 44795
rect 45787 44792 45799 44795
rect 46477 44795 46535 44801
rect 46477 44792 46489 44795
rect 45787 44764 46489 44792
rect 45787 44761 45799 44764
rect 45741 44755 45799 44761
rect 46477 44761 46489 44764
rect 46523 44761 46535 44795
rect 46477 44755 46535 44761
rect 28813 44727 28871 44733
rect 28813 44693 28825 44727
rect 28859 44724 28871 44727
rect 38654 44724 38660 44736
rect 28859 44696 38660 44724
rect 28859 44693 28871 44696
rect 28813 44687 28871 44693
rect 38654 44684 38660 44696
rect 38712 44684 38718 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 41598 44520 41604 44532
rect 41559 44492 41604 44520
rect 41598 44480 41604 44492
rect 41656 44480 41662 44532
rect 46934 44520 46940 44532
rect 46895 44492 46940 44520
rect 46934 44480 46940 44492
rect 46992 44480 46998 44532
rect 41509 44387 41567 44393
rect 41509 44353 41521 44387
rect 41555 44353 41567 44387
rect 41509 44347 41567 44353
rect 41524 44316 41552 44347
rect 45554 44344 45560 44396
rect 45612 44384 45618 44396
rect 45649 44387 45707 44393
rect 45649 44384 45661 44387
rect 45612 44356 45661 44384
rect 45612 44344 45618 44356
rect 45649 44353 45661 44356
rect 45695 44353 45707 44387
rect 45649 44347 45707 44353
rect 46290 44344 46296 44396
rect 46348 44384 46354 44396
rect 46385 44387 46443 44393
rect 46385 44384 46397 44387
rect 46348 44356 46397 44384
rect 46348 44344 46354 44356
rect 46385 44353 46397 44356
rect 46431 44353 46443 44387
rect 46842 44384 46848 44396
rect 46803 44356 46848 44384
rect 46385 44347 46443 44353
rect 46842 44344 46848 44356
rect 46900 44344 46906 44396
rect 47486 44344 47492 44396
rect 47544 44384 47550 44396
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 47544 44356 47593 44384
rect 47544 44344 47550 44356
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 47302 44316 47308 44328
rect 41524 44288 47308 44316
rect 47302 44276 47308 44288
rect 47360 44276 47366 44328
rect 45830 44140 45836 44192
rect 45888 44180 45894 44192
rect 46566 44180 46572 44192
rect 45888 44152 46572 44180
rect 45888 44140 45894 44152
rect 46566 44140 46572 44152
rect 46624 44140 46630 44192
rect 47670 44180 47676 44192
rect 47631 44152 47676 44180
rect 47670 44140 47676 44152
rect 47728 44140 47734 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 45186 43936 45192 43988
rect 45244 43976 45250 43988
rect 45833 43979 45891 43985
rect 45833 43976 45845 43979
rect 45244 43948 45845 43976
rect 45244 43936 45250 43948
rect 45833 43945 45845 43948
rect 45879 43945 45891 43979
rect 45833 43939 45891 43945
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 47670 43840 47676 43852
rect 46523 43812 47676 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 47670 43800 47676 43812
rect 47728 43800 47734 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 46290 43772 46296 43784
rect 46251 43744 46296 43772
rect 46290 43732 46296 43744
rect 46348 43732 46354 43784
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 46290 43256 46296 43308
rect 46348 43296 46354 43308
rect 47029 43299 47087 43305
rect 47029 43296 47041 43299
rect 46348 43268 47041 43296
rect 46348 43256 46354 43268
rect 47029 43265 47041 43268
rect 47075 43265 47087 43299
rect 47029 43259 47087 43265
rect 1486 43188 1492 43240
rect 1544 43228 1550 43240
rect 1581 43231 1639 43237
rect 1581 43228 1593 43231
rect 1544 43200 1593 43228
rect 1544 43188 1550 43200
rect 1581 43197 1593 43200
rect 1627 43197 1639 43231
rect 1581 43191 1639 43197
rect 46750 43188 46756 43240
rect 46808 43228 46814 43240
rect 47765 43231 47823 43237
rect 47765 43228 47777 43231
rect 46808 43200 47777 43228
rect 46808 43188 46814 43200
rect 47765 43197 47777 43200
rect 47811 43197 47823 43231
rect 47765 43191 47823 43197
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46290 42684 46296 42696
rect 46251 42656 46296 42684
rect 46290 42644 46296 42656
rect 46348 42644 46354 42696
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 47670 42616 47676 42628
rect 46523 42588 47676 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 47670 42576 47676 42588
rect 47728 42576 47734 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 47670 42344 47676 42356
rect 47631 42316 47676 42344
rect 47670 42304 47676 42316
rect 47728 42304 47734 42356
rect 46290 42168 46296 42220
rect 46348 42208 46354 42220
rect 47029 42211 47087 42217
rect 47029 42208 47041 42211
rect 46348 42180 47041 42208
rect 46348 42168 46354 42180
rect 47029 42177 47041 42180
rect 47075 42177 47087 42211
rect 47029 42171 47087 42177
rect 47302 42168 47308 42220
rect 47360 42208 47366 42220
rect 47581 42211 47639 42217
rect 47581 42208 47593 42211
rect 47360 42180 47593 42208
rect 47360 42168 47366 42180
rect 47581 42177 47593 42180
rect 47627 42177 47639 42211
rect 47581 42171 47639 42177
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41664 46351 41667
rect 47670 41664 47676 41676
rect 46339 41636 47676 41664
rect 46339 41633 46351 41636
rect 46293 41627 46351 41633
rect 47670 41624 47676 41636
rect 47728 41624 47734 41676
rect 48130 41596 48136 41608
rect 48091 41568 48136 41596
rect 48130 41556 48136 41568
rect 48188 41556 48194 41608
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46477 41531 46535 41537
rect 46477 41497 46489 41531
rect 46523 41528 46535 41531
rect 46934 41528 46940 41540
rect 46523 41500 46940 41528
rect 46523 41497 46535 41500
rect 46477 41491 46535 41497
rect 46934 41488 46940 41500
rect 46992 41488 46998 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2225 41259 2283 41265
rect 2225 41256 2237 41259
rect 1636 41228 2237 41256
rect 1636 41216 1642 41228
rect 2225 41225 2237 41228
rect 2271 41225 2283 41259
rect 46934 41256 46940 41268
rect 46895 41228 46940 41256
rect 2225 41219 2283 41225
rect 46934 41216 46940 41228
rect 46992 41216 46998 41268
rect 2130 41120 2136 41132
rect 2091 41092 2136 41120
rect 2130 41080 2136 41092
rect 2188 41080 2194 41132
rect 46842 41120 46848 41132
rect 46803 41092 46848 41120
rect 46842 41080 46848 41092
rect 46900 41080 46906 41132
rect 47946 41120 47952 41132
rect 47907 41092 47952 41120
rect 47946 41080 47952 41092
rect 48004 41080 48010 41132
rect 48038 40916 48044 40928
rect 47999 40888 48044 40916
rect 48038 40876 48044 40888
rect 48096 40876 48102 40928
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 47670 40712 47676 40724
rect 47631 40684 47676 40712
rect 47670 40672 47676 40684
rect 47728 40672 47734 40724
rect 1394 40508 1400 40520
rect 1355 40480 1400 40508
rect 1394 40468 1400 40480
rect 1452 40468 1458 40520
rect 1581 40375 1639 40381
rect 1581 40341 1593 40375
rect 1627 40372 1639 40375
rect 1670 40372 1676 40384
rect 1627 40344 1676 40372
rect 1627 40341 1639 40344
rect 1581 40335 1639 40341
rect 1670 40332 1676 40344
rect 1728 40332 1734 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 46290 39788 46296 39840
rect 46348 39828 46354 39840
rect 47765 39831 47823 39837
rect 47765 39828 47777 39831
rect 46348 39800 47777 39828
rect 46348 39788 46354 39800
rect 47765 39797 47777 39800
rect 47811 39797 47823 39831
rect 47765 39791 47823 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 40221 39491 40279 39497
rect 40221 39457 40233 39491
rect 40267 39488 40279 39491
rect 40770 39488 40776 39500
rect 40267 39460 40776 39488
rect 40267 39457 40279 39460
rect 40221 39451 40279 39457
rect 40770 39448 40776 39460
rect 40828 39488 40834 39500
rect 40954 39488 40960 39500
rect 40828 39460 40960 39488
rect 40828 39448 40834 39460
rect 40954 39448 40960 39460
rect 41012 39448 41018 39500
rect 46290 39488 46296 39500
rect 46251 39460 46296 39488
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 39945 39423 40003 39429
rect 39945 39389 39957 39423
rect 39991 39420 40003 39423
rect 40126 39420 40132 39432
rect 39991 39392 40132 39420
rect 39991 39389 40003 39392
rect 39945 39383 40003 39389
rect 40126 39380 40132 39392
rect 40184 39380 40190 39432
rect 46477 39355 46535 39361
rect 46477 39321 46489 39355
rect 46523 39352 46535 39355
rect 46934 39352 46940 39364
rect 46523 39324 46940 39352
rect 46523 39321 46535 39324
rect 46477 39315 46535 39321
rect 46934 39312 46940 39324
rect 46992 39312 46998 39364
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 46934 39080 46940 39092
rect 46895 39052 46940 39080
rect 46934 39040 46940 39052
rect 46992 39040 46998 39092
rect 3510 38972 3516 39024
rect 3568 39012 3574 39024
rect 7558 39012 7564 39024
rect 3568 38984 7564 39012
rect 3568 38972 3574 38984
rect 7558 38972 7564 38984
rect 7616 38972 7622 39024
rect 40126 38944 40132 38956
rect 40087 38916 40132 38944
rect 40126 38904 40132 38916
rect 40184 38904 40190 38956
rect 46750 38904 46756 38956
rect 46808 38944 46814 38956
rect 46845 38947 46903 38953
rect 46845 38944 46857 38947
rect 46808 38916 46857 38944
rect 46808 38904 46814 38916
rect 46845 38913 46857 38916
rect 46891 38913 46903 38947
rect 47670 38944 47676 38956
rect 47631 38916 47676 38944
rect 46845 38907 46903 38913
rect 47670 38904 47676 38916
rect 47728 38904 47734 38956
rect 3326 38836 3332 38888
rect 3384 38876 3390 38888
rect 3510 38876 3516 38888
rect 3384 38848 3516 38876
rect 3384 38836 3390 38848
rect 3510 38836 3516 38848
rect 3568 38836 3574 38888
rect 40310 38836 40316 38888
rect 40368 38876 40374 38888
rect 40405 38879 40463 38885
rect 40405 38876 40417 38879
rect 40368 38848 40417 38876
rect 40368 38836 40374 38848
rect 40405 38845 40417 38848
rect 40451 38845 40463 38879
rect 40405 38839 40463 38845
rect 40420 38808 40448 38839
rect 44174 38836 44180 38888
rect 44232 38876 44238 38888
rect 45462 38876 45468 38888
rect 44232 38848 45468 38876
rect 44232 38836 44238 38848
rect 45462 38836 45468 38848
rect 45520 38876 45526 38888
rect 47857 38879 47915 38885
rect 47857 38876 47869 38879
rect 45520 38848 47869 38876
rect 45520 38836 45526 38848
rect 47857 38845 47869 38848
rect 47903 38845 47915 38879
rect 47857 38839 47915 38845
rect 45646 38808 45652 38820
rect 40420 38780 45652 38808
rect 45646 38768 45652 38780
rect 45704 38808 45710 38820
rect 46842 38808 46848 38820
rect 45704 38780 46848 38808
rect 45704 38768 45710 38780
rect 46842 38768 46848 38780
rect 46900 38768 46906 38820
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 41322 38360 41328 38412
rect 41380 38400 41386 38412
rect 41969 38403 42027 38409
rect 41969 38400 41981 38403
rect 41380 38372 41981 38400
rect 41380 38360 41386 38372
rect 41969 38369 41981 38372
rect 42015 38400 42027 38403
rect 45002 38400 45008 38412
rect 42015 38372 45008 38400
rect 42015 38369 42027 38372
rect 41969 38363 42027 38369
rect 45002 38360 45008 38372
rect 45060 38360 45066 38412
rect 39025 38335 39083 38341
rect 39025 38301 39037 38335
rect 39071 38332 39083 38335
rect 44174 38332 44180 38344
rect 39071 38304 44180 38332
rect 39071 38301 39083 38304
rect 39025 38295 39083 38301
rect 44174 38292 44180 38304
rect 44232 38292 44238 38344
rect 46290 38332 46296 38344
rect 46251 38304 46296 38332
rect 46290 38292 46296 38304
rect 46348 38292 46354 38344
rect 40126 38264 40132 38276
rect 39224 38236 40132 38264
rect 39224 38205 39252 38236
rect 40126 38224 40132 38236
rect 40184 38264 40190 38276
rect 40221 38267 40279 38273
rect 40221 38264 40233 38267
rect 40184 38236 40233 38264
rect 40184 38224 40190 38236
rect 40221 38233 40233 38236
rect 40267 38233 40279 38267
rect 40221 38227 40279 38233
rect 46477 38267 46535 38273
rect 46477 38233 46489 38267
rect 46523 38264 46535 38267
rect 47670 38264 47676 38276
rect 46523 38236 47676 38264
rect 46523 38233 46535 38236
rect 46477 38227 46535 38233
rect 47670 38224 47676 38236
rect 47728 38224 47734 38276
rect 48130 38264 48136 38276
rect 48091 38236 48136 38264
rect 48130 38224 48136 38236
rect 48188 38224 48194 38276
rect 39209 38199 39267 38205
rect 39209 38165 39221 38199
rect 39255 38165 39267 38199
rect 39209 38159 39267 38165
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 47670 37992 47676 38004
rect 47631 37964 47676 37992
rect 47670 37952 47676 37964
rect 47728 37952 47734 38004
rect 40126 37856 40132 37868
rect 40087 37828 40132 37856
rect 40126 37816 40132 37828
rect 40184 37816 40190 37868
rect 47578 37856 47584 37868
rect 45526 37828 47584 37856
rect 20714 37748 20720 37800
rect 20772 37788 20778 37800
rect 40405 37791 40463 37797
rect 40405 37788 40417 37791
rect 20772 37760 40417 37788
rect 20772 37748 20778 37760
rect 40405 37757 40417 37760
rect 40451 37788 40463 37791
rect 45526 37788 45554 37828
rect 47578 37816 47584 37828
rect 47636 37816 47642 37868
rect 40451 37760 45554 37788
rect 40451 37757 40463 37760
rect 40405 37751 40463 37757
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 46290 37408 46296 37460
rect 46348 37448 46354 37460
rect 47673 37451 47731 37457
rect 47673 37448 47685 37451
rect 46348 37420 47685 37448
rect 46348 37408 46354 37420
rect 47673 37417 47685 37420
rect 47719 37417 47731 37451
rect 47673 37411 47731 37417
rect 1946 37204 1952 37256
rect 2004 37244 2010 37256
rect 2225 37247 2283 37253
rect 2225 37244 2237 37247
rect 2004 37216 2237 37244
rect 2004 37204 2010 37216
rect 2225 37213 2237 37216
rect 2271 37213 2283 37247
rect 2225 37207 2283 37213
rect 12434 37204 12440 37256
rect 12492 37244 12498 37256
rect 25685 37247 25743 37253
rect 25685 37244 25697 37247
rect 12492 37216 25697 37244
rect 12492 37204 12498 37216
rect 25685 37213 25697 37216
rect 25731 37213 25743 37247
rect 40126 37244 40132 37256
rect 40087 37216 40132 37244
rect 25685 37207 25743 37213
rect 40126 37204 40132 37216
rect 40184 37204 40190 37256
rect 25869 37179 25927 37185
rect 25869 37145 25881 37179
rect 25915 37176 25927 37179
rect 27522 37176 27528 37188
rect 25915 37148 27528 37176
rect 25915 37145 25927 37148
rect 25869 37139 25927 37145
rect 27522 37136 27528 37148
rect 27580 37136 27586 37188
rect 40310 37136 40316 37188
rect 40368 37176 40374 37188
rect 40497 37179 40555 37185
rect 40497 37176 40509 37179
rect 40368 37148 40509 37176
rect 40368 37136 40374 37148
rect 40497 37145 40509 37148
rect 40543 37145 40555 37179
rect 40497 37139 40555 37145
rect 25774 37068 25780 37120
rect 25832 37108 25838 37120
rect 26053 37111 26111 37117
rect 26053 37108 26065 37111
rect 25832 37080 26065 37108
rect 25832 37068 25838 37080
rect 26053 37077 26065 37080
rect 26099 37077 26111 37111
rect 26053 37071 26111 37077
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 27338 36904 27344 36916
rect 27299 36876 27344 36904
rect 27338 36864 27344 36876
rect 27396 36864 27402 36916
rect 40310 36904 40316 36916
rect 35866 36876 40316 36904
rect 25314 36796 25320 36848
rect 25372 36836 25378 36848
rect 35866 36836 35894 36876
rect 40310 36864 40316 36876
rect 40368 36904 40374 36916
rect 40678 36904 40684 36916
rect 40368 36876 40684 36904
rect 40368 36864 40374 36876
rect 40678 36864 40684 36876
rect 40736 36864 40742 36916
rect 25372 36808 35894 36836
rect 25372 36796 25378 36808
rect 1946 36768 1952 36780
rect 1907 36740 1952 36768
rect 1946 36728 1952 36740
rect 2004 36728 2010 36780
rect 23201 36771 23259 36777
rect 23201 36737 23213 36771
rect 23247 36737 23259 36771
rect 23201 36731 23259 36737
rect 2133 36703 2191 36709
rect 2133 36669 2145 36703
rect 2179 36700 2191 36703
rect 2866 36700 2872 36712
rect 2179 36672 2872 36700
rect 2179 36669 2191 36672
rect 2133 36663 2191 36669
rect 2866 36660 2872 36672
rect 2924 36660 2930 36712
rect 2958 36660 2964 36712
rect 3016 36700 3022 36712
rect 3016 36672 3061 36700
rect 3016 36660 3022 36672
rect 23216 36632 23244 36731
rect 25682 36728 25688 36780
rect 25740 36768 25746 36780
rect 26053 36771 26111 36777
rect 26053 36768 26065 36771
rect 25740 36740 26065 36768
rect 25740 36728 25746 36740
rect 26053 36737 26065 36740
rect 26099 36737 26111 36771
rect 26053 36731 26111 36737
rect 26145 36703 26203 36709
rect 26145 36669 26157 36703
rect 26191 36700 26203 36703
rect 26326 36700 26332 36712
rect 26191 36672 26332 36700
rect 26191 36669 26203 36672
rect 26145 36663 26203 36669
rect 26326 36660 26332 36672
rect 26384 36660 26390 36712
rect 26421 36703 26479 36709
rect 26421 36669 26433 36703
rect 26467 36700 26479 36703
rect 27433 36703 27491 36709
rect 27433 36700 27445 36703
rect 26467 36672 27445 36700
rect 26467 36669 26479 36672
rect 26421 36663 26479 36669
rect 27433 36669 27445 36672
rect 27479 36669 27491 36703
rect 27433 36663 27491 36669
rect 27522 36660 27528 36712
rect 27580 36700 27586 36712
rect 27580 36672 27625 36700
rect 27580 36660 27586 36672
rect 26973 36635 27031 36641
rect 26973 36632 26985 36635
rect 23216 36604 26985 36632
rect 26973 36601 26985 36604
rect 27019 36601 27031 36635
rect 26973 36595 27031 36601
rect 22370 36524 22376 36576
rect 22428 36564 22434 36576
rect 23017 36567 23075 36573
rect 23017 36564 23029 36567
rect 22428 36536 23029 36564
rect 22428 36524 22434 36536
rect 23017 36533 23029 36536
rect 23063 36533 23075 36567
rect 23017 36527 23075 36533
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 2866 36360 2872 36372
rect 2827 36332 2872 36360
rect 2866 36320 2872 36332
rect 2924 36320 2930 36372
rect 6886 36332 31754 36360
rect 2777 36159 2835 36165
rect 2777 36125 2789 36159
rect 2823 36156 2835 36159
rect 6638 36156 6644 36168
rect 2823 36128 6644 36156
rect 2823 36125 2835 36128
rect 2777 36119 2835 36125
rect 6638 36116 6644 36128
rect 6696 36156 6702 36168
rect 6886 36156 6914 36332
rect 22097 36227 22155 36233
rect 22097 36193 22109 36227
rect 22143 36224 22155 36227
rect 31726 36224 31754 36332
rect 37090 36224 37096 36236
rect 22143 36196 24440 36224
rect 31726 36196 37096 36224
rect 22143 36193 22155 36196
rect 22097 36187 22155 36193
rect 24412 36168 24440 36196
rect 37090 36184 37096 36196
rect 37148 36184 37154 36236
rect 24394 36156 24400 36168
rect 6696 36128 6914 36156
rect 24355 36128 24400 36156
rect 6696 36116 6702 36128
rect 24394 36116 24400 36128
rect 24452 36116 24458 36168
rect 28166 36116 28172 36168
rect 28224 36156 28230 36168
rect 28537 36159 28595 36165
rect 28537 36156 28549 36159
rect 28224 36128 28549 36156
rect 28224 36116 28230 36128
rect 28537 36125 28549 36128
rect 28583 36125 28595 36159
rect 33410 36156 33416 36168
rect 33371 36128 33416 36156
rect 28537 36119 28595 36125
rect 33410 36116 33416 36128
rect 33468 36116 33474 36168
rect 22370 36088 22376 36100
rect 22331 36060 22376 36088
rect 22370 36048 22376 36060
rect 22428 36048 22434 36100
rect 22830 36048 22836 36100
rect 22888 36048 22894 36100
rect 24673 36091 24731 36097
rect 24673 36057 24685 36091
rect 24719 36088 24731 36091
rect 24946 36088 24952 36100
rect 24719 36060 24952 36088
rect 24719 36057 24731 36060
rect 24673 36051 24731 36057
rect 24946 36048 24952 36060
rect 25004 36048 25010 36100
rect 25130 36048 25136 36100
rect 25188 36048 25194 36100
rect 23845 36023 23903 36029
rect 23845 35989 23857 36023
rect 23891 36020 23903 36023
rect 25682 36020 25688 36032
rect 23891 35992 25688 36020
rect 23891 35989 23903 35992
rect 23845 35983 23903 35989
rect 25682 35980 25688 35992
rect 25740 35980 25746 36032
rect 26142 36020 26148 36032
rect 26103 35992 26148 36020
rect 26142 35980 26148 35992
rect 26200 35980 26206 36032
rect 28534 35980 28540 36032
rect 28592 36020 28598 36032
rect 28629 36023 28687 36029
rect 28629 36020 28641 36023
rect 28592 35992 28641 36020
rect 28592 35980 28598 35992
rect 28629 35989 28641 35992
rect 28675 35989 28687 36023
rect 28629 35983 28687 35989
rect 33229 36023 33287 36029
rect 33229 35989 33241 36023
rect 33275 36020 33287 36023
rect 33318 36020 33324 36032
rect 33275 35992 33324 36020
rect 33275 35989 33287 35992
rect 33229 35983 33287 35989
rect 33318 35980 33324 35992
rect 33376 35980 33382 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 22649 35819 22707 35825
rect 22649 35785 22661 35819
rect 22695 35816 22707 35819
rect 22830 35816 22836 35828
rect 22695 35788 22836 35816
rect 22695 35785 22707 35788
rect 22649 35779 22707 35785
rect 22830 35776 22836 35788
rect 22888 35776 22894 35828
rect 24946 35776 24952 35828
rect 25004 35816 25010 35828
rect 25593 35819 25651 35825
rect 25593 35816 25605 35819
rect 25004 35788 25605 35816
rect 25004 35776 25010 35788
rect 25593 35785 25605 35788
rect 25639 35785 25651 35819
rect 29914 35816 29920 35828
rect 25593 35779 25651 35785
rect 25700 35788 29920 35816
rect 22370 35708 22376 35760
rect 22428 35748 22434 35760
rect 25700 35748 25728 35788
rect 29914 35776 29920 35788
rect 29972 35776 29978 35828
rect 33321 35819 33379 35825
rect 33321 35785 33333 35819
rect 33367 35816 33379 35819
rect 33410 35816 33416 35828
rect 33367 35788 33416 35816
rect 33367 35785 33379 35788
rect 33321 35779 33379 35785
rect 33410 35776 33416 35788
rect 33468 35776 33474 35828
rect 33686 35816 33692 35828
rect 33647 35788 33692 35816
rect 33686 35776 33692 35788
rect 33744 35776 33750 35828
rect 26142 35748 26148 35760
rect 22428 35720 25728 35748
rect 25977 35720 26148 35748
rect 22428 35708 22434 35720
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 22002 35640 22008 35692
rect 22060 35680 22066 35692
rect 25977 35689 26005 35720
rect 26142 35708 26148 35720
rect 26200 35708 26206 35760
rect 29270 35708 29276 35760
rect 29328 35748 29334 35760
rect 29641 35751 29699 35757
rect 29641 35748 29653 35751
rect 29328 35720 29653 35748
rect 29328 35708 29334 35720
rect 29641 35717 29653 35720
rect 29687 35717 29699 35751
rect 29641 35711 29699 35717
rect 30650 35708 30656 35760
rect 30708 35708 30714 35760
rect 22557 35683 22615 35689
rect 22557 35680 22569 35683
rect 22060 35652 22569 35680
rect 22060 35640 22066 35652
rect 22557 35649 22569 35652
rect 22603 35649 22615 35683
rect 22557 35643 22615 35649
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35649 24455 35683
rect 24397 35643 24455 35649
rect 25961 35683 26019 35689
rect 25961 35649 25973 35683
rect 26007 35649 26019 35683
rect 25961 35643 26019 35649
rect 20530 35572 20536 35624
rect 20588 35612 20594 35624
rect 24412 35612 24440 35643
rect 28534 35640 28540 35692
rect 28592 35640 28598 35692
rect 25774 35612 25780 35624
rect 20588 35584 24440 35612
rect 25735 35584 25780 35612
rect 20588 35572 20594 35584
rect 25774 35572 25780 35584
rect 25832 35572 25838 35624
rect 25869 35615 25927 35621
rect 25869 35581 25881 35615
rect 25915 35581 25927 35615
rect 25869 35575 25927 35581
rect 26053 35615 26111 35621
rect 26053 35581 26065 35615
rect 26099 35612 26111 35615
rect 26234 35612 26240 35624
rect 26099 35584 26240 35612
rect 26099 35581 26111 35584
rect 26053 35575 26111 35581
rect 25590 35504 25596 35556
rect 25648 35544 25654 35556
rect 25884 35544 25912 35575
rect 26234 35572 26240 35584
rect 26292 35572 26298 35624
rect 27154 35612 27160 35624
rect 27115 35584 27160 35612
rect 27154 35572 27160 35584
rect 27212 35572 27218 35624
rect 27433 35615 27491 35621
rect 27433 35581 27445 35615
rect 27479 35612 27491 35615
rect 28442 35612 28448 35624
rect 27479 35584 28448 35612
rect 27479 35581 27491 35584
rect 27433 35575 27491 35581
rect 28442 35572 28448 35584
rect 28500 35572 28506 35624
rect 29365 35615 29423 35621
rect 29365 35581 29377 35615
rect 29411 35612 29423 35615
rect 29411 35584 29500 35612
rect 29411 35581 29423 35584
rect 29365 35575 29423 35581
rect 25648 35516 25912 35544
rect 25648 35504 25654 35516
rect 1394 35476 1400 35488
rect 1355 35448 1400 35476
rect 1394 35436 1400 35448
rect 1452 35436 1458 35488
rect 24578 35476 24584 35488
rect 24539 35448 24584 35476
rect 24578 35436 24584 35448
rect 24636 35476 24642 35488
rect 25866 35476 25872 35488
rect 24636 35448 25872 35476
rect 24636 35436 24642 35448
rect 25866 35436 25872 35448
rect 25924 35436 25930 35488
rect 26050 35436 26056 35488
rect 26108 35476 26114 35488
rect 28166 35476 28172 35488
rect 26108 35448 28172 35476
rect 26108 35436 26114 35448
rect 28166 35436 28172 35448
rect 28224 35436 28230 35488
rect 28534 35436 28540 35488
rect 28592 35476 28598 35488
rect 28905 35479 28963 35485
rect 28905 35476 28917 35479
rect 28592 35448 28917 35476
rect 28592 35436 28598 35448
rect 28905 35445 28917 35448
rect 28951 35445 28963 35479
rect 29472 35476 29500 35584
rect 33502 35572 33508 35624
rect 33560 35612 33566 35624
rect 33781 35615 33839 35621
rect 33781 35612 33793 35615
rect 33560 35584 33793 35612
rect 33560 35572 33566 35584
rect 33781 35581 33793 35584
rect 33827 35581 33839 35615
rect 33781 35575 33839 35581
rect 33873 35615 33931 35621
rect 33873 35581 33885 35615
rect 33919 35581 33931 35615
rect 33873 35575 33931 35581
rect 33410 35504 33416 35556
rect 33468 35544 33474 35556
rect 33888 35544 33916 35575
rect 33468 35516 33916 35544
rect 33468 35504 33474 35516
rect 30374 35476 30380 35488
rect 29472 35448 30380 35476
rect 28905 35439 28963 35445
rect 30374 35436 30380 35448
rect 30432 35436 30438 35488
rect 30834 35436 30840 35488
rect 30892 35476 30898 35488
rect 31113 35479 31171 35485
rect 31113 35476 31125 35479
rect 30892 35448 31125 35476
rect 30892 35436 30898 35448
rect 31113 35445 31125 35448
rect 31159 35445 31171 35479
rect 31113 35439 31171 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 24765 35275 24823 35281
rect 24765 35241 24777 35275
rect 24811 35272 24823 35275
rect 25130 35272 25136 35284
rect 24811 35244 25136 35272
rect 24811 35241 24823 35244
rect 24765 35235 24823 35241
rect 25130 35232 25136 35244
rect 25188 35232 25194 35284
rect 26053 35275 26111 35281
rect 26053 35241 26065 35275
rect 26099 35272 26111 35275
rect 26234 35272 26240 35284
rect 26099 35244 26240 35272
rect 26099 35241 26111 35244
rect 26053 35235 26111 35241
rect 26234 35232 26240 35244
rect 26292 35232 26298 35284
rect 26326 35232 26332 35284
rect 26384 35272 26390 35284
rect 26421 35275 26479 35281
rect 26421 35272 26433 35275
rect 26384 35244 26433 35272
rect 26384 35232 26390 35244
rect 26421 35241 26433 35244
rect 26467 35241 26479 35275
rect 26421 35235 26479 35241
rect 27157 35275 27215 35281
rect 27157 35241 27169 35275
rect 27203 35272 27215 35275
rect 27246 35272 27252 35284
rect 27203 35244 27252 35272
rect 27203 35241 27215 35244
rect 27157 35235 27215 35241
rect 26436 35204 26464 35235
rect 27246 35232 27252 35244
rect 27304 35232 27310 35284
rect 28074 35272 28080 35284
rect 28035 35244 28080 35272
rect 28074 35232 28080 35244
rect 28132 35232 28138 35284
rect 30469 35275 30527 35281
rect 30469 35241 30481 35275
rect 30515 35272 30527 35275
rect 30650 35272 30656 35284
rect 30515 35244 30656 35272
rect 30515 35241 30527 35244
rect 30469 35235 30527 35241
rect 30650 35232 30656 35244
rect 30708 35232 30714 35284
rect 33502 35272 33508 35284
rect 33463 35244 33508 35272
rect 33502 35232 33508 35244
rect 33560 35232 33566 35284
rect 27341 35207 27399 35213
rect 27341 35204 27353 35207
rect 26436 35176 27353 35204
rect 27341 35173 27353 35176
rect 27387 35173 27399 35207
rect 27341 35167 27399 35173
rect 25593 35139 25651 35145
rect 25593 35105 25605 35139
rect 25639 35136 25651 35139
rect 25958 35136 25964 35148
rect 25639 35108 25964 35136
rect 25639 35105 25651 35108
rect 25593 35099 25651 35105
rect 25958 35096 25964 35108
rect 26016 35136 26022 35148
rect 26142 35136 26148 35148
rect 26016 35108 26148 35136
rect 26016 35096 26022 35108
rect 26142 35096 26148 35108
rect 26200 35096 26206 35148
rect 28092 35136 28120 35232
rect 26344 35108 28120 35136
rect 20254 35028 20260 35080
rect 20312 35068 20318 35080
rect 20530 35068 20536 35080
rect 20312 35040 20536 35068
rect 20312 35028 20318 35040
rect 20530 35028 20536 35040
rect 20588 35028 20594 35080
rect 24578 35028 24584 35080
rect 24636 35068 24642 35080
rect 24673 35071 24731 35077
rect 24673 35068 24685 35071
rect 24636 35040 24685 35068
rect 24636 35028 24642 35040
rect 24673 35037 24685 35040
rect 24719 35037 24731 35071
rect 25314 35068 25320 35080
rect 25275 35040 25320 35068
rect 24673 35031 24731 35037
rect 25314 35028 25320 35040
rect 25372 35028 25378 35080
rect 25406 35028 25412 35080
rect 25464 35068 25470 35080
rect 25464 35040 25509 35068
rect 25464 35028 25470 35040
rect 25774 35028 25780 35080
rect 25832 35068 25838 35080
rect 26237 35071 26295 35077
rect 26237 35068 26249 35071
rect 25832 35040 26249 35068
rect 25832 35028 25838 35040
rect 26237 35037 26249 35040
rect 26283 35037 26295 35071
rect 26237 35031 26295 35037
rect 25130 34960 25136 35012
rect 25188 35000 25194 35012
rect 26344 35000 26372 35108
rect 31110 35096 31116 35148
rect 31168 35136 31174 35148
rect 33045 35139 33103 35145
rect 33045 35136 33057 35139
rect 31168 35108 33057 35136
rect 31168 35096 31174 35108
rect 33045 35105 33057 35108
rect 33091 35105 33103 35139
rect 33045 35099 33103 35105
rect 26513 35071 26571 35077
rect 26513 35037 26525 35071
rect 26559 35068 26571 35071
rect 28166 35068 28172 35080
rect 26559 35040 28172 35068
rect 26559 35037 26571 35040
rect 26513 35031 26571 35037
rect 28166 35028 28172 35040
rect 28224 35028 28230 35080
rect 28258 35028 28264 35080
rect 28316 35068 28322 35080
rect 30377 35071 30435 35077
rect 30377 35068 30389 35071
rect 28316 35040 30389 35068
rect 28316 35028 28322 35040
rect 30377 35037 30389 35040
rect 30423 35068 30435 35071
rect 31021 35071 31079 35077
rect 31021 35068 31033 35071
rect 30423 35040 31033 35068
rect 30423 35037 30435 35040
rect 30377 35031 30435 35037
rect 31021 35037 31033 35040
rect 31067 35037 31079 35071
rect 31021 35031 31079 35037
rect 33137 35071 33195 35077
rect 33137 35037 33149 35071
rect 33183 35068 33195 35071
rect 34606 35068 34612 35080
rect 33183 35040 34612 35068
rect 33183 35037 33195 35040
rect 33137 35031 33195 35037
rect 34606 35028 34612 35040
rect 34664 35028 34670 35080
rect 48130 35068 48136 35080
rect 48091 35040 48136 35068
rect 48130 35028 48136 35040
rect 48188 35028 48194 35080
rect 25188 34972 26372 35000
rect 26973 35003 27031 35009
rect 25188 34960 25194 34972
rect 26973 34969 26985 35003
rect 27019 35000 27031 35003
rect 27614 35000 27620 35012
rect 27019 34972 27620 35000
rect 27019 34969 27031 34972
rect 26973 34963 27031 34969
rect 27614 34960 27620 34972
rect 27672 34960 27678 35012
rect 27985 35003 28043 35009
rect 27985 34969 27997 35003
rect 28031 34969 28043 35003
rect 27985 34963 28043 34969
rect 20717 34935 20775 34941
rect 20717 34901 20729 34935
rect 20763 34932 20775 34935
rect 20806 34932 20812 34944
rect 20763 34904 20812 34932
rect 20763 34901 20775 34904
rect 20717 34895 20775 34901
rect 20806 34892 20812 34904
rect 20864 34892 20870 34944
rect 25317 34935 25375 34941
rect 25317 34901 25329 34935
rect 25363 34932 25375 34935
rect 27173 34935 27231 34941
rect 27173 34932 27185 34935
rect 25363 34904 27185 34932
rect 25363 34901 25375 34904
rect 25317 34895 25375 34901
rect 27173 34901 27185 34904
rect 27219 34901 27231 34935
rect 27173 34895 27231 34901
rect 27338 34892 27344 34944
rect 27396 34932 27402 34944
rect 28000 34932 28028 34963
rect 27396 34904 28028 34932
rect 31113 34935 31171 34941
rect 27396 34892 27402 34904
rect 31113 34901 31125 34935
rect 31159 34932 31171 34935
rect 31754 34932 31760 34944
rect 31159 34904 31760 34932
rect 31159 34901 31171 34904
rect 31113 34895 31171 34901
rect 31754 34892 31760 34904
rect 31812 34892 31818 34944
rect 47118 34892 47124 34944
rect 47176 34932 47182 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47176 34904 47961 34932
rect 47176 34892 47182 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 25682 34688 25688 34740
rect 25740 34688 25746 34740
rect 28994 34728 29000 34740
rect 28955 34700 29000 34728
rect 28994 34688 29000 34700
rect 29052 34688 29058 34740
rect 29270 34728 29276 34740
rect 29231 34700 29276 34728
rect 29270 34688 29276 34700
rect 29328 34688 29334 34740
rect 29454 34728 29460 34740
rect 29415 34700 29460 34728
rect 29454 34688 29460 34700
rect 29512 34688 29518 34740
rect 31110 34728 31116 34740
rect 31071 34700 31116 34728
rect 31110 34688 31116 34700
rect 31168 34688 31174 34740
rect 25700 34660 25728 34688
rect 29012 34660 29040 34688
rect 30745 34663 30803 34669
rect 25700 34632 26004 34660
rect 29012 34632 29868 34660
rect 20806 34552 20812 34604
rect 20864 34592 20870 34604
rect 22002 34592 22008 34604
rect 20864 34564 22008 34592
rect 20864 34552 20870 34564
rect 22002 34552 22008 34564
rect 22060 34592 22066 34604
rect 22097 34595 22155 34601
rect 22097 34592 22109 34595
rect 22060 34564 22109 34592
rect 22060 34552 22066 34564
rect 22097 34561 22109 34564
rect 22143 34561 22155 34595
rect 22097 34555 22155 34561
rect 24854 34552 24860 34604
rect 24912 34552 24918 34604
rect 25976 34601 26004 34632
rect 25685 34595 25743 34601
rect 25685 34592 25697 34595
rect 25240 34564 25697 34592
rect 25240 34536 25268 34564
rect 25685 34561 25697 34564
rect 25731 34561 25743 34595
rect 25685 34555 25743 34561
rect 25961 34595 26019 34601
rect 25961 34561 25973 34595
rect 26007 34561 26019 34595
rect 25961 34555 26019 34561
rect 29454 34595 29512 34601
rect 29454 34561 29466 34595
rect 29500 34592 29512 34595
rect 29546 34592 29552 34604
rect 29500 34564 29552 34592
rect 29500 34561 29512 34564
rect 29454 34555 29512 34561
rect 29546 34552 29552 34564
rect 29604 34552 29610 34604
rect 29840 34601 29868 34632
rect 30745 34629 30757 34663
rect 30791 34629 30803 34663
rect 30745 34623 30803 34629
rect 30961 34663 31019 34669
rect 30961 34629 30973 34663
rect 31007 34660 31019 34663
rect 31294 34660 31300 34672
rect 31007 34632 31300 34660
rect 31007 34629 31019 34632
rect 30961 34623 31019 34629
rect 29825 34595 29883 34601
rect 29825 34561 29837 34595
rect 29871 34561 29883 34595
rect 29825 34555 29883 34561
rect 29914 34552 29920 34604
rect 29972 34592 29978 34604
rect 29972 34564 30017 34592
rect 29972 34552 29978 34564
rect 22186 34524 22192 34536
rect 22147 34496 22192 34524
rect 22186 34484 22192 34496
rect 22244 34484 22250 34536
rect 23474 34524 23480 34536
rect 23435 34496 23480 34524
rect 23474 34484 23480 34496
rect 23532 34484 23538 34536
rect 23750 34524 23756 34536
rect 23711 34496 23756 34524
rect 23750 34484 23756 34496
rect 23808 34484 23814 34536
rect 25222 34524 25228 34536
rect 25183 34496 25228 34524
rect 25222 34484 25228 34496
rect 25280 34484 25286 34536
rect 25406 34484 25412 34536
rect 25464 34524 25470 34536
rect 25774 34524 25780 34536
rect 25464 34496 25780 34524
rect 25464 34484 25470 34496
rect 25774 34484 25780 34496
rect 25832 34484 25838 34536
rect 27614 34484 27620 34536
rect 27672 34524 27678 34536
rect 28074 34524 28080 34536
rect 27672 34496 28080 34524
rect 27672 34484 27678 34496
rect 28074 34484 28080 34496
rect 28132 34524 28138 34536
rect 30760 34524 30788 34623
rect 31294 34620 31300 34632
rect 31352 34620 31358 34672
rect 33318 34660 33324 34672
rect 33279 34632 33324 34660
rect 33318 34620 33324 34632
rect 33376 34620 33382 34672
rect 34790 34660 34796 34672
rect 34546 34632 34796 34660
rect 34790 34620 34796 34632
rect 34848 34620 34854 34672
rect 48130 34592 48136 34604
rect 48091 34564 48136 34592
rect 48130 34552 48136 34564
rect 48188 34552 48194 34604
rect 28132 34496 30788 34524
rect 28132 34484 28138 34496
rect 31662 34484 31668 34536
rect 31720 34524 31726 34536
rect 33045 34527 33103 34533
rect 33045 34524 33057 34527
rect 31720 34496 33057 34524
rect 31720 34484 31726 34496
rect 33045 34493 33057 34496
rect 33091 34493 33103 34527
rect 33045 34487 33103 34493
rect 34606 34484 34612 34536
rect 34664 34524 34670 34536
rect 34793 34527 34851 34533
rect 34793 34524 34805 34527
rect 34664 34496 34805 34524
rect 34664 34484 34670 34496
rect 34793 34493 34805 34496
rect 34839 34493 34851 34527
rect 34793 34487 34851 34493
rect 27154 34456 27160 34468
rect 25792 34428 27160 34456
rect 23474 34348 23480 34400
rect 23532 34388 23538 34400
rect 24394 34388 24400 34400
rect 23532 34360 24400 34388
rect 23532 34348 23538 34360
rect 24394 34348 24400 34360
rect 24452 34388 24458 34400
rect 25792 34388 25820 34428
rect 27154 34416 27160 34428
rect 27212 34416 27218 34468
rect 25958 34388 25964 34400
rect 24452 34360 25820 34388
rect 25919 34360 25964 34388
rect 24452 34348 24458 34360
rect 25958 34348 25964 34360
rect 26016 34348 26022 34400
rect 26142 34388 26148 34400
rect 26103 34360 26148 34388
rect 26142 34348 26148 34360
rect 26200 34348 26206 34400
rect 27246 34348 27252 34400
rect 27304 34388 27310 34400
rect 30929 34391 30987 34397
rect 30929 34388 30941 34391
rect 27304 34360 30941 34388
rect 27304 34348 27310 34360
rect 30929 34357 30941 34360
rect 30975 34357 30987 34391
rect 30929 34351 30987 34357
rect 47854 34348 47860 34400
rect 47912 34388 47918 34400
rect 47949 34391 48007 34397
rect 47949 34388 47961 34391
rect 47912 34360 47961 34388
rect 47912 34348 47918 34360
rect 47949 34357 47961 34360
rect 47995 34357 48007 34391
rect 47949 34351 48007 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 24673 34187 24731 34193
rect 24673 34153 24685 34187
rect 24719 34184 24731 34187
rect 24854 34184 24860 34196
rect 24719 34156 24860 34184
rect 24719 34153 24731 34156
rect 24673 34147 24731 34153
rect 24854 34144 24860 34156
rect 24912 34144 24918 34196
rect 26050 34184 26056 34196
rect 26011 34156 26056 34184
rect 26050 34144 26056 34156
rect 26108 34144 26114 34196
rect 29546 34144 29552 34196
rect 29604 34184 29610 34196
rect 29917 34187 29975 34193
rect 29917 34184 29929 34187
rect 29604 34156 29929 34184
rect 29604 34144 29610 34156
rect 29917 34153 29929 34156
rect 29963 34153 29975 34187
rect 30926 34184 30932 34196
rect 29917 34147 29975 34153
rect 30024 34156 30932 34184
rect 25590 34076 25596 34128
rect 25648 34116 25654 34128
rect 26237 34119 26295 34125
rect 26237 34116 26249 34119
rect 25648 34088 26249 34116
rect 25648 34076 25654 34088
rect 26237 34085 26249 34088
rect 26283 34085 26295 34119
rect 26237 34079 26295 34085
rect 28626 34076 28632 34128
rect 28684 34116 28690 34128
rect 30024 34116 30052 34156
rect 30926 34144 30932 34156
rect 30984 34144 30990 34196
rect 34790 34184 34796 34196
rect 34751 34156 34796 34184
rect 34790 34144 34796 34156
rect 34848 34144 34854 34196
rect 28684 34088 30052 34116
rect 28684 34076 28690 34088
rect 20070 34008 20076 34060
rect 20128 34048 20134 34060
rect 21361 34051 21419 34057
rect 21361 34048 21373 34051
rect 20128 34020 21373 34048
rect 20128 34008 20134 34020
rect 21361 34017 21373 34020
rect 21407 34048 21419 34051
rect 23474 34048 23480 34060
rect 21407 34020 23480 34048
rect 21407 34017 21419 34020
rect 21361 34011 21419 34017
rect 23474 34008 23480 34020
rect 23532 34008 23538 34060
rect 25774 34008 25780 34060
rect 25832 34048 25838 34060
rect 25961 34051 26019 34057
rect 25961 34048 25973 34051
rect 25832 34020 25973 34048
rect 25832 34008 25838 34020
rect 25961 34017 25973 34020
rect 26007 34017 26019 34051
rect 25961 34011 26019 34017
rect 28445 34051 28503 34057
rect 28445 34017 28457 34051
rect 28491 34048 28503 34051
rect 29086 34048 29092 34060
rect 28491 34020 29092 34048
rect 28491 34017 28503 34020
rect 28445 34011 28503 34017
rect 29086 34008 29092 34020
rect 29144 34008 29150 34060
rect 30374 34008 30380 34060
rect 30432 34048 30438 34060
rect 30469 34051 30527 34057
rect 30469 34048 30481 34051
rect 30432 34020 30481 34048
rect 30432 34008 30438 34020
rect 30469 34017 30481 34020
rect 30515 34048 30527 34051
rect 31478 34048 31484 34060
rect 30515 34020 31484 34048
rect 30515 34017 30527 34020
rect 30469 34011 30527 34017
rect 31478 34008 31484 34020
rect 31536 34008 31542 34060
rect 20533 33983 20591 33989
rect 20533 33949 20545 33983
rect 20579 33980 20591 33983
rect 20806 33980 20812 33992
rect 20579 33952 20812 33980
rect 20579 33949 20591 33952
rect 20533 33943 20591 33949
rect 20806 33940 20812 33952
rect 20864 33940 20870 33992
rect 24578 33980 24584 33992
rect 24539 33952 24584 33980
rect 24578 33940 24584 33952
rect 24636 33940 24642 33992
rect 25314 33940 25320 33992
rect 25372 33980 25378 33992
rect 25866 33980 25872 33992
rect 25372 33952 25872 33980
rect 25372 33940 25378 33952
rect 25866 33940 25872 33952
rect 25924 33940 25930 33992
rect 28166 33980 28172 33992
rect 28127 33952 28172 33980
rect 28166 33940 28172 33952
rect 28224 33940 28230 33992
rect 28261 33983 28319 33989
rect 28261 33949 28273 33983
rect 28307 33980 28319 33983
rect 28810 33980 28816 33992
rect 28307 33952 28816 33980
rect 28307 33949 28319 33952
rect 28261 33943 28319 33949
rect 28810 33940 28816 33952
rect 28868 33940 28874 33992
rect 29825 33983 29883 33989
rect 29825 33949 29837 33983
rect 29871 33949 29883 33983
rect 29825 33943 29883 33949
rect 30009 33983 30067 33989
rect 30009 33949 30021 33983
rect 30055 33980 30067 33983
rect 34701 33983 34759 33989
rect 30055 33952 30512 33980
rect 30055 33949 30067 33952
rect 30009 33943 30067 33949
rect 21634 33912 21640 33924
rect 21595 33884 21640 33912
rect 21634 33872 21640 33884
rect 21692 33872 21698 33924
rect 22186 33872 22192 33924
rect 22244 33872 22250 33924
rect 24762 33872 24768 33924
rect 24820 33912 24826 33924
rect 28445 33915 28503 33921
rect 28445 33912 28457 33915
rect 24820 33884 28457 33912
rect 24820 33872 24826 33884
rect 28445 33881 28457 33884
rect 28491 33881 28503 33915
rect 29840 33912 29868 33943
rect 30374 33912 30380 33924
rect 29840 33884 30380 33912
rect 28445 33875 28503 33881
rect 30374 33872 30380 33884
rect 30432 33872 30438 33924
rect 20530 33804 20536 33856
rect 20588 33844 20594 33856
rect 20625 33847 20683 33853
rect 20625 33844 20637 33847
rect 20588 33816 20637 33844
rect 20588 33804 20594 33816
rect 20625 33813 20637 33816
rect 20671 33813 20683 33847
rect 20625 33807 20683 33813
rect 23109 33847 23167 33853
rect 23109 33813 23121 33847
rect 23155 33844 23167 33847
rect 23566 33844 23572 33856
rect 23155 33816 23572 33844
rect 23155 33813 23167 33816
rect 23109 33807 23167 33813
rect 23566 33804 23572 33816
rect 23624 33844 23630 33856
rect 24670 33844 24676 33856
rect 23624 33816 24676 33844
rect 23624 33804 23630 33816
rect 24670 33804 24676 33816
rect 24728 33804 24734 33856
rect 30484 33844 30512 33952
rect 34701 33949 34713 33983
rect 34747 33980 34759 33983
rect 35342 33980 35348 33992
rect 34747 33952 35348 33980
rect 34747 33949 34759 33952
rect 34701 33943 34759 33949
rect 35342 33940 35348 33952
rect 35400 33940 35406 33992
rect 47857 33983 47915 33989
rect 47857 33949 47869 33983
rect 47903 33980 47915 33983
rect 47946 33980 47952 33992
rect 47903 33952 47952 33980
rect 47903 33949 47915 33952
rect 47857 33943 47915 33949
rect 47946 33940 47952 33952
rect 48004 33940 48010 33992
rect 30742 33912 30748 33924
rect 30703 33884 30748 33912
rect 30742 33872 30748 33884
rect 30800 33872 30806 33924
rect 31754 33872 31760 33924
rect 31812 33872 31818 33924
rect 32674 33912 32680 33924
rect 32048 33884 32680 33912
rect 30834 33844 30840 33856
rect 30484 33816 30840 33844
rect 30834 33804 30840 33816
rect 30892 33804 30898 33856
rect 30926 33804 30932 33856
rect 30984 33844 30990 33856
rect 32048 33844 32076 33884
rect 32674 33872 32680 33884
rect 32732 33872 32738 33924
rect 32214 33844 32220 33856
rect 30984 33816 32076 33844
rect 32175 33816 32220 33844
rect 30984 33804 30990 33816
rect 32214 33804 32220 33816
rect 32272 33804 32278 33856
rect 48038 33844 48044 33856
rect 47999 33816 48044 33844
rect 48038 33804 48044 33816
rect 48096 33804 48102 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 21634 33600 21640 33652
rect 21692 33640 21698 33652
rect 22557 33643 22615 33649
rect 22557 33640 22569 33643
rect 21692 33612 22569 33640
rect 21692 33600 21698 33612
rect 22557 33609 22569 33612
rect 22603 33609 22615 33643
rect 22557 33603 22615 33609
rect 23750 33600 23756 33652
rect 23808 33640 23814 33652
rect 24949 33643 25007 33649
rect 24949 33640 24961 33643
rect 23808 33612 24961 33640
rect 23808 33600 23814 33612
rect 24949 33609 24961 33612
rect 24995 33609 25007 33643
rect 28442 33640 28448 33652
rect 28403 33612 28448 33640
rect 24949 33603 25007 33609
rect 28442 33600 28448 33612
rect 28500 33600 28506 33652
rect 29273 33643 29331 33649
rect 29273 33609 29285 33643
rect 29319 33640 29331 33643
rect 29454 33640 29460 33652
rect 29319 33612 29460 33640
rect 29319 33609 29331 33612
rect 29273 33603 29331 33609
rect 29454 33600 29460 33612
rect 29512 33600 29518 33652
rect 32585 33643 32643 33649
rect 32585 33640 32597 33643
rect 29564 33612 32597 33640
rect 15838 33572 15844 33584
rect 15799 33544 15844 33572
rect 15838 33532 15844 33544
rect 15896 33532 15902 33584
rect 20070 33572 20076 33584
rect 19536 33544 20076 33572
rect 1394 33464 1400 33516
rect 1452 33504 1458 33516
rect 19536 33513 19564 33544
rect 20070 33532 20076 33544
rect 20128 33532 20134 33584
rect 20530 33532 20536 33584
rect 20588 33532 20594 33584
rect 22186 33572 22192 33584
rect 21836 33544 22192 33572
rect 21836 33513 21864 33544
rect 22186 33532 22192 33544
rect 22244 33532 22250 33584
rect 23566 33572 23572 33584
rect 22296 33544 23572 33572
rect 1949 33507 2007 33513
rect 1949 33504 1961 33507
rect 1452 33476 1961 33504
rect 1452 33464 1458 33476
rect 1949 33473 1961 33476
rect 1995 33473 2007 33507
rect 1949 33467 2007 33473
rect 19521 33507 19579 33513
rect 19521 33473 19533 33507
rect 19567 33473 19579 33507
rect 19521 33467 19579 33473
rect 21821 33507 21879 33513
rect 21821 33473 21833 33507
rect 21867 33473 21879 33507
rect 21821 33467 21879 33473
rect 21910 33464 21916 33516
rect 21968 33504 21974 33516
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 21968 33476 22017 33504
rect 21968 33464 21974 33476
rect 22005 33473 22017 33476
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 22097 33507 22155 33513
rect 22097 33473 22109 33507
rect 22143 33504 22155 33507
rect 22296 33504 22324 33544
rect 23566 33532 23572 33544
rect 23624 33532 23630 33584
rect 25593 33575 25651 33581
rect 25593 33541 25605 33575
rect 25639 33572 25651 33575
rect 26142 33572 26148 33584
rect 25639 33544 26148 33572
rect 25639 33541 25651 33544
rect 25593 33535 25651 33541
rect 26142 33532 26148 33544
rect 26200 33532 26206 33584
rect 28718 33572 28724 33584
rect 27540 33544 28724 33572
rect 22143 33476 22324 33504
rect 22143 33473 22155 33476
rect 22097 33467 22155 33473
rect 22370 33464 22376 33516
rect 22428 33504 22434 33516
rect 22830 33504 22836 33516
rect 22428 33476 22836 33504
rect 22428 33464 22434 33476
rect 22830 33464 22836 33476
rect 22888 33464 22894 33516
rect 24762 33504 24768 33516
rect 24723 33476 24768 33504
rect 24762 33464 24768 33476
rect 24820 33464 24826 33516
rect 25682 33464 25688 33516
rect 25740 33504 25746 33516
rect 25777 33507 25835 33513
rect 25777 33504 25789 33507
rect 25740 33476 25789 33504
rect 25740 33464 25746 33476
rect 25777 33473 25789 33476
rect 25823 33504 25835 33507
rect 27540 33504 27568 33544
rect 28718 33532 28724 33544
rect 28776 33572 28782 33584
rect 29564 33572 29592 33612
rect 32585 33609 32597 33612
rect 32631 33609 32643 33643
rect 32585 33603 32643 33609
rect 32674 33600 32680 33652
rect 32732 33640 32738 33652
rect 48038 33640 48044 33652
rect 32732 33612 48044 33640
rect 32732 33600 32738 33612
rect 48038 33600 48044 33612
rect 48096 33600 48102 33652
rect 28776 33544 29592 33572
rect 29825 33575 29883 33581
rect 28776 33532 28782 33544
rect 29825 33541 29837 33575
rect 29871 33572 29883 33575
rect 30098 33572 30104 33584
rect 29871 33544 30104 33572
rect 29871 33541 29883 33544
rect 29825 33535 29883 33541
rect 30098 33532 30104 33544
rect 30156 33572 30162 33584
rect 30745 33575 30803 33581
rect 30745 33572 30757 33575
rect 30156 33544 30757 33572
rect 30156 33532 30162 33544
rect 30745 33541 30757 33544
rect 30791 33541 30803 33575
rect 30745 33535 30803 33541
rect 32125 33575 32183 33581
rect 32125 33541 32137 33575
rect 32171 33572 32183 33575
rect 32171 33544 32536 33572
rect 32171 33541 32183 33544
rect 32125 33535 32183 33541
rect 32508 33516 32536 33544
rect 46106 33532 46112 33584
rect 46164 33572 46170 33584
rect 46164 33544 47624 33572
rect 46164 33532 46170 33544
rect 27706 33504 27712 33516
rect 25823 33476 27568 33504
rect 27667 33476 27712 33504
rect 25823 33473 25835 33476
rect 25777 33467 25835 33473
rect 27706 33464 27712 33476
rect 27764 33464 27770 33516
rect 27893 33507 27951 33513
rect 27893 33504 27905 33507
rect 27816 33476 27905 33504
rect 2133 33439 2191 33445
rect 2133 33405 2145 33439
rect 2179 33436 2191 33439
rect 3694 33436 3700 33448
rect 2179 33408 3700 33436
rect 2179 33405 2191 33408
rect 2133 33399 2191 33405
rect 3694 33396 3700 33408
rect 3752 33396 3758 33448
rect 3789 33439 3847 33445
rect 3789 33405 3801 33439
rect 3835 33436 3847 33439
rect 4614 33436 4620 33448
rect 3835 33408 4620 33436
rect 3835 33405 3847 33408
rect 3789 33399 3847 33405
rect 4614 33396 4620 33408
rect 4672 33396 4678 33448
rect 13354 33396 13360 33448
rect 13412 33436 13418 33448
rect 14001 33439 14059 33445
rect 14001 33436 14013 33439
rect 13412 33408 14013 33436
rect 13412 33396 13418 33408
rect 14001 33405 14013 33408
rect 14047 33405 14059 33439
rect 14182 33436 14188 33448
rect 14143 33408 14188 33436
rect 14001 33399 14059 33405
rect 14182 33396 14188 33408
rect 14240 33396 14246 33448
rect 19797 33439 19855 33445
rect 19797 33405 19809 33439
rect 19843 33436 19855 33439
rect 20990 33436 20996 33448
rect 19843 33408 20996 33436
rect 19843 33405 19855 33408
rect 19797 33399 19855 33405
rect 20990 33396 20996 33408
rect 21048 33396 21054 33448
rect 22189 33439 22247 33445
rect 22189 33405 22201 33439
rect 22235 33405 22247 33439
rect 22189 33399 22247 33405
rect 22204 33368 22232 33399
rect 24118 33396 24124 33448
rect 24176 33436 24182 33448
rect 24305 33439 24363 33445
rect 24305 33436 24317 33439
rect 24176 33408 24317 33436
rect 24176 33396 24182 33408
rect 24305 33405 24317 33408
rect 24351 33405 24363 33439
rect 24305 33399 24363 33405
rect 24673 33439 24731 33445
rect 24673 33405 24685 33439
rect 24719 33436 24731 33439
rect 25222 33436 25228 33448
rect 24719 33408 25228 33436
rect 24719 33405 24731 33408
rect 24673 33399 24731 33405
rect 25222 33396 25228 33408
rect 25280 33396 25286 33448
rect 27816 33436 27844 33476
rect 27893 33473 27905 33476
rect 27939 33473 27951 33507
rect 28258 33504 28264 33516
rect 28219 33476 28264 33504
rect 27893 33467 27951 33473
rect 28258 33464 28264 33476
rect 28316 33464 28322 33516
rect 29086 33464 29092 33516
rect 29144 33504 29150 33516
rect 29549 33507 29607 33513
rect 29549 33504 29561 33507
rect 29144 33476 29561 33504
rect 29144 33464 29150 33476
rect 29549 33473 29561 33476
rect 29595 33473 29607 33507
rect 30374 33504 30380 33516
rect 29549 33467 29607 33473
rect 29840 33476 30236 33504
rect 30335 33476 30380 33504
rect 27982 33436 27988 33448
rect 25332 33408 27844 33436
rect 27943 33408 27988 33436
rect 20824 33340 22232 33368
rect 16942 33260 16948 33312
rect 17000 33300 17006 33312
rect 20824 33300 20852 33340
rect 22370 33328 22376 33380
rect 22428 33368 22434 33380
rect 25332 33368 25360 33408
rect 22428 33340 25360 33368
rect 22428 33328 22434 33340
rect 25406 33328 25412 33380
rect 25464 33368 25470 33380
rect 27816 33368 27844 33408
rect 27982 33396 27988 33408
rect 28040 33396 28046 33448
rect 28077 33439 28135 33445
rect 28077 33405 28089 33439
rect 28123 33436 28135 33439
rect 28350 33436 28356 33448
rect 28123 33408 28356 33436
rect 28123 33405 28135 33408
rect 28077 33399 28135 33405
rect 28350 33396 28356 33408
rect 28408 33396 28414 33448
rect 29457 33439 29515 33445
rect 29457 33405 29469 33439
rect 29503 33436 29515 33439
rect 29840 33436 29868 33476
rect 29503 33408 29868 33436
rect 29917 33439 29975 33445
rect 29503 33405 29515 33408
rect 29457 33399 29515 33405
rect 29917 33405 29929 33439
rect 29963 33405 29975 33439
rect 30208 33436 30236 33476
rect 30374 33464 30380 33476
rect 30432 33464 30438 33516
rect 30561 33507 30619 33513
rect 30561 33473 30573 33507
rect 30607 33504 30619 33507
rect 30834 33504 30840 33516
rect 30607 33476 30840 33504
rect 30607 33473 30619 33476
rect 30561 33467 30619 33473
rect 30576 33436 30604 33467
rect 30834 33464 30840 33476
rect 30892 33464 30898 33516
rect 30926 33464 30932 33516
rect 30984 33504 30990 33516
rect 32214 33504 32220 33516
rect 30984 33476 32220 33504
rect 30984 33464 30990 33476
rect 32214 33464 32220 33476
rect 32272 33504 32278 33516
rect 32401 33507 32459 33513
rect 32401 33504 32413 33507
rect 32272 33476 32413 33504
rect 32272 33464 32278 33476
rect 32401 33473 32413 33476
rect 32447 33473 32459 33507
rect 32401 33467 32459 33473
rect 32490 33464 32496 33516
rect 32548 33504 32554 33516
rect 33045 33507 33103 33513
rect 33045 33504 33057 33507
rect 32548 33476 33057 33504
rect 32548 33464 32554 33476
rect 33045 33473 33057 33476
rect 33091 33473 33103 33507
rect 35342 33504 35348 33516
rect 35303 33476 35348 33504
rect 33045 33467 33103 33473
rect 35342 33464 35348 33476
rect 35400 33464 35406 33516
rect 47596 33513 47624 33544
rect 47029 33507 47087 33513
rect 47029 33473 47041 33507
rect 47075 33473 47087 33507
rect 47029 33467 47087 33473
rect 47581 33507 47639 33513
rect 47581 33473 47593 33507
rect 47627 33473 47639 33507
rect 47581 33467 47639 33473
rect 30208 33408 30604 33436
rect 32309 33439 32367 33445
rect 29917 33399 29975 33405
rect 32309 33405 32321 33439
rect 32355 33436 32367 33439
rect 33321 33439 33379 33445
rect 33321 33436 33333 33439
rect 32355 33408 33333 33436
rect 32355 33405 32367 33408
rect 32309 33399 32367 33405
rect 28442 33368 28448 33380
rect 25464 33340 26096 33368
rect 27816 33340 28448 33368
rect 25464 33328 25470 33340
rect 17000 33272 20852 33300
rect 17000 33260 17006 33272
rect 21082 33260 21088 33312
rect 21140 33300 21146 33312
rect 21269 33303 21327 33309
rect 21269 33300 21281 33303
rect 21140 33272 21281 33300
rect 21140 33260 21146 33272
rect 21269 33269 21281 33272
rect 21315 33269 21327 33303
rect 21269 33263 21327 33269
rect 22186 33260 22192 33312
rect 22244 33300 22250 33312
rect 22922 33300 22928 33312
rect 22244 33272 22928 33300
rect 22244 33260 22250 33272
rect 22922 33260 22928 33272
rect 22980 33260 22986 33312
rect 25038 33260 25044 33312
rect 25096 33300 25102 33312
rect 25961 33303 26019 33309
rect 25961 33300 25973 33303
rect 25096 33272 25973 33300
rect 25096 33260 25102 33272
rect 25961 33269 25973 33272
rect 26007 33269 26019 33303
rect 26068 33300 26096 33340
rect 28442 33328 28448 33340
rect 28500 33328 28506 33380
rect 29932 33300 29960 33399
rect 33060 33380 33088 33408
rect 33321 33405 33333 33408
rect 33367 33405 33379 33439
rect 47044 33436 47072 33467
rect 48041 33439 48099 33445
rect 48041 33436 48053 33439
rect 47044 33408 48053 33436
rect 33321 33399 33379 33405
rect 48041 33405 48053 33408
rect 48087 33405 48099 33439
rect 48041 33399 48099 33405
rect 33042 33328 33048 33380
rect 33100 33328 33106 33380
rect 26068 33272 29960 33300
rect 25961 33263 26019 33269
rect 30834 33260 30840 33312
rect 30892 33300 30898 33312
rect 32125 33303 32183 33309
rect 32125 33300 32137 33303
rect 30892 33272 32137 33300
rect 30892 33260 30898 33272
rect 32125 33269 32137 33272
rect 32171 33269 32183 33303
rect 33134 33300 33140 33312
rect 33095 33272 33140 33300
rect 32125 33263 32183 33269
rect 33134 33260 33140 33272
rect 33192 33260 33198 33312
rect 33229 33303 33287 33309
rect 33229 33269 33241 33303
rect 33275 33300 33287 33303
rect 33318 33300 33324 33312
rect 33275 33272 33324 33300
rect 33275 33269 33287 33272
rect 33229 33263 33287 33269
rect 33318 33260 33324 33272
rect 33376 33260 33382 33312
rect 35437 33303 35495 33309
rect 35437 33269 35449 33303
rect 35483 33300 35495 33303
rect 35986 33300 35992 33312
rect 35483 33272 35992 33300
rect 35483 33269 35495 33272
rect 35437 33263 35495 33269
rect 35986 33260 35992 33272
rect 36044 33260 36050 33312
rect 46845 33303 46903 33309
rect 46845 33269 46857 33303
rect 46891 33300 46903 33303
rect 47210 33300 47216 33312
rect 46891 33272 47216 33300
rect 46891 33269 46903 33272
rect 46845 33263 46903 33269
rect 47210 33260 47216 33272
rect 47268 33260 47274 33312
rect 47854 33300 47860 33312
rect 47815 33272 47860 33300
rect 47854 33260 47860 33272
rect 47912 33260 47918 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1670 33056 1676 33108
rect 1728 33096 1734 33108
rect 2777 33099 2835 33105
rect 2777 33096 2789 33099
rect 1728 33068 2789 33096
rect 1728 33056 1734 33068
rect 2777 33065 2789 33068
rect 2823 33065 2835 33099
rect 2777 33059 2835 33065
rect 3694 33056 3700 33108
rect 3752 33096 3758 33108
rect 3789 33099 3847 33105
rect 3789 33096 3801 33099
rect 3752 33068 3801 33096
rect 3752 33056 3758 33068
rect 3789 33065 3801 33068
rect 3835 33065 3847 33099
rect 3789 33059 3847 33065
rect 20990 33056 20996 33108
rect 21048 33096 21054 33108
rect 22649 33099 22707 33105
rect 22649 33096 22661 33099
rect 21048 33068 22661 33096
rect 21048 33056 21054 33068
rect 22649 33065 22661 33068
rect 22695 33065 22707 33099
rect 25038 33096 25044 33108
rect 24999 33068 25044 33096
rect 22649 33059 22707 33065
rect 25038 33056 25044 33068
rect 25096 33056 25102 33108
rect 25869 33099 25927 33105
rect 25869 33065 25881 33099
rect 25915 33096 25927 33099
rect 26234 33096 26240 33108
rect 25915 33068 26240 33096
rect 25915 33065 25927 33068
rect 25869 33059 25927 33065
rect 26234 33056 26240 33068
rect 26292 33056 26298 33108
rect 27706 33056 27712 33108
rect 27764 33096 27770 33108
rect 28353 33099 28411 33105
rect 28353 33096 28365 33099
rect 27764 33068 28365 33096
rect 27764 33056 27770 33068
rect 28353 33065 28365 33068
rect 28399 33065 28411 33099
rect 28810 33096 28816 33108
rect 28771 33068 28816 33096
rect 28353 33059 28411 33065
rect 28810 33056 28816 33068
rect 28868 33056 28874 33108
rect 30650 33096 30656 33108
rect 30300 33068 30656 33096
rect 21453 33031 21511 33037
rect 21453 32997 21465 33031
rect 21499 33028 21511 33031
rect 21499 33000 22232 33028
rect 21499 32997 21511 33000
rect 21453 32991 21511 32997
rect 1394 32960 1400 32972
rect 1355 32932 1400 32960
rect 1394 32920 1400 32932
rect 1452 32920 1458 32972
rect 3145 32963 3203 32969
rect 3145 32929 3157 32963
rect 3191 32960 3203 32963
rect 3191 32932 4016 32960
rect 3191 32929 3203 32932
rect 3145 32923 3203 32929
rect 1673 32895 1731 32901
rect 1673 32861 1685 32895
rect 1719 32892 1731 32895
rect 2685 32895 2743 32901
rect 2685 32892 2697 32895
rect 1719 32864 2697 32892
rect 1719 32861 1731 32864
rect 1673 32855 1731 32861
rect 2685 32861 2697 32864
rect 2731 32892 2743 32895
rect 2774 32892 2780 32904
rect 2731 32864 2780 32892
rect 2731 32861 2743 32864
rect 2685 32855 2743 32861
rect 2774 32852 2780 32864
rect 2832 32852 2838 32904
rect 3988 32901 4016 32932
rect 13262 32920 13268 32972
rect 13320 32960 13326 32972
rect 14093 32963 14151 32969
rect 14093 32960 14105 32963
rect 13320 32932 14105 32960
rect 13320 32920 13326 32932
rect 14093 32929 14105 32932
rect 14139 32929 14151 32963
rect 15930 32960 15936 32972
rect 15891 32932 15936 32960
rect 14093 32923 14151 32929
rect 15930 32920 15936 32932
rect 15988 32920 15994 32972
rect 21177 32963 21235 32969
rect 21177 32929 21189 32963
rect 21223 32960 21235 32963
rect 21542 32960 21548 32972
rect 21223 32932 21548 32960
rect 21223 32929 21235 32932
rect 21177 32923 21235 32929
rect 21542 32920 21548 32932
rect 21600 32960 21606 32972
rect 22002 32960 22008 32972
rect 21600 32932 22008 32960
rect 21600 32920 21606 32932
rect 22002 32920 22008 32932
rect 22060 32920 22066 32972
rect 22204 32969 22232 33000
rect 25958 32988 25964 33040
rect 26016 33028 26022 33040
rect 26145 33031 26203 33037
rect 26145 33028 26157 33031
rect 26016 33000 26157 33028
rect 26016 32988 26022 33000
rect 26145 32997 26157 33000
rect 26191 33028 26203 33031
rect 27249 33031 27307 33037
rect 26191 33000 26832 33028
rect 26191 32997 26203 33000
rect 26145 32991 26203 32997
rect 22189 32963 22247 32969
rect 22189 32929 22201 32963
rect 22235 32929 22247 32963
rect 22189 32923 22247 32929
rect 22281 32963 22339 32969
rect 22281 32929 22293 32963
rect 22327 32960 22339 32963
rect 24578 32960 24584 32972
rect 22327 32932 24584 32960
rect 22327 32929 22339 32932
rect 22281 32923 22339 32929
rect 24578 32920 24584 32932
rect 24636 32920 24642 32972
rect 25590 32920 25596 32972
rect 25648 32960 25654 32972
rect 26804 32969 26832 33000
rect 27249 32997 27261 33031
rect 27295 33028 27307 33031
rect 27982 33028 27988 33040
rect 27295 33000 27988 33028
rect 27295 32997 27307 33000
rect 27249 32991 27307 32997
rect 27982 32988 27988 33000
rect 28040 32988 28046 33040
rect 28258 32988 28264 33040
rect 28316 33028 28322 33040
rect 30300 33028 30328 33068
rect 30650 33056 30656 33068
rect 30708 33056 30714 33108
rect 30742 33056 30748 33108
rect 30800 33096 30806 33108
rect 31021 33099 31079 33105
rect 31021 33096 31033 33099
rect 30800 33068 31033 33096
rect 30800 33056 30806 33068
rect 31021 33065 31033 33068
rect 31067 33065 31079 33099
rect 31021 33059 31079 33065
rect 32306 33056 32312 33108
rect 32364 33096 32370 33108
rect 32490 33096 32496 33108
rect 32364 33068 32496 33096
rect 32364 33056 32370 33068
rect 32490 33056 32496 33068
rect 32548 33056 32554 33108
rect 28316 33000 30328 33028
rect 28316 32988 28322 33000
rect 30374 32988 30380 33040
rect 30432 33028 30438 33040
rect 32858 33028 32864 33040
rect 30432 33000 32864 33028
rect 30432 32988 30438 33000
rect 32858 32988 32864 33000
rect 32916 32988 32922 33040
rect 47026 32988 47032 33040
rect 47084 33028 47090 33040
rect 47084 33000 47440 33028
rect 47084 32988 47090 33000
rect 25777 32963 25835 32969
rect 25777 32960 25789 32963
rect 25648 32932 25789 32960
rect 25648 32920 25654 32932
rect 25777 32929 25789 32932
rect 25823 32929 25835 32963
rect 25777 32923 25835 32929
rect 26789 32963 26847 32969
rect 26789 32929 26801 32963
rect 26835 32929 26847 32963
rect 26789 32923 26847 32929
rect 28000 32932 29132 32960
rect 3973 32895 4031 32901
rect 3973 32861 3985 32895
rect 4019 32861 4031 32895
rect 3973 32855 4031 32861
rect 9582 32852 9588 32904
rect 9640 32892 9646 32904
rect 13357 32895 13415 32901
rect 13357 32892 13369 32895
rect 9640 32864 13369 32892
rect 9640 32852 9646 32864
rect 13357 32861 13369 32864
rect 13403 32892 13415 32895
rect 13998 32892 14004 32904
rect 13403 32864 14004 32892
rect 13403 32861 13415 32864
rect 13357 32855 13415 32861
rect 13998 32852 14004 32864
rect 14056 32852 14062 32904
rect 21082 32892 21088 32904
rect 21043 32864 21088 32892
rect 21082 32852 21088 32864
rect 21140 32852 21146 32904
rect 21266 32852 21272 32904
rect 21324 32892 21330 32904
rect 21913 32895 21971 32901
rect 21913 32892 21925 32895
rect 21324 32864 21925 32892
rect 21324 32852 21330 32864
rect 21913 32861 21925 32864
rect 21959 32861 21971 32895
rect 21913 32855 21971 32861
rect 22097 32895 22155 32901
rect 22097 32861 22109 32895
rect 22143 32892 22155 32895
rect 22370 32892 22376 32904
rect 22143 32864 22376 32892
rect 22143 32861 22155 32864
rect 22097 32855 22155 32861
rect 22370 32852 22376 32864
rect 22428 32852 22434 32904
rect 22465 32895 22523 32901
rect 22465 32861 22477 32895
rect 22511 32892 22523 32895
rect 22554 32892 22560 32904
rect 22511 32864 22560 32892
rect 22511 32861 22523 32864
rect 22465 32855 22523 32861
rect 22554 32852 22560 32864
rect 22612 32852 22618 32904
rect 24762 32852 24768 32904
rect 24820 32892 24826 32904
rect 24857 32895 24915 32901
rect 24857 32892 24869 32895
rect 24820 32864 24869 32892
rect 24820 32852 24826 32864
rect 24857 32861 24869 32864
rect 24903 32861 24915 32895
rect 24857 32855 24915 32861
rect 25133 32895 25191 32901
rect 25133 32861 25145 32895
rect 25179 32861 25191 32895
rect 25133 32855 25191 32861
rect 13449 32827 13507 32833
rect 13449 32793 13461 32827
rect 13495 32824 13507 32827
rect 14277 32827 14335 32833
rect 14277 32824 14289 32827
rect 13495 32796 14289 32824
rect 13495 32793 13507 32796
rect 13449 32787 13507 32793
rect 14277 32793 14289 32796
rect 14323 32793 14335 32827
rect 14277 32787 14335 32793
rect 22738 32716 22744 32768
rect 22796 32756 22802 32768
rect 24673 32759 24731 32765
rect 24673 32756 24685 32759
rect 22796 32728 24685 32756
rect 22796 32716 22802 32728
rect 24673 32725 24685 32728
rect 24719 32725 24731 32759
rect 25148 32756 25176 32855
rect 25222 32852 25228 32904
rect 25280 32892 25286 32904
rect 28000 32901 28028 32932
rect 29104 32904 29132 32932
rect 29546 32920 29552 32972
rect 29604 32960 29610 32972
rect 30561 32963 30619 32969
rect 29604 32932 30512 32960
rect 29604 32920 29610 32932
rect 25961 32895 26019 32901
rect 25961 32892 25973 32895
rect 25280 32864 25973 32892
rect 25280 32852 25286 32864
rect 25961 32861 25973 32864
rect 26007 32861 26019 32895
rect 25961 32855 26019 32861
rect 26881 32895 26939 32901
rect 26881 32861 26893 32895
rect 26927 32861 26939 32895
rect 26881 32855 26939 32861
rect 27985 32895 28043 32901
rect 27985 32861 27997 32895
rect 28031 32861 28043 32895
rect 27985 32855 28043 32861
rect 28169 32895 28227 32901
rect 28169 32861 28181 32895
rect 28215 32892 28227 32895
rect 28534 32892 28540 32904
rect 28215 32864 28540 32892
rect 28215 32861 28227 32864
rect 28169 32855 28227 32861
rect 25682 32824 25688 32836
rect 25643 32796 25688 32824
rect 25682 32784 25688 32796
rect 25740 32784 25746 32836
rect 25774 32784 25780 32836
rect 25832 32824 25838 32836
rect 26896 32824 26924 32855
rect 28184 32824 28212 32855
rect 28534 32852 28540 32864
rect 28592 32852 28598 32904
rect 28718 32852 28724 32904
rect 28776 32892 28782 32904
rect 28813 32895 28871 32901
rect 28813 32892 28825 32895
rect 28776 32864 28825 32892
rect 28776 32852 28782 32864
rect 28813 32861 28825 32864
rect 28859 32861 28871 32895
rect 28813 32855 28871 32861
rect 28997 32895 29055 32901
rect 28997 32861 29009 32895
rect 29043 32861 29055 32895
rect 28997 32855 29055 32861
rect 25832 32796 28212 32824
rect 29012 32824 29040 32855
rect 29086 32852 29092 32904
rect 29144 32892 29150 32904
rect 29144 32864 29189 32892
rect 29144 32852 29150 32864
rect 29914 32852 29920 32904
rect 29972 32892 29978 32904
rect 30484 32901 30512 32932
rect 30561 32929 30573 32963
rect 30607 32960 30619 32963
rect 30926 32960 30932 32972
rect 30607 32932 30932 32960
rect 30607 32929 30619 32932
rect 30561 32923 30619 32929
rect 30926 32920 30932 32932
rect 30984 32920 30990 32972
rect 33134 32960 33140 32972
rect 32508 32932 33140 32960
rect 32508 32904 32536 32932
rect 33134 32920 33140 32932
rect 33192 32920 33198 32972
rect 34974 32960 34980 32972
rect 33428 32932 34980 32960
rect 30285 32895 30343 32901
rect 30285 32892 30297 32895
rect 29972 32864 30297 32892
rect 29972 32852 29978 32864
rect 30285 32861 30297 32864
rect 30331 32861 30343 32895
rect 30285 32855 30343 32861
rect 30469 32895 30527 32901
rect 30469 32861 30481 32895
rect 30515 32861 30527 32895
rect 30469 32855 30527 32861
rect 30650 32852 30656 32904
rect 30708 32892 30714 32904
rect 30708 32864 30753 32892
rect 30708 32852 30714 32864
rect 30834 32852 30840 32904
rect 30892 32892 30898 32904
rect 32490 32892 32496 32904
rect 30892 32864 31754 32892
rect 32451 32864 32496 32892
rect 30892 32852 30898 32864
rect 30009 32827 30067 32833
rect 29012 32796 29684 32824
rect 25832 32784 25838 32796
rect 29012 32756 29040 32796
rect 25148 32728 29040 32756
rect 29273 32759 29331 32765
rect 24673 32719 24731 32725
rect 29273 32725 29285 32759
rect 29319 32756 29331 32759
rect 29546 32756 29552 32768
rect 29319 32728 29552 32756
rect 29319 32725 29331 32728
rect 29273 32719 29331 32725
rect 29546 32716 29552 32728
rect 29604 32716 29610 32768
rect 29656 32756 29684 32796
rect 30009 32793 30021 32827
rect 30055 32824 30067 32827
rect 30668 32824 30696 32852
rect 30055 32796 30696 32824
rect 31726 32824 31754 32864
rect 32490 32852 32496 32864
rect 32548 32852 32554 32904
rect 32677 32895 32735 32901
rect 32677 32861 32689 32895
rect 32723 32892 32735 32895
rect 33042 32892 33048 32904
rect 32723 32864 33048 32892
rect 32723 32861 32735 32864
rect 32677 32855 32735 32861
rect 33042 32852 33048 32864
rect 33100 32852 33106 32904
rect 33428 32824 33456 32932
rect 34974 32920 34980 32932
rect 35032 32920 35038 32972
rect 47118 32960 47124 32972
rect 47079 32932 47124 32960
rect 47118 32920 47124 32932
rect 47176 32920 47182 32972
rect 47412 32969 47440 33000
rect 47397 32963 47455 32969
rect 47397 32929 47409 32963
rect 47443 32929 47455 32963
rect 47397 32923 47455 32929
rect 33502 32852 33508 32904
rect 33560 32892 33566 32904
rect 34701 32895 34759 32901
rect 34701 32892 34713 32895
rect 33560 32864 34713 32892
rect 33560 32852 33566 32864
rect 34701 32861 34713 32864
rect 34747 32861 34759 32895
rect 34701 32855 34759 32861
rect 46290 32852 46296 32904
rect 46348 32892 46354 32904
rect 46569 32895 46627 32901
rect 46569 32892 46581 32895
rect 46348 32864 46581 32892
rect 46348 32852 46354 32864
rect 46569 32861 46581 32864
rect 46615 32861 46627 32895
rect 46569 32855 46627 32861
rect 33778 32824 33784 32836
rect 31726 32796 33456 32824
rect 33739 32796 33784 32824
rect 30055 32793 30067 32796
rect 30009 32787 30067 32793
rect 33778 32784 33784 32796
rect 33836 32784 33842 32836
rect 33965 32827 34023 32833
rect 33965 32793 33977 32827
rect 34011 32824 34023 32827
rect 34977 32827 35035 32833
rect 34011 32796 34560 32824
rect 34011 32793 34023 32796
rect 33965 32787 34023 32793
rect 30558 32756 30564 32768
rect 29656 32728 30564 32756
rect 30558 32716 30564 32728
rect 30616 32716 30622 32768
rect 30742 32716 30748 32768
rect 30800 32756 30806 32768
rect 32950 32756 32956 32768
rect 30800 32728 32956 32756
rect 30800 32716 30806 32728
rect 32950 32716 32956 32728
rect 33008 32716 33014 32768
rect 33042 32716 33048 32768
rect 33100 32756 33106 32768
rect 33980 32756 34008 32787
rect 33100 32728 34008 32756
rect 34149 32759 34207 32765
rect 33100 32716 33106 32728
rect 34149 32725 34161 32759
rect 34195 32756 34207 32759
rect 34422 32756 34428 32768
rect 34195 32728 34428 32756
rect 34195 32725 34207 32728
rect 34149 32719 34207 32725
rect 34422 32716 34428 32728
rect 34480 32716 34486 32768
rect 34532 32756 34560 32796
rect 34977 32793 34989 32827
rect 35023 32824 35035 32827
rect 35066 32824 35072 32836
rect 35023 32796 35072 32824
rect 35023 32793 35035 32796
rect 34977 32787 35035 32793
rect 35066 32784 35072 32796
rect 35124 32784 35130 32836
rect 35986 32784 35992 32836
rect 36044 32784 36050 32836
rect 47210 32784 47216 32836
rect 47268 32824 47274 32836
rect 47268 32796 47313 32824
rect 47268 32784 47274 32796
rect 36449 32759 36507 32765
rect 36449 32756 36461 32759
rect 34532 32728 36461 32756
rect 36449 32725 36461 32728
rect 36495 32725 36507 32759
rect 36449 32719 36507 32725
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 3142 32512 3148 32564
rect 3200 32552 3206 32564
rect 41138 32552 41144 32564
rect 3200 32524 41144 32552
rect 3200 32512 3206 32524
rect 41138 32512 41144 32524
rect 41196 32512 41202 32564
rect 2774 32484 2780 32496
rect 2735 32456 2780 32484
rect 2774 32444 2780 32456
rect 2832 32444 2838 32496
rect 8294 32444 8300 32496
rect 8352 32484 8358 32496
rect 8352 32456 10548 32484
rect 8352 32444 8358 32456
rect 2590 32348 2596 32360
rect 2551 32320 2596 32348
rect 2590 32308 2596 32320
rect 2648 32308 2654 32360
rect 4433 32351 4491 32357
rect 4433 32317 4445 32351
rect 4479 32348 4491 32351
rect 4614 32348 4620 32360
rect 4479 32320 4620 32348
rect 4479 32317 4491 32320
rect 4433 32311 4491 32317
rect 4614 32308 4620 32320
rect 4672 32308 4678 32360
rect 9125 32351 9183 32357
rect 9125 32317 9137 32351
rect 9171 32317 9183 32351
rect 9125 32311 9183 32317
rect 9309 32351 9367 32357
rect 9309 32317 9321 32351
rect 9355 32348 9367 32351
rect 9766 32348 9772 32360
rect 9355 32320 9772 32348
rect 9355 32317 9367 32320
rect 9309 32311 9367 32317
rect 2038 32172 2044 32224
rect 2096 32212 2102 32224
rect 2133 32215 2191 32221
rect 2133 32212 2145 32215
rect 2096 32184 2145 32212
rect 2096 32172 2102 32184
rect 2133 32181 2145 32184
rect 2179 32181 2191 32215
rect 9140 32212 9168 32311
rect 9766 32308 9772 32320
rect 9824 32308 9830 32360
rect 10520 32357 10548 32456
rect 12526 32444 12532 32496
rect 12584 32444 12590 32496
rect 14093 32487 14151 32493
rect 14093 32453 14105 32487
rect 14139 32484 14151 32487
rect 14182 32484 14188 32496
rect 14139 32456 14188 32484
rect 14139 32453 14151 32456
rect 14093 32447 14151 32453
rect 14182 32444 14188 32456
rect 14240 32444 14246 32496
rect 20346 32444 20352 32496
rect 20404 32484 20410 32496
rect 20901 32487 20959 32493
rect 20901 32484 20913 32487
rect 20404 32456 20913 32484
rect 20404 32444 20410 32456
rect 20901 32453 20913 32456
rect 20947 32453 20959 32487
rect 21266 32484 21272 32496
rect 21227 32456 21272 32484
rect 20901 32447 20959 32453
rect 21266 32444 21272 32456
rect 21324 32444 21330 32496
rect 21450 32444 21456 32496
rect 21508 32484 21514 32496
rect 22005 32487 22063 32493
rect 22005 32484 22017 32487
rect 21508 32456 22017 32484
rect 21508 32444 21514 32456
rect 22005 32453 22017 32456
rect 22051 32453 22063 32487
rect 22005 32447 22063 32453
rect 22094 32444 22100 32496
rect 22152 32484 22158 32496
rect 22189 32487 22247 32493
rect 22189 32484 22201 32487
rect 22152 32456 22201 32484
rect 22152 32444 22158 32456
rect 22189 32453 22201 32456
rect 22235 32453 22247 32487
rect 22189 32447 22247 32453
rect 25038 32444 25044 32496
rect 25096 32484 25102 32496
rect 25133 32487 25191 32493
rect 25133 32484 25145 32487
rect 25096 32456 25145 32484
rect 25096 32444 25102 32456
rect 25133 32453 25145 32456
rect 25179 32453 25191 32487
rect 25133 32447 25191 32453
rect 25498 32444 25504 32496
rect 25556 32484 25562 32496
rect 25958 32484 25964 32496
rect 25556 32456 25964 32484
rect 25556 32444 25562 32456
rect 25958 32444 25964 32456
rect 26016 32444 26022 32496
rect 27154 32484 27160 32496
rect 27115 32456 27160 32484
rect 27154 32444 27160 32456
rect 27212 32444 27218 32496
rect 29638 32484 29644 32496
rect 27264 32456 29644 32484
rect 13998 32416 14004 32428
rect 13959 32388 14004 32416
rect 13998 32376 14004 32388
rect 14056 32376 14062 32428
rect 21085 32419 21143 32425
rect 21085 32385 21097 32419
rect 21131 32416 21143 32419
rect 21726 32416 21732 32428
rect 21131 32388 21732 32416
rect 21131 32385 21143 32388
rect 21085 32379 21143 32385
rect 21726 32376 21732 32388
rect 21784 32376 21790 32428
rect 21821 32419 21879 32425
rect 21821 32385 21833 32419
rect 21867 32416 21879 32419
rect 21910 32416 21916 32428
rect 21867 32388 21916 32416
rect 21867 32385 21879 32388
rect 21821 32379 21879 32385
rect 21910 32376 21916 32388
rect 21968 32376 21974 32428
rect 24762 32376 24768 32428
rect 24820 32416 24826 32428
rect 25409 32419 25467 32425
rect 25409 32416 25421 32419
rect 24820 32388 25421 32416
rect 24820 32376 24826 32388
rect 25409 32385 25421 32388
rect 25455 32385 25467 32419
rect 25409 32379 25467 32385
rect 25590 32376 25596 32428
rect 25648 32376 25654 32428
rect 26973 32419 27031 32425
rect 26973 32385 26985 32419
rect 27019 32416 27031 32419
rect 27264 32416 27292 32456
rect 29638 32444 29644 32456
rect 29696 32444 29702 32496
rect 29914 32484 29920 32496
rect 29875 32456 29920 32484
rect 29914 32444 29920 32456
rect 29972 32444 29978 32496
rect 30926 32484 30932 32496
rect 30208 32456 30932 32484
rect 27019 32388 27292 32416
rect 27019 32385 27031 32388
rect 26973 32379 27031 32385
rect 10505 32351 10563 32357
rect 10505 32317 10517 32351
rect 10551 32317 10563 32351
rect 10505 32311 10563 32317
rect 10778 32308 10784 32360
rect 10836 32348 10842 32360
rect 11517 32351 11575 32357
rect 11517 32348 11529 32351
rect 10836 32320 11529 32348
rect 10836 32308 10842 32320
rect 11517 32317 11529 32320
rect 11563 32317 11575 32351
rect 11790 32348 11796 32360
rect 11751 32320 11796 32348
rect 11517 32311 11575 32317
rect 11790 32308 11796 32320
rect 11848 32308 11854 32360
rect 13262 32348 13268 32360
rect 13223 32320 13268 32348
rect 13262 32308 13268 32320
rect 13320 32348 13326 32360
rect 13538 32348 13544 32360
rect 13320 32320 13544 32348
rect 13320 32308 13326 32320
rect 13538 32308 13544 32320
rect 13596 32308 13602 32360
rect 25317 32351 25375 32357
rect 25317 32317 25329 32351
rect 25363 32348 25375 32351
rect 25608 32348 25636 32376
rect 26988 32348 27016 32379
rect 27982 32376 27988 32428
rect 28040 32416 28046 32428
rect 28353 32419 28411 32425
rect 28353 32416 28365 32419
rect 28040 32388 28365 32416
rect 28040 32376 28046 32388
rect 28353 32385 28365 32388
rect 28399 32416 28411 32419
rect 28626 32416 28632 32428
rect 28399 32388 28632 32416
rect 28399 32385 28411 32388
rect 28353 32379 28411 32385
rect 28626 32376 28632 32388
rect 28684 32376 28690 32428
rect 28997 32419 29055 32425
rect 28997 32385 29009 32419
rect 29043 32416 29055 32419
rect 29086 32416 29092 32428
rect 29043 32388 29092 32416
rect 29043 32385 29055 32388
rect 28997 32379 29055 32385
rect 29086 32376 29092 32388
rect 29144 32376 29150 32428
rect 30098 32416 30104 32428
rect 30059 32388 30104 32416
rect 30098 32376 30104 32388
rect 30156 32376 30162 32428
rect 30208 32425 30236 32456
rect 30926 32444 30932 32456
rect 30984 32444 30990 32496
rect 32858 32444 32864 32496
rect 32916 32484 32922 32496
rect 32916 32456 33548 32484
rect 32916 32444 32922 32456
rect 30193 32419 30251 32425
rect 30193 32385 30205 32419
rect 30239 32385 30251 32419
rect 30193 32379 30251 32385
rect 30377 32419 30435 32425
rect 30377 32385 30389 32419
rect 30423 32385 30435 32419
rect 30377 32379 30435 32385
rect 25363 32320 27016 32348
rect 25363 32317 25375 32320
rect 25317 32311 25375 32317
rect 27890 32308 27896 32360
rect 27948 32348 27954 32360
rect 28074 32348 28080 32360
rect 27948 32320 28080 32348
rect 27948 32308 27954 32320
rect 28074 32308 28080 32320
rect 28132 32348 28138 32360
rect 28537 32351 28595 32357
rect 28537 32348 28549 32351
rect 28132 32320 28549 32348
rect 28132 32308 28138 32320
rect 28537 32317 28549 32320
rect 28583 32317 28595 32351
rect 28537 32311 28595 32317
rect 28810 32308 28816 32360
rect 28868 32348 28874 32360
rect 30392 32348 30420 32379
rect 30466 32376 30472 32428
rect 30524 32416 30530 32428
rect 31021 32419 31079 32425
rect 31021 32416 31033 32419
rect 30524 32388 31033 32416
rect 30524 32376 30530 32388
rect 31021 32385 31033 32388
rect 31067 32385 31079 32419
rect 32306 32416 32312 32428
rect 32267 32388 32312 32416
rect 31021 32379 31079 32385
rect 32306 32376 32312 32388
rect 32364 32376 32370 32428
rect 33318 32416 33324 32428
rect 33279 32388 33324 32416
rect 33318 32376 33324 32388
rect 33376 32376 33382 32428
rect 33520 32425 33548 32456
rect 35066 32444 35072 32496
rect 35124 32484 35130 32496
rect 35161 32487 35219 32493
rect 35161 32484 35173 32487
rect 35124 32456 35173 32484
rect 35124 32444 35130 32456
rect 35161 32453 35173 32456
rect 35207 32453 35219 32487
rect 35161 32447 35219 32453
rect 33505 32419 33563 32425
rect 33505 32385 33517 32419
rect 33551 32385 33563 32419
rect 34422 32416 34428 32428
rect 34383 32388 34428 32416
rect 33505 32379 33563 32385
rect 34422 32376 34428 32388
rect 34480 32376 34486 32428
rect 34514 32376 34520 32428
rect 34572 32416 34578 32428
rect 34609 32419 34667 32425
rect 34609 32416 34621 32419
rect 34572 32388 34621 32416
rect 34572 32376 34578 32388
rect 34609 32385 34621 32388
rect 34655 32385 34667 32419
rect 34974 32416 34980 32428
rect 34935 32388 34980 32416
rect 34609 32379 34667 32385
rect 34974 32376 34980 32388
rect 35032 32416 35038 32428
rect 35434 32416 35440 32428
rect 35032 32388 35440 32416
rect 35032 32376 35038 32388
rect 35434 32376 35440 32388
rect 35492 32376 35498 32428
rect 46477 32419 46535 32425
rect 46477 32416 46489 32419
rect 35866 32388 46489 32416
rect 28868 32320 30420 32348
rect 28868 32308 28874 32320
rect 30558 32308 30564 32360
rect 30616 32348 30622 32360
rect 32217 32351 32275 32357
rect 32217 32348 32229 32351
rect 30616 32320 32229 32348
rect 30616 32308 30622 32320
rect 32217 32317 32229 32320
rect 32263 32348 32275 32351
rect 32490 32348 32496 32360
rect 32263 32320 32496 32348
rect 32263 32317 32275 32320
rect 32217 32311 32275 32317
rect 32490 32308 32496 32320
rect 32548 32308 32554 32360
rect 33413 32351 33471 32357
rect 33413 32317 33425 32351
rect 33459 32348 33471 32351
rect 34701 32351 34759 32357
rect 34701 32348 34713 32351
rect 33459 32320 34713 32348
rect 33459 32317 33471 32320
rect 33413 32311 33471 32317
rect 34701 32317 34713 32320
rect 34747 32317 34759 32351
rect 34701 32311 34759 32317
rect 34793 32351 34851 32357
rect 34793 32317 34805 32351
rect 34839 32348 34851 32351
rect 35866 32348 35894 32388
rect 46477 32385 46489 32388
rect 46523 32385 46535 32419
rect 46477 32379 46535 32385
rect 47486 32376 47492 32428
rect 47544 32416 47550 32428
rect 47581 32419 47639 32425
rect 47581 32416 47593 32419
rect 47544 32388 47593 32416
rect 47544 32376 47550 32388
rect 47581 32385 47593 32388
rect 47627 32385 47639 32419
rect 47581 32379 47639 32385
rect 46198 32348 46204 32360
rect 34839 32320 35894 32348
rect 46159 32320 46204 32348
rect 34839 32317 34851 32320
rect 34793 32311 34851 32317
rect 46198 32308 46204 32320
rect 46256 32308 46262 32360
rect 22278 32240 22284 32292
rect 22336 32280 22342 32292
rect 25593 32283 25651 32289
rect 25593 32280 25605 32283
rect 22336 32252 25605 32280
rect 22336 32240 22342 32252
rect 25593 32249 25605 32252
rect 25639 32249 25651 32283
rect 25593 32243 25651 32249
rect 25958 32240 25964 32292
rect 26016 32280 26022 32292
rect 27341 32283 27399 32289
rect 26016 32252 27016 32280
rect 26016 32240 26022 32252
rect 12986 32212 12992 32224
rect 9140 32184 12992 32212
rect 2133 32175 2191 32181
rect 12986 32172 12992 32184
rect 13044 32212 13050 32224
rect 14550 32212 14556 32224
rect 13044 32184 14556 32212
rect 13044 32172 13050 32184
rect 14550 32172 14556 32184
rect 14608 32172 14614 32224
rect 22554 32172 22560 32224
rect 22612 32212 22618 32224
rect 23382 32212 23388 32224
rect 22612 32184 23388 32212
rect 22612 32172 22618 32184
rect 23382 32172 23388 32184
rect 23440 32172 23446 32224
rect 25409 32215 25467 32221
rect 25409 32181 25421 32215
rect 25455 32212 25467 32215
rect 26786 32212 26792 32224
rect 25455 32184 26792 32212
rect 25455 32181 25467 32184
rect 25409 32175 25467 32181
rect 26786 32172 26792 32184
rect 26844 32172 26850 32224
rect 26988 32212 27016 32252
rect 27341 32249 27353 32283
rect 27387 32280 27399 32283
rect 30576 32280 30604 32308
rect 34514 32280 34520 32292
rect 27387 32252 30604 32280
rect 31220 32252 34520 32280
rect 27387 32249 27399 32252
rect 27341 32243 27399 32249
rect 31220 32224 31248 32252
rect 34514 32240 34520 32252
rect 34572 32240 34578 32292
rect 29181 32215 29239 32221
rect 29181 32212 29193 32215
rect 26988 32184 29193 32212
rect 29181 32181 29193 32184
rect 29227 32212 29239 32215
rect 30742 32212 30748 32224
rect 29227 32184 30748 32212
rect 29227 32181 29239 32184
rect 29181 32175 29239 32181
rect 30742 32172 30748 32184
rect 30800 32172 30806 32224
rect 31202 32212 31208 32224
rect 31163 32184 31208 32212
rect 31202 32172 31208 32184
rect 31260 32172 31266 32224
rect 31294 32172 31300 32224
rect 31352 32212 31358 32224
rect 32677 32215 32735 32221
rect 32677 32212 32689 32215
rect 31352 32184 32689 32212
rect 31352 32172 31358 32184
rect 32677 32181 32689 32184
rect 32723 32181 32735 32215
rect 32677 32175 32735 32181
rect 46474 32172 46480 32224
rect 46532 32212 46538 32224
rect 47673 32215 47731 32221
rect 47673 32212 47685 32215
rect 46532 32184 47685 32212
rect 46532 32172 46538 32184
rect 47673 32181 47685 32184
rect 47719 32181 47731 32215
rect 47673 32175 47731 32181
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1397 32011 1455 32017
rect 1397 31977 1409 32011
rect 1443 32008 1455 32011
rect 1670 32008 1676 32020
rect 1443 31980 1676 32008
rect 1443 31977 1455 31980
rect 1397 31971 1455 31977
rect 1670 31968 1676 31980
rect 1728 31968 1734 32020
rect 9766 32008 9772 32020
rect 9727 31980 9772 32008
rect 9766 31968 9772 31980
rect 9824 31968 9830 32020
rect 10778 32008 10784 32020
rect 10739 31980 10784 32008
rect 10778 31968 10784 31980
rect 10836 31968 10842 32020
rect 11790 32008 11796 32020
rect 11751 31980 11796 32008
rect 11790 31968 11796 31980
rect 11848 31968 11854 32020
rect 12526 31968 12532 32020
rect 12584 32008 12590 32020
rect 12621 32011 12679 32017
rect 12621 32008 12633 32011
rect 12584 31980 12633 32008
rect 12584 31968 12590 31980
rect 12621 31977 12633 31980
rect 12667 31977 12679 32011
rect 15102 32008 15108 32020
rect 15063 31980 15108 32008
rect 12621 31971 12679 31977
rect 15102 31968 15108 31980
rect 15160 31968 15166 32020
rect 21082 31968 21088 32020
rect 21140 32008 21146 32020
rect 21453 32011 21511 32017
rect 21453 32008 21465 32011
rect 21140 31980 21465 32008
rect 21140 31968 21146 31980
rect 21453 31977 21465 31980
rect 21499 32008 21511 32011
rect 22554 32008 22560 32020
rect 21499 31980 22560 32008
rect 21499 31977 21511 31980
rect 21453 31971 21511 31977
rect 22554 31968 22560 31980
rect 22612 31968 22618 32020
rect 22738 32008 22744 32020
rect 22699 31980 22744 32008
rect 22738 31968 22744 31980
rect 22796 31968 22802 32020
rect 22922 32008 22928 32020
rect 22883 31980 22928 32008
rect 22922 31968 22928 31980
rect 22980 31968 22986 32020
rect 24578 31968 24584 32020
rect 24636 32008 24642 32020
rect 25958 32008 25964 32020
rect 24636 31980 25964 32008
rect 24636 31968 24642 31980
rect 25958 31968 25964 31980
rect 26016 31968 26022 32020
rect 26142 31968 26148 32020
rect 26200 32008 26206 32020
rect 26881 32011 26939 32017
rect 26881 32008 26893 32011
rect 26200 31980 26893 32008
rect 26200 31968 26206 31980
rect 26881 31977 26893 31980
rect 26927 32008 26939 32011
rect 27154 32008 27160 32020
rect 26927 31980 27160 32008
rect 26927 31977 26939 31980
rect 26881 31971 26939 31977
rect 27154 31968 27160 31980
rect 27212 31968 27218 32020
rect 27617 32011 27675 32017
rect 27617 31977 27629 32011
rect 27663 32008 27675 32011
rect 28258 32008 28264 32020
rect 27663 31980 28264 32008
rect 27663 31977 27675 31980
rect 27617 31971 27675 31977
rect 28258 31968 28264 31980
rect 28316 31968 28322 32020
rect 28537 32011 28595 32017
rect 28537 31977 28549 32011
rect 28583 32008 28595 32011
rect 29086 32008 29092 32020
rect 28583 31980 29092 32008
rect 28583 31977 28595 31980
rect 28537 31971 28595 31977
rect 29086 31968 29092 31980
rect 29144 31968 29150 32020
rect 31570 32008 31576 32020
rect 29196 31980 31576 32008
rect 11698 31900 11704 31952
rect 11756 31940 11762 31952
rect 11756 31912 22876 31940
rect 11756 31900 11762 31912
rect 11609 31875 11667 31881
rect 11609 31841 11621 31875
rect 11655 31872 11667 31875
rect 13265 31875 13323 31881
rect 13265 31872 13277 31875
rect 11655 31844 13277 31872
rect 11655 31841 11667 31844
rect 11609 31835 11667 31841
rect 13265 31841 13277 31844
rect 13311 31841 13323 31875
rect 14550 31872 14556 31884
rect 14511 31844 14556 31872
rect 13265 31835 13323 31841
rect 14550 31832 14556 31844
rect 14608 31832 14614 31884
rect 20806 31872 20812 31884
rect 19996 31844 20812 31872
rect 1578 31804 1584 31816
rect 1539 31776 1584 31804
rect 1578 31764 1584 31776
rect 1636 31764 1642 31816
rect 2869 31807 2927 31813
rect 2869 31773 2881 31807
rect 2915 31804 2927 31807
rect 3142 31804 3148 31816
rect 2915 31776 3148 31804
rect 2915 31773 2927 31776
rect 2869 31767 2927 31773
rect 3142 31764 3148 31776
rect 3200 31764 3206 31816
rect 9582 31764 9588 31816
rect 9640 31804 9646 31816
rect 9677 31807 9735 31813
rect 9677 31804 9689 31807
rect 9640 31776 9689 31804
rect 9640 31764 9646 31776
rect 9677 31773 9689 31776
rect 9723 31773 9735 31807
rect 10686 31804 10692 31816
rect 10647 31776 10692 31804
rect 9677 31767 9735 31773
rect 10686 31764 10692 31776
rect 10744 31764 10750 31816
rect 11517 31807 11575 31813
rect 11517 31773 11529 31807
rect 11563 31804 11575 31807
rect 12434 31804 12440 31816
rect 11563 31776 12440 31804
rect 11563 31773 11575 31776
rect 11517 31767 11575 31773
rect 12434 31764 12440 31776
rect 12492 31764 12498 31816
rect 12529 31807 12587 31813
rect 12529 31773 12541 31807
rect 12575 31804 12587 31807
rect 13170 31804 13176 31816
rect 12575 31776 12609 31804
rect 13131 31776 13176 31804
rect 12575 31773 12587 31776
rect 12529 31767 12587 31773
rect 12250 31696 12256 31748
rect 12308 31736 12314 31748
rect 12544 31736 12572 31767
rect 13170 31764 13176 31776
rect 13228 31764 13234 31816
rect 13354 31804 13360 31816
rect 13315 31776 13360 31804
rect 13354 31764 13360 31776
rect 13412 31764 13418 31816
rect 14274 31804 14280 31816
rect 14235 31776 14280 31804
rect 14274 31764 14280 31776
rect 14332 31764 14338 31816
rect 14458 31804 14464 31816
rect 14419 31776 14464 31804
rect 14458 31764 14464 31776
rect 14516 31764 14522 31816
rect 19996 31813 20024 31844
rect 20806 31832 20812 31844
rect 20864 31832 20870 31884
rect 21450 31872 21456 31884
rect 21284 31844 21456 31872
rect 15013 31807 15071 31813
rect 15013 31773 15025 31807
rect 15059 31804 15071 31807
rect 19981 31807 20039 31813
rect 15059 31776 15093 31804
rect 15059 31773 15071 31776
rect 15013 31767 15071 31773
rect 19981 31773 19993 31807
rect 20027 31773 20039 31807
rect 19981 31767 20039 31773
rect 20073 31807 20131 31813
rect 20073 31773 20085 31807
rect 20119 31804 20131 31807
rect 20162 31804 20168 31816
rect 20119 31776 20168 31804
rect 20119 31773 20131 31776
rect 20073 31767 20131 31773
rect 15028 31736 15056 31767
rect 20162 31764 20168 31776
rect 20220 31764 20226 31816
rect 21284 31813 21312 31844
rect 21450 31832 21456 31844
rect 21508 31832 21514 31884
rect 22094 31832 22100 31884
rect 22152 31872 22158 31884
rect 22554 31872 22560 31884
rect 22152 31844 22560 31872
rect 22152 31832 22158 31844
rect 21269 31807 21327 31813
rect 21269 31773 21281 31807
rect 21315 31773 21327 31807
rect 21269 31767 21327 31773
rect 21358 31764 21364 31816
rect 21416 31804 21422 31816
rect 22388 31813 22416 31844
rect 22554 31832 22560 31844
rect 22612 31832 22618 31884
rect 22848 31872 22876 31912
rect 25038 31900 25044 31952
rect 25096 31940 25102 31952
rect 25866 31940 25872 31952
rect 25096 31912 25872 31940
rect 25096 31900 25102 31912
rect 25866 31900 25872 31912
rect 25924 31940 25930 31952
rect 29196 31940 29224 31980
rect 31570 31968 31576 31980
rect 31628 31968 31634 32020
rect 25924 31912 29224 31940
rect 25924 31900 25930 31912
rect 29270 31900 29276 31952
rect 29328 31940 29334 31952
rect 31202 31940 31208 31952
rect 29328 31912 31208 31940
rect 29328 31900 29334 31912
rect 31202 31900 31208 31912
rect 31260 31900 31266 31952
rect 31294 31900 31300 31952
rect 31352 31900 31358 31952
rect 31849 31943 31907 31949
rect 31849 31909 31861 31943
rect 31895 31940 31907 31943
rect 32674 31940 32680 31952
rect 31895 31912 32680 31940
rect 31895 31909 31907 31912
rect 31849 31903 31907 31909
rect 32674 31900 32680 31912
rect 32732 31900 32738 31952
rect 32769 31943 32827 31949
rect 32769 31909 32781 31943
rect 32815 31940 32827 31943
rect 33226 31940 33232 31952
rect 32815 31912 33232 31940
rect 32815 31909 32827 31912
rect 32769 31903 32827 31909
rect 33226 31900 33232 31912
rect 33284 31900 33290 31952
rect 22848 31844 24624 31872
rect 22373 31807 22431 31813
rect 21416 31776 21461 31804
rect 21416 31764 21422 31776
rect 22373 31773 22385 31807
rect 22419 31804 22431 31807
rect 22738 31804 22744 31816
rect 22419 31776 22453 31804
rect 22699 31776 22744 31804
rect 22419 31773 22431 31776
rect 22373 31767 22431 31773
rect 22738 31764 22744 31776
rect 22796 31764 22802 31816
rect 16850 31736 16856 31748
rect 12308 31708 16856 31736
rect 12308 31696 12314 31708
rect 16850 31696 16856 31708
rect 16908 31696 16914 31748
rect 24596 31736 24624 31844
rect 24688 31844 26280 31872
rect 24688 31813 24716 31844
rect 24673 31807 24731 31813
rect 24673 31773 24685 31807
rect 24719 31773 24731 31807
rect 24949 31807 25007 31813
rect 24949 31804 24961 31807
rect 24673 31767 24731 31773
rect 24780 31776 24961 31804
rect 24780 31736 24808 31776
rect 24949 31773 24961 31776
rect 24995 31773 25007 31807
rect 24949 31767 25007 31773
rect 25038 31764 25044 31816
rect 25096 31764 25102 31816
rect 25406 31764 25412 31816
rect 25464 31804 25470 31816
rect 25682 31804 25688 31816
rect 25464 31776 25544 31804
rect 25643 31776 25688 31804
rect 25464 31764 25470 31776
rect 24596 31708 24808 31736
rect 24857 31739 24915 31745
rect 24857 31705 24869 31739
rect 24903 31736 24915 31739
rect 25056 31736 25084 31764
rect 24903 31708 25084 31736
rect 25516 31736 25544 31776
rect 25682 31764 25688 31776
rect 25740 31764 25746 31816
rect 25774 31764 25780 31816
rect 25832 31804 25838 31816
rect 26050 31804 26056 31816
rect 25832 31776 26056 31804
rect 25832 31764 25838 31776
rect 26050 31764 26056 31776
rect 26108 31764 26114 31816
rect 25869 31739 25927 31745
rect 25869 31736 25881 31739
rect 25516 31708 25881 31736
rect 24903 31705 24915 31708
rect 24857 31699 24915 31705
rect 25869 31705 25881 31708
rect 25915 31705 25927 31739
rect 25869 31699 25927 31705
rect 25961 31739 26019 31745
rect 25961 31705 25973 31739
rect 26007 31705 26019 31739
rect 25961 31699 26019 31705
rect 2958 31668 2964 31680
rect 2919 31640 2964 31668
rect 2958 31628 2964 31640
rect 3016 31628 3022 31680
rect 12434 31628 12440 31680
rect 12492 31668 12498 31680
rect 13538 31668 13544 31680
rect 12492 31640 13544 31668
rect 12492 31628 12498 31640
rect 13538 31628 13544 31640
rect 13596 31628 13602 31680
rect 14090 31668 14096 31680
rect 14051 31640 14096 31668
rect 14090 31628 14096 31640
rect 14148 31628 14154 31680
rect 21634 31668 21640 31680
rect 21595 31640 21640 31668
rect 21634 31628 21640 31640
rect 21692 31628 21698 31680
rect 24486 31668 24492 31680
rect 24447 31640 24492 31668
rect 24486 31628 24492 31640
rect 24544 31628 24550 31680
rect 25976 31668 26004 31699
rect 26050 31668 26056 31680
rect 25976 31640 26056 31668
rect 26050 31628 26056 31640
rect 26108 31628 26114 31680
rect 26252 31677 26280 31844
rect 27890 31832 27896 31884
rect 27948 31872 27954 31884
rect 28258 31872 28264 31884
rect 27948 31844 28264 31872
rect 27948 31832 27954 31844
rect 28258 31832 28264 31844
rect 28316 31832 28322 31884
rect 28442 31832 28448 31884
rect 28500 31872 28506 31884
rect 30466 31872 30472 31884
rect 28500 31844 30472 31872
rect 28500 31832 28506 31844
rect 30466 31832 30472 31844
rect 30524 31872 30530 31884
rect 30524 31844 31156 31872
rect 30524 31832 30530 31844
rect 26786 31804 26792 31816
rect 26747 31776 26792 31804
rect 26786 31764 26792 31776
rect 26844 31764 26850 31816
rect 27798 31764 27804 31816
rect 27856 31804 27862 31816
rect 28721 31807 28779 31813
rect 28721 31804 28733 31807
rect 27856 31776 28733 31804
rect 27856 31764 27862 31776
rect 28721 31773 28733 31776
rect 28767 31804 28779 31807
rect 28767 31776 30052 31804
rect 28767 31773 28779 31776
rect 28721 31767 28779 31773
rect 27522 31736 27528 31748
rect 27483 31708 27528 31736
rect 27522 31696 27528 31708
rect 27580 31696 27586 31748
rect 26237 31671 26295 31677
rect 26237 31637 26249 31671
rect 26283 31637 26295 31671
rect 30024 31668 30052 31776
rect 31128 31736 31156 31844
rect 31312 31813 31340 31900
rect 31389 31875 31447 31881
rect 31389 31841 31401 31875
rect 31435 31872 31447 31875
rect 35342 31872 35348 31884
rect 31435 31844 32168 31872
rect 31435 31841 31447 31844
rect 31389 31835 31447 31841
rect 31297 31807 31355 31813
rect 31297 31773 31309 31807
rect 31343 31773 31355 31807
rect 31481 31807 31539 31813
rect 31481 31804 31493 31807
rect 31297 31767 31355 31773
rect 31404 31776 31493 31804
rect 31404 31736 31432 31776
rect 31481 31773 31493 31776
rect 31527 31773 31539 31807
rect 31481 31767 31539 31773
rect 31570 31764 31576 31816
rect 31628 31804 31634 31816
rect 32140 31813 32168 31844
rect 34716 31844 35348 31872
rect 32306 31813 32312 31816
rect 32125 31807 32183 31813
rect 31628 31776 32076 31804
rect 31628 31764 31634 31776
rect 31128 31708 31432 31736
rect 32048 31736 32076 31776
rect 32125 31773 32137 31807
rect 32171 31773 32183 31807
rect 32125 31767 32183 31773
rect 32273 31807 32312 31813
rect 32273 31773 32285 31807
rect 32273 31767 32312 31773
rect 32306 31764 32312 31767
rect 32364 31764 32370 31816
rect 32401 31807 32459 31813
rect 32401 31773 32413 31807
rect 32447 31773 32459 31807
rect 32401 31767 32459 31773
rect 32416 31736 32444 31767
rect 32490 31764 32496 31816
rect 32548 31804 32554 31816
rect 32674 31813 32680 31816
rect 32631 31807 32680 31813
rect 32548 31776 32593 31804
rect 32548 31764 32554 31776
rect 32631 31773 32643 31807
rect 32677 31773 32680 31807
rect 32631 31767 32680 31773
rect 32674 31764 32680 31767
rect 32732 31764 32738 31816
rect 34716 31813 34744 31844
rect 35342 31832 35348 31844
rect 35400 31832 35406 31884
rect 46290 31872 46296 31884
rect 46251 31844 46296 31872
rect 46290 31832 46296 31844
rect 46348 31832 46354 31884
rect 46474 31872 46480 31884
rect 46435 31844 46480 31872
rect 46474 31832 46480 31844
rect 46532 31832 46538 31884
rect 48130 31872 48136 31884
rect 48091 31844 48136 31872
rect 48130 31832 48136 31844
rect 48188 31832 48194 31884
rect 34701 31807 34759 31813
rect 34701 31773 34713 31807
rect 34747 31773 34759 31807
rect 34701 31767 34759 31773
rect 34790 31764 34796 31816
rect 34848 31804 34854 31816
rect 34848 31776 34893 31804
rect 34848 31764 34854 31776
rect 32048 31708 32444 31736
rect 33778 31668 33784 31680
rect 30024 31640 33784 31668
rect 26237 31631 26295 31637
rect 33778 31628 33784 31640
rect 33836 31628 33842 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 14642 31424 14648 31476
rect 14700 31464 14706 31476
rect 15473 31467 15531 31473
rect 15473 31464 15485 31467
rect 14700 31436 15485 31464
rect 14700 31424 14706 31436
rect 15473 31433 15485 31436
rect 15519 31433 15531 31467
rect 15473 31427 15531 31433
rect 20625 31467 20683 31473
rect 20625 31433 20637 31467
rect 20671 31464 20683 31467
rect 20898 31464 20904 31476
rect 20671 31436 20904 31464
rect 20671 31433 20683 31436
rect 20625 31427 20683 31433
rect 20898 31424 20904 31436
rect 20956 31464 20962 31476
rect 21450 31464 21456 31476
rect 20956 31436 21456 31464
rect 20956 31424 20962 31436
rect 21450 31424 21456 31436
rect 21508 31424 21514 31476
rect 21726 31424 21732 31476
rect 21784 31464 21790 31476
rect 23569 31467 23627 31473
rect 23569 31464 23581 31467
rect 21784 31436 23581 31464
rect 21784 31424 21790 31436
rect 23569 31433 23581 31436
rect 23615 31464 23627 31467
rect 27154 31464 27160 31476
rect 23615 31436 27160 31464
rect 23615 31433 23627 31436
rect 23569 31427 23627 31433
rect 27154 31424 27160 31436
rect 27212 31464 27218 31476
rect 27522 31464 27528 31476
rect 27212 31436 27528 31464
rect 27212 31424 27218 31436
rect 27522 31424 27528 31436
rect 27580 31424 27586 31476
rect 31202 31424 31208 31476
rect 31260 31464 31266 31476
rect 31570 31464 31576 31476
rect 31260 31436 31576 31464
rect 31260 31424 31266 31436
rect 31570 31424 31576 31436
rect 31628 31424 31634 31476
rect 32306 31424 32312 31476
rect 32364 31464 32370 31476
rect 34701 31467 34759 31473
rect 34701 31464 34713 31467
rect 32364 31436 34713 31464
rect 32364 31424 32370 31436
rect 34701 31433 34713 31436
rect 34747 31433 34759 31467
rect 34701 31427 34759 31433
rect 2225 31399 2283 31405
rect 2225 31365 2237 31399
rect 2271 31396 2283 31399
rect 2958 31396 2964 31408
rect 2271 31368 2964 31396
rect 2271 31365 2283 31368
rect 2225 31359 2283 31365
rect 2958 31356 2964 31368
rect 3016 31356 3022 31408
rect 14001 31399 14059 31405
rect 14001 31365 14013 31399
rect 14047 31396 14059 31399
rect 14090 31396 14096 31408
rect 14047 31368 14096 31396
rect 14047 31365 14059 31368
rect 14001 31359 14059 31365
rect 14090 31356 14096 31368
rect 14148 31356 14154 31408
rect 20162 31356 20168 31408
rect 20220 31356 20226 31408
rect 23474 31356 23480 31408
rect 23532 31396 23538 31408
rect 24670 31396 24676 31408
rect 23532 31368 24676 31396
rect 23532 31356 23538 31368
rect 2038 31328 2044 31340
rect 1999 31300 2044 31328
rect 2038 31288 2044 31300
rect 2096 31288 2102 31340
rect 10686 31288 10692 31340
rect 10744 31328 10750 31340
rect 10870 31328 10876 31340
rect 10744 31300 10876 31328
rect 10744 31288 10750 31300
rect 10870 31288 10876 31300
rect 10928 31288 10934 31340
rect 12250 31328 12256 31340
rect 12211 31300 12256 31328
rect 12250 31288 12256 31300
rect 12308 31288 12314 31340
rect 15102 31288 15108 31340
rect 15160 31288 15166 31340
rect 15286 31288 15292 31340
rect 15344 31328 15350 31340
rect 15933 31331 15991 31337
rect 15933 31328 15945 31331
rect 15344 31300 15945 31328
rect 15344 31288 15350 31300
rect 15933 31297 15945 31300
rect 15979 31297 15991 31331
rect 15933 31291 15991 31297
rect 16669 31331 16727 31337
rect 16669 31297 16681 31331
rect 16715 31328 16727 31331
rect 16850 31328 16856 31340
rect 16715 31300 16856 31328
rect 16715 31297 16727 31300
rect 16669 31291 16727 31297
rect 16850 31288 16856 31300
rect 16908 31288 16914 31340
rect 20806 31288 20812 31340
rect 20864 31328 20870 31340
rect 21085 31331 21143 31337
rect 21085 31328 21097 31331
rect 20864 31300 21097 31328
rect 20864 31288 20870 31300
rect 21085 31297 21097 31300
rect 21131 31297 21143 31331
rect 21085 31291 21143 31297
rect 21266 31288 21272 31340
rect 21324 31328 21330 31340
rect 21913 31331 21971 31337
rect 21913 31328 21925 31331
rect 21324 31300 21925 31328
rect 21324 31288 21330 31300
rect 21913 31297 21925 31300
rect 21959 31328 21971 31331
rect 22278 31328 22284 31340
rect 21959 31300 22284 31328
rect 21959 31297 21971 31300
rect 21913 31291 21971 31297
rect 22278 31288 22284 31300
rect 22336 31288 22342 31340
rect 22922 31288 22928 31340
rect 22980 31328 22986 31340
rect 24136 31337 24164 31368
rect 24670 31356 24676 31368
rect 24728 31356 24734 31408
rect 33502 31396 33508 31408
rect 32968 31368 33508 31396
rect 23385 31331 23443 31337
rect 23385 31328 23397 31331
rect 22980 31300 23397 31328
rect 22980 31288 22986 31300
rect 23385 31297 23397 31300
rect 23431 31297 23443 31331
rect 23385 31291 23443 31297
rect 23661 31331 23719 31337
rect 23661 31297 23673 31331
rect 23707 31297 23719 31331
rect 23661 31291 23719 31297
rect 24121 31331 24179 31337
rect 24121 31297 24133 31331
rect 24167 31297 24179 31331
rect 26326 31328 26332 31340
rect 25530 31300 26332 31328
rect 24121 31291 24179 31297
rect 2774 31220 2780 31272
rect 2832 31260 2838 31272
rect 13725 31263 13783 31269
rect 2832 31232 2877 31260
rect 2832 31220 2838 31232
rect 13725 31229 13737 31263
rect 13771 31260 13783 31263
rect 16025 31263 16083 31269
rect 16025 31260 16037 31263
rect 13771 31232 16037 31260
rect 13771 31229 13783 31232
rect 13725 31223 13783 31229
rect 16025 31229 16037 31232
rect 16071 31229 16083 31263
rect 18874 31260 18880 31272
rect 18835 31232 18880 31260
rect 16025 31223 16083 31229
rect 18874 31220 18880 31232
rect 18932 31220 18938 31272
rect 19153 31263 19211 31269
rect 19153 31229 19165 31263
rect 19199 31260 19211 31263
rect 20622 31260 20628 31272
rect 19199 31232 20628 31260
rect 19199 31229 19211 31232
rect 19153 31223 19211 31229
rect 20622 31220 20628 31232
rect 20680 31220 20686 31272
rect 22189 31263 22247 31269
rect 22189 31229 22201 31263
rect 22235 31260 22247 31263
rect 22462 31260 22468 31272
rect 22235 31232 22468 31260
rect 22235 31229 22247 31232
rect 22189 31223 22247 31229
rect 22462 31220 22468 31232
rect 22520 31260 22526 31272
rect 23676 31260 23704 31291
rect 26326 31288 26332 31300
rect 26384 31288 26390 31340
rect 31570 31288 31576 31340
rect 31628 31328 31634 31340
rect 32968 31337 32996 31368
rect 33502 31356 33508 31368
rect 33560 31356 33566 31408
rect 34790 31396 34796 31408
rect 34454 31368 34796 31396
rect 34790 31356 34796 31368
rect 34848 31356 34854 31408
rect 46106 31396 46112 31408
rect 46067 31368 46112 31396
rect 46106 31356 46112 31368
rect 46164 31356 46170 31408
rect 32953 31331 33011 31337
rect 32953 31328 32965 31331
rect 31628 31300 32965 31328
rect 31628 31288 31634 31300
rect 32953 31297 32965 31300
rect 32999 31297 33011 31331
rect 32953 31291 33011 31297
rect 22520 31232 23704 31260
rect 24397 31263 24455 31269
rect 22520 31220 22526 31232
rect 24397 31229 24409 31263
rect 24443 31260 24455 31263
rect 24486 31260 24492 31272
rect 24443 31232 24492 31260
rect 24443 31229 24455 31232
rect 24397 31223 24455 31229
rect 24486 31220 24492 31232
rect 24544 31220 24550 31272
rect 33226 31260 33232 31272
rect 33187 31232 33232 31260
rect 33226 31220 33232 31232
rect 33284 31220 33290 31272
rect 46014 31260 46020 31272
rect 45975 31232 46020 31260
rect 46014 31220 46020 31232
rect 46072 31220 46078 31272
rect 46845 31263 46903 31269
rect 46845 31229 46857 31263
rect 46891 31260 46903 31263
rect 47026 31260 47032 31272
rect 46891 31232 47032 31260
rect 46891 31229 46903 31232
rect 46845 31223 46903 31229
rect 47026 31220 47032 31232
rect 47084 31220 47090 31272
rect 22278 31152 22284 31204
rect 22336 31192 22342 31204
rect 22738 31192 22744 31204
rect 22336 31164 22744 31192
rect 22336 31152 22342 31164
rect 22738 31152 22744 31164
rect 22796 31192 22802 31204
rect 22796 31164 24256 31192
rect 22796 31152 22802 31164
rect 10778 31084 10784 31136
rect 10836 31124 10842 31136
rect 10873 31127 10931 31133
rect 10873 31124 10885 31127
rect 10836 31096 10885 31124
rect 10836 31084 10842 31096
rect 10873 31093 10885 31096
rect 10919 31093 10931 31127
rect 12342 31124 12348 31136
rect 12303 31096 12348 31124
rect 10873 31087 10931 31093
rect 12342 31084 12348 31096
rect 12400 31084 12406 31136
rect 16666 31084 16672 31136
rect 16724 31124 16730 31136
rect 16761 31127 16819 31133
rect 16761 31124 16773 31127
rect 16724 31096 16773 31124
rect 16724 31084 16730 31096
rect 16761 31093 16773 31096
rect 16807 31093 16819 31127
rect 21174 31124 21180 31136
rect 21135 31096 21180 31124
rect 16761 31087 16819 31093
rect 21174 31084 21180 31096
rect 21232 31084 21238 31136
rect 21726 31084 21732 31136
rect 21784 31124 21790 31136
rect 23201 31127 23259 31133
rect 23201 31124 23213 31127
rect 21784 31096 23213 31124
rect 21784 31084 21790 31096
rect 23201 31093 23213 31096
rect 23247 31093 23259 31127
rect 24228 31124 24256 31164
rect 24946 31124 24952 31136
rect 24228 31096 24952 31124
rect 23201 31087 23259 31093
rect 24946 31084 24952 31096
rect 25004 31084 25010 31136
rect 25869 31127 25927 31133
rect 25869 31093 25881 31127
rect 25915 31124 25927 31127
rect 26050 31124 26056 31136
rect 25915 31096 26056 31124
rect 25915 31093 25927 31096
rect 25869 31087 25927 31093
rect 26050 31084 26056 31096
rect 26108 31084 26114 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 20993 30923 21051 30929
rect 20993 30889 21005 30923
rect 21039 30920 21051 30923
rect 21358 30920 21364 30932
rect 21039 30892 21364 30920
rect 21039 30889 21051 30892
rect 20993 30883 21051 30889
rect 21358 30880 21364 30892
rect 21416 30880 21422 30932
rect 22281 30923 22339 30929
rect 22281 30889 22293 30923
rect 22327 30920 22339 30923
rect 22925 30923 22983 30929
rect 22925 30920 22937 30923
rect 22327 30892 22937 30920
rect 22327 30889 22339 30892
rect 22281 30883 22339 30889
rect 22925 30889 22937 30892
rect 22971 30889 22983 30923
rect 25682 30920 25688 30932
rect 25643 30892 25688 30920
rect 22925 30883 22983 30889
rect 25682 30880 25688 30892
rect 25740 30880 25746 30932
rect 26326 30920 26332 30932
rect 26287 30892 26332 30920
rect 26326 30880 26332 30892
rect 26384 30880 26390 30932
rect 26786 30880 26792 30932
rect 26844 30920 26850 30932
rect 28537 30923 28595 30929
rect 28537 30920 28549 30923
rect 26844 30892 28549 30920
rect 26844 30880 26850 30892
rect 28537 30889 28549 30892
rect 28583 30889 28595 30923
rect 28537 30883 28595 30889
rect 28994 30880 29000 30932
rect 29052 30920 29058 30932
rect 29549 30923 29607 30929
rect 29549 30920 29561 30923
rect 29052 30892 29561 30920
rect 29052 30880 29058 30892
rect 29549 30889 29561 30892
rect 29595 30889 29607 30923
rect 29549 30883 29607 30889
rect 29638 30880 29644 30932
rect 29696 30920 29702 30932
rect 30009 30923 30067 30929
rect 30009 30920 30021 30923
rect 29696 30892 30021 30920
rect 29696 30880 29702 30892
rect 30009 30889 30021 30892
rect 30055 30889 30067 30923
rect 30009 30883 30067 30889
rect 12986 30852 12992 30864
rect 12947 30824 12992 30852
rect 12986 30812 12992 30824
rect 13044 30812 13050 30864
rect 21542 30812 21548 30864
rect 21600 30852 21606 30864
rect 23293 30855 23351 30861
rect 23293 30852 23305 30855
rect 21600 30824 23305 30852
rect 21600 30812 21606 30824
rect 23293 30821 23305 30824
rect 23339 30821 23351 30855
rect 35802 30852 35808 30864
rect 23293 30815 23351 30821
rect 26252 30824 31754 30852
rect 10778 30784 10784 30796
rect 10739 30756 10784 30784
rect 10778 30744 10784 30756
rect 10836 30744 10842 30796
rect 14274 30744 14280 30796
rect 14332 30784 14338 30796
rect 14645 30787 14703 30793
rect 14645 30784 14657 30787
rect 14332 30756 14657 30784
rect 14332 30744 14338 30756
rect 14645 30753 14657 30756
rect 14691 30753 14703 30787
rect 17405 30787 17463 30793
rect 17405 30784 17417 30787
rect 14645 30747 14703 30753
rect 14752 30756 17417 30784
rect 13265 30719 13323 30725
rect 13265 30685 13277 30719
rect 13311 30716 13323 30719
rect 13538 30716 13544 30728
rect 13311 30688 13544 30716
rect 13311 30685 13323 30688
rect 13265 30679 13323 30685
rect 13538 30676 13544 30688
rect 13596 30676 13602 30728
rect 14366 30676 14372 30728
rect 14424 30716 14430 30728
rect 14752 30725 14780 30756
rect 17405 30753 17417 30756
rect 17451 30753 17463 30787
rect 17405 30747 17463 30753
rect 18874 30744 18880 30796
rect 18932 30784 18938 30796
rect 19245 30787 19303 30793
rect 19245 30784 19257 30787
rect 18932 30756 19257 30784
rect 18932 30744 18938 30756
rect 19245 30753 19257 30756
rect 19291 30784 19303 30787
rect 20070 30784 20076 30796
rect 19291 30756 20076 30784
rect 19291 30753 19303 30756
rect 19245 30747 19303 30753
rect 20070 30744 20076 30756
rect 20128 30744 20134 30796
rect 25501 30787 25559 30793
rect 25501 30753 25513 30787
rect 25547 30784 25559 30787
rect 26142 30784 26148 30796
rect 25547 30756 26148 30784
rect 25547 30753 25559 30756
rect 25501 30747 25559 30753
rect 26142 30744 26148 30756
rect 26200 30744 26206 30796
rect 26252 30728 26280 30824
rect 28534 30744 28540 30796
rect 28592 30784 28598 30796
rect 29641 30787 29699 30793
rect 29641 30784 29653 30787
rect 28592 30756 29653 30784
rect 28592 30744 28598 30756
rect 29641 30753 29653 30756
rect 29687 30753 29699 30787
rect 31386 30784 31392 30796
rect 29641 30747 29699 30753
rect 29840 30756 31392 30784
rect 14737 30719 14795 30725
rect 14737 30716 14749 30719
rect 14424 30688 14749 30716
rect 14424 30676 14430 30688
rect 14737 30685 14749 30688
rect 14783 30685 14795 30719
rect 15654 30716 15660 30728
rect 15615 30688 15660 30716
rect 14737 30679 14795 30685
rect 15654 30676 15660 30688
rect 15712 30676 15718 30728
rect 21174 30716 21180 30728
rect 20654 30688 21180 30716
rect 21174 30676 21180 30688
rect 21232 30676 21238 30728
rect 21913 30719 21971 30725
rect 21913 30685 21925 30719
rect 21959 30716 21971 30719
rect 22278 30716 22284 30728
rect 21959 30688 22094 30716
rect 22239 30688 22284 30716
rect 21959 30685 21971 30688
rect 21913 30679 21971 30685
rect 11054 30648 11060 30660
rect 11015 30620 11060 30648
rect 11054 30608 11060 30620
rect 11112 30608 11118 30660
rect 12342 30648 12348 30660
rect 12282 30620 12348 30648
rect 12342 30608 12348 30620
rect 12400 30608 12406 30660
rect 13354 30648 13360 30660
rect 13315 30620 13360 30648
rect 13354 30608 13360 30620
rect 13412 30608 13418 30660
rect 15933 30651 15991 30657
rect 15933 30617 15945 30651
rect 15979 30617 15991 30651
rect 15933 30611 15991 30617
rect 12529 30583 12587 30589
rect 12529 30549 12541 30583
rect 12575 30580 12587 30583
rect 12618 30580 12624 30592
rect 12575 30552 12624 30580
rect 12575 30549 12587 30552
rect 12529 30543 12587 30549
rect 12618 30540 12624 30552
rect 12676 30580 12682 30592
rect 13173 30583 13231 30589
rect 13173 30580 13185 30583
rect 12676 30552 13185 30580
rect 12676 30540 12682 30552
rect 13173 30549 13185 30552
rect 13219 30549 13231 30583
rect 13173 30543 13231 30549
rect 13541 30583 13599 30589
rect 13541 30549 13553 30583
rect 13587 30580 13599 30583
rect 14182 30580 14188 30592
rect 13587 30552 14188 30580
rect 13587 30549 13599 30552
rect 13541 30543 13599 30549
rect 14182 30540 14188 30552
rect 14240 30540 14246 30592
rect 15105 30583 15163 30589
rect 15105 30549 15117 30583
rect 15151 30580 15163 30583
rect 15948 30580 15976 30611
rect 16666 30608 16672 30660
rect 16724 30608 16730 30660
rect 19521 30651 19579 30657
rect 19521 30617 19533 30651
rect 19567 30617 19579 30651
rect 21358 30648 21364 30660
rect 19521 30611 19579 30617
rect 20916 30620 21364 30648
rect 15151 30552 15976 30580
rect 19536 30580 19564 30611
rect 20916 30580 20944 30620
rect 21358 30608 21364 30620
rect 21416 30608 21422 30660
rect 22066 30648 22094 30688
rect 22278 30676 22284 30688
rect 22336 30676 22342 30728
rect 22370 30676 22376 30728
rect 22428 30716 22434 30728
rect 23109 30719 23167 30725
rect 23109 30716 23121 30719
rect 22428 30688 23121 30716
rect 22428 30676 22434 30688
rect 23109 30685 23121 30688
rect 23155 30685 23167 30719
rect 23109 30679 23167 30685
rect 23382 30676 23388 30728
rect 23440 30716 23446 30728
rect 25409 30719 25467 30725
rect 23440 30688 23485 30716
rect 23440 30676 23446 30688
rect 25409 30685 25421 30719
rect 25455 30716 25467 30719
rect 26050 30716 26056 30728
rect 25455 30688 26056 30716
rect 25455 30685 25467 30688
rect 25409 30679 25467 30685
rect 26050 30676 26056 30688
rect 26108 30676 26114 30728
rect 26234 30676 26240 30728
rect 26292 30716 26298 30728
rect 28169 30719 28227 30725
rect 26292 30688 26385 30716
rect 26292 30676 26298 30688
rect 28169 30685 28181 30719
rect 28215 30716 28227 30719
rect 28718 30716 28724 30728
rect 28215 30688 28724 30716
rect 28215 30685 28227 30688
rect 28169 30679 28227 30685
rect 28718 30676 28724 30688
rect 28776 30676 28782 30728
rect 29840 30725 29868 30756
rect 31386 30744 31392 30756
rect 31444 30744 31450 30796
rect 31726 30784 31754 30824
rect 32140 30824 35808 30852
rect 32140 30784 32168 30824
rect 35802 30812 35808 30824
rect 35860 30812 35866 30864
rect 31726 30756 32168 30784
rect 29825 30719 29883 30725
rect 29825 30685 29837 30719
rect 29871 30685 29883 30719
rect 29825 30679 29883 30685
rect 30466 30676 30472 30728
rect 30524 30716 30530 30728
rect 30561 30719 30619 30725
rect 30561 30716 30573 30719
rect 30524 30688 30573 30716
rect 30524 30676 30530 30688
rect 30561 30685 30573 30688
rect 30607 30685 30619 30719
rect 30561 30679 30619 30685
rect 30745 30719 30803 30725
rect 30745 30685 30757 30719
rect 30791 30716 30803 30719
rect 31018 30716 31024 30728
rect 30791 30688 31024 30716
rect 30791 30685 30803 30688
rect 30745 30679 30803 30685
rect 31018 30676 31024 30688
rect 31076 30716 31082 30728
rect 31294 30716 31300 30728
rect 31076 30688 31300 30716
rect 31076 30676 31082 30688
rect 31294 30676 31300 30688
rect 31352 30676 31358 30728
rect 32140 30725 32168 30756
rect 34514 30744 34520 30796
rect 34572 30784 34578 30796
rect 35253 30787 35311 30793
rect 34572 30756 35112 30784
rect 34572 30744 34578 30756
rect 32125 30719 32183 30725
rect 32125 30685 32137 30719
rect 32171 30685 32183 30719
rect 33778 30716 33784 30728
rect 33739 30688 33784 30716
rect 32125 30679 32183 30685
rect 33778 30676 33784 30688
rect 33836 30676 33842 30728
rect 35084 30725 35112 30756
rect 35253 30753 35265 30787
rect 35299 30784 35311 30787
rect 44358 30784 44364 30796
rect 35299 30756 44364 30784
rect 35299 30753 35311 30756
rect 35253 30747 35311 30753
rect 44358 30744 44364 30756
rect 44416 30744 44422 30796
rect 34149 30719 34207 30725
rect 34149 30685 34161 30719
rect 34195 30716 34207 30719
rect 34885 30719 34943 30725
rect 34885 30716 34897 30719
rect 34195 30688 34897 30716
rect 34195 30685 34207 30688
rect 34149 30679 34207 30685
rect 34885 30685 34897 30688
rect 34931 30685 34943 30719
rect 34885 30679 34943 30685
rect 35069 30719 35127 30725
rect 35069 30685 35081 30719
rect 35115 30685 35127 30719
rect 35069 30679 35127 30685
rect 35158 30676 35164 30728
rect 35216 30716 35222 30728
rect 35434 30716 35440 30728
rect 35216 30688 35261 30716
rect 35347 30688 35440 30716
rect 35216 30676 35222 30688
rect 35434 30676 35440 30688
rect 35492 30676 35498 30728
rect 22554 30648 22560 30660
rect 22066 30620 22560 30648
rect 22554 30608 22560 30620
rect 22612 30608 22618 30660
rect 24581 30651 24639 30657
rect 24581 30617 24593 30651
rect 24627 30648 24639 30651
rect 24854 30648 24860 30660
rect 24627 30620 24860 30648
rect 24627 30617 24639 30620
rect 24581 30611 24639 30617
rect 24854 30608 24860 30620
rect 24912 30608 24918 30660
rect 28353 30651 28411 30657
rect 28353 30617 28365 30651
rect 28399 30648 28411 30651
rect 28626 30648 28632 30660
rect 28399 30620 28632 30648
rect 28399 30617 28411 30620
rect 28353 30611 28411 30617
rect 28626 30608 28632 30620
rect 28684 30608 28690 30660
rect 29549 30651 29607 30657
rect 29549 30617 29561 30651
rect 29595 30648 29607 30651
rect 31110 30648 31116 30660
rect 29595 30620 31116 30648
rect 29595 30617 29607 30620
rect 29549 30611 29607 30617
rect 31110 30608 31116 30620
rect 31168 30608 31174 30660
rect 31481 30651 31539 30657
rect 31481 30617 31493 30651
rect 31527 30648 31539 30651
rect 32306 30648 32312 30660
rect 31527 30620 32312 30648
rect 31527 30617 31539 30620
rect 31481 30611 31539 30617
rect 32306 30608 32312 30620
rect 32364 30608 32370 30660
rect 33965 30651 34023 30657
rect 33965 30617 33977 30651
rect 34011 30617 34023 30651
rect 33965 30611 34023 30617
rect 19536 30552 20944 30580
rect 15151 30549 15163 30552
rect 15105 30543 15163 30549
rect 21910 30540 21916 30592
rect 21968 30580 21974 30592
rect 22465 30583 22523 30589
rect 22465 30580 22477 30583
rect 21968 30552 22477 30580
rect 21968 30540 21974 30552
rect 22465 30549 22477 30552
rect 22511 30549 22523 30583
rect 24670 30580 24676 30592
rect 24631 30552 24676 30580
rect 22465 30543 22523 30549
rect 24670 30540 24676 30552
rect 24728 30540 24734 30592
rect 30650 30580 30656 30592
rect 30611 30552 30656 30580
rect 30650 30540 30656 30552
rect 30708 30540 30714 30592
rect 31570 30580 31576 30592
rect 31531 30552 31576 30580
rect 31570 30540 31576 30552
rect 31628 30540 31634 30592
rect 32214 30580 32220 30592
rect 32175 30552 32220 30580
rect 32214 30540 32220 30552
rect 32272 30540 32278 30592
rect 33980 30580 34008 30611
rect 34514 30608 34520 30660
rect 34572 30648 34578 30660
rect 35452 30648 35480 30676
rect 34572 30620 35480 30648
rect 34572 30608 34578 30620
rect 34146 30580 34152 30592
rect 33980 30552 34152 30580
rect 34146 30540 34152 30552
rect 34204 30540 34210 30592
rect 35250 30540 35256 30592
rect 35308 30580 35314 30592
rect 35621 30583 35679 30589
rect 35621 30580 35633 30583
rect 35308 30552 35633 30580
rect 35308 30540 35314 30552
rect 35621 30549 35633 30552
rect 35667 30549 35679 30583
rect 35621 30543 35679 30549
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 11054 30336 11060 30388
rect 11112 30376 11118 30388
rect 11701 30379 11759 30385
rect 11701 30376 11713 30379
rect 11112 30348 11713 30376
rect 11112 30336 11118 30348
rect 11701 30345 11713 30348
rect 11747 30345 11759 30379
rect 12618 30376 12624 30388
rect 11701 30339 11759 30345
rect 12406 30348 12624 30376
rect 12253 30311 12311 30317
rect 12253 30308 12265 30311
rect 10980 30280 12265 30308
rect 10980 30252 11008 30280
rect 12253 30277 12265 30280
rect 12299 30308 12311 30311
rect 12406 30308 12434 30348
rect 12618 30336 12624 30348
rect 12676 30336 12682 30388
rect 14274 30376 14280 30388
rect 14235 30348 14280 30376
rect 14274 30336 14280 30348
rect 14332 30336 14338 30388
rect 15654 30336 15660 30388
rect 15712 30376 15718 30388
rect 15749 30379 15807 30385
rect 15749 30376 15761 30379
rect 15712 30348 15761 30376
rect 15712 30336 15718 30348
rect 15749 30345 15761 30348
rect 15795 30345 15807 30379
rect 15749 30339 15807 30345
rect 21450 30336 21456 30388
rect 21508 30376 21514 30388
rect 22370 30376 22376 30388
rect 21508 30348 22376 30376
rect 21508 30336 21514 30348
rect 22370 30336 22376 30348
rect 22428 30336 22434 30388
rect 24305 30379 24363 30385
rect 24305 30345 24317 30379
rect 24351 30345 24363 30379
rect 31570 30376 31576 30388
rect 24305 30339 24363 30345
rect 30484 30348 31576 30376
rect 12299 30280 12434 30308
rect 12529 30311 12587 30317
rect 12299 30277 12311 30280
rect 12253 30271 12311 30277
rect 12529 30277 12541 30311
rect 12575 30308 12587 30311
rect 12710 30308 12716 30320
rect 12575 30280 12716 30308
rect 12575 30277 12587 30280
rect 12529 30271 12587 30277
rect 12710 30268 12716 30280
rect 12768 30308 12774 30320
rect 13354 30308 13360 30320
rect 12768 30280 13360 30308
rect 12768 30268 12774 30280
rect 13354 30268 13360 30280
rect 13412 30268 13418 30320
rect 20622 30268 20628 30320
rect 20680 30308 20686 30320
rect 21177 30311 21235 30317
rect 21177 30308 21189 30311
rect 20680 30280 21189 30308
rect 20680 30268 20686 30280
rect 21177 30277 21189 30280
rect 21223 30277 21235 30311
rect 21177 30271 21235 30277
rect 21818 30268 21824 30320
rect 21876 30308 21882 30320
rect 23014 30308 23020 30320
rect 21876 30280 23020 30308
rect 21876 30268 21882 30280
rect 10594 30240 10600 30252
rect 10555 30212 10600 30240
rect 10594 30200 10600 30212
rect 10652 30200 10658 30252
rect 10686 30200 10692 30252
rect 10744 30240 10750 30252
rect 10962 30240 10968 30252
rect 10744 30212 10789 30240
rect 10923 30212 10968 30240
rect 10744 30200 10750 30212
rect 10962 30200 10968 30212
rect 11020 30200 11026 30252
rect 11609 30243 11667 30249
rect 11609 30209 11621 30243
rect 11655 30209 11667 30243
rect 11609 30203 11667 30209
rect 11793 30243 11851 30249
rect 11793 30209 11805 30243
rect 11839 30209 11851 30243
rect 11793 30203 11851 30209
rect 10781 30175 10839 30181
rect 10781 30141 10793 30175
rect 10827 30141 10839 30175
rect 11624 30172 11652 30203
rect 10781 30135 10839 30141
rect 10980 30144 11652 30172
rect 11808 30172 11836 30203
rect 12434 30200 12440 30252
rect 12492 30240 12498 30252
rect 12621 30243 12679 30249
rect 12492 30212 12537 30240
rect 12492 30200 12498 30212
rect 12621 30209 12633 30243
rect 12667 30240 12679 30243
rect 13170 30240 13176 30252
rect 12667 30212 13176 30240
rect 12667 30209 12679 30212
rect 12621 30203 12679 30209
rect 13170 30200 13176 30212
rect 13228 30240 13234 30252
rect 14093 30243 14151 30249
rect 14093 30240 14105 30243
rect 13228 30212 14105 30240
rect 13228 30200 13234 30212
rect 14093 30209 14105 30212
rect 14139 30209 14151 30243
rect 14093 30203 14151 30209
rect 14182 30200 14188 30252
rect 14240 30240 14246 30252
rect 14277 30243 14335 30249
rect 14277 30240 14289 30243
rect 14240 30212 14289 30240
rect 14240 30200 14246 30212
rect 14277 30209 14289 30212
rect 14323 30209 14335 30243
rect 14277 30203 14335 30209
rect 15286 30200 15292 30252
rect 15344 30240 15350 30252
rect 15565 30243 15623 30249
rect 15565 30240 15577 30243
rect 15344 30212 15577 30240
rect 15344 30200 15350 30212
rect 15565 30209 15577 30212
rect 15611 30209 15623 30243
rect 20898 30240 20904 30252
rect 20859 30212 20904 30240
rect 15565 30203 15623 30209
rect 20898 30200 20904 30212
rect 20956 30200 20962 30252
rect 20993 30243 21051 30249
rect 20993 30209 21005 30243
rect 21039 30240 21051 30243
rect 21726 30240 21732 30252
rect 21039 30212 21732 30240
rect 21039 30209 21051 30212
rect 20993 30203 21051 30209
rect 21726 30200 21732 30212
rect 21784 30200 21790 30252
rect 21910 30240 21916 30252
rect 21871 30212 21916 30240
rect 21910 30200 21916 30212
rect 21968 30200 21974 30252
rect 22112 30249 22140 30280
rect 23014 30268 23020 30280
rect 23072 30268 23078 30320
rect 24320 30308 24348 30339
rect 25682 30308 25688 30320
rect 23768 30280 24348 30308
rect 24688 30280 25688 30308
rect 22097 30243 22155 30249
rect 22097 30209 22109 30243
rect 22143 30209 22155 30243
rect 22097 30203 22155 30209
rect 22189 30243 22247 30249
rect 22189 30209 22201 30243
rect 22235 30240 22247 30243
rect 22370 30240 22376 30252
rect 22235 30212 22376 30240
rect 22235 30209 22247 30212
rect 22189 30203 22247 30209
rect 22370 30200 22376 30212
rect 22428 30200 22434 30252
rect 22465 30243 22523 30249
rect 22465 30209 22477 30243
rect 22511 30240 22523 30243
rect 22646 30240 22652 30252
rect 22511 30212 22652 30240
rect 22511 30209 22523 30212
rect 22465 30203 22523 30209
rect 22646 30200 22652 30212
rect 22704 30200 22710 30252
rect 12805 30175 12863 30181
rect 12805 30172 12817 30175
rect 11808 30144 12817 30172
rect 10796 30036 10824 30135
rect 10980 30113 11008 30144
rect 12805 30141 12817 30144
rect 12851 30172 12863 30175
rect 14458 30172 14464 30184
rect 12851 30144 14464 30172
rect 12851 30141 12863 30144
rect 12805 30135 12863 30141
rect 14458 30132 14464 30144
rect 14516 30132 14522 30184
rect 20530 30172 20536 30184
rect 20491 30144 20536 30172
rect 20530 30132 20536 30144
rect 20588 30132 20594 30184
rect 22278 30132 22284 30184
rect 22336 30172 22342 30184
rect 22336 30144 22381 30172
rect 22336 30132 22342 30144
rect 10965 30107 11023 30113
rect 10965 30073 10977 30107
rect 11011 30073 11023 30107
rect 10965 30067 11023 30073
rect 17126 30064 17132 30116
rect 17184 30104 17190 30116
rect 17184 30076 21312 30104
rect 17184 30064 17190 30076
rect 12434 30036 12440 30048
rect 10796 30008 12440 30036
rect 12434 29996 12440 30008
rect 12492 29996 12498 30048
rect 21284 30036 21312 30076
rect 21358 30064 21364 30116
rect 21416 30104 21422 30116
rect 22649 30107 22707 30113
rect 22649 30104 22661 30107
rect 21416 30076 22661 30104
rect 21416 30064 21422 30076
rect 22649 30073 22661 30076
rect 22695 30073 22707 30107
rect 22649 30067 22707 30073
rect 23768 30045 23796 30280
rect 24210 30200 24216 30252
rect 24268 30249 24274 30252
rect 24688 30249 24716 30280
rect 25682 30268 25688 30280
rect 25740 30268 25746 30320
rect 25958 30268 25964 30320
rect 26016 30308 26022 30320
rect 26237 30311 26295 30317
rect 26237 30308 26249 30311
rect 26016 30280 26249 30308
rect 26016 30268 26022 30280
rect 26237 30277 26249 30280
rect 26283 30277 26295 30311
rect 26237 30271 26295 30277
rect 27706 30268 27712 30320
rect 27764 30308 27770 30320
rect 28166 30308 28172 30320
rect 27764 30280 28172 30308
rect 27764 30268 27770 30280
rect 28166 30268 28172 30280
rect 28224 30268 28230 30320
rect 30484 30308 30512 30348
rect 31570 30336 31576 30348
rect 31628 30336 31634 30388
rect 34517 30379 34575 30385
rect 34517 30345 34529 30379
rect 34563 30376 34575 30379
rect 35158 30376 35164 30388
rect 34563 30348 35164 30376
rect 34563 30345 34575 30348
rect 34517 30339 34575 30345
rect 35158 30336 35164 30348
rect 35216 30336 35222 30388
rect 32214 30308 32220 30320
rect 29840 30280 30512 30308
rect 31326 30280 32220 30308
rect 24268 30243 24304 30249
rect 24292 30209 24304 30243
rect 24268 30203 24304 30209
rect 24673 30243 24731 30249
rect 24673 30209 24685 30243
rect 24719 30209 24731 30243
rect 25406 30240 25412 30252
rect 25367 30212 25412 30240
rect 24673 30203 24731 30209
rect 24268 30200 24274 30203
rect 25406 30200 25412 30212
rect 25464 30200 25470 30252
rect 26050 30240 26056 30252
rect 26011 30212 26056 30240
rect 26050 30200 26056 30212
rect 26108 30200 26114 30252
rect 27522 30240 27528 30252
rect 27483 30212 27528 30240
rect 27522 30200 27528 30212
rect 27580 30240 27586 30252
rect 28537 30243 28595 30249
rect 27580 30212 28488 30240
rect 27580 30200 27586 30212
rect 24762 30172 24768 30184
rect 24723 30144 24768 30172
rect 24762 30132 24768 30144
rect 24820 30132 24826 30184
rect 25038 30132 25044 30184
rect 25096 30172 25102 30184
rect 27433 30175 27491 30181
rect 27433 30172 27445 30175
rect 25096 30144 27445 30172
rect 25096 30132 25102 30144
rect 27433 30141 27445 30144
rect 27479 30172 27491 30175
rect 28166 30172 28172 30184
rect 27479 30144 28172 30172
rect 27479 30141 27491 30144
rect 27433 30135 27491 30141
rect 28166 30132 28172 30144
rect 28224 30132 28230 30184
rect 28460 30172 28488 30212
rect 28537 30209 28549 30243
rect 28583 30240 28595 30243
rect 28994 30240 29000 30252
rect 28583 30212 29000 30240
rect 28583 30209 28595 30212
rect 28537 30203 28595 30209
rect 28994 30200 29000 30212
rect 29052 30200 29058 30252
rect 29840 30249 29868 30280
rect 32214 30268 32220 30280
rect 32272 30268 32278 30320
rect 33137 30311 33195 30317
rect 33137 30277 33149 30311
rect 33183 30308 33195 30311
rect 33183 30280 33456 30308
rect 33183 30277 33195 30280
rect 33137 30271 33195 30277
rect 29825 30243 29883 30249
rect 29825 30209 29837 30243
rect 29871 30209 29883 30243
rect 33318 30240 33324 30252
rect 33279 30212 33324 30240
rect 29825 30203 29883 30209
rect 33318 30200 33324 30212
rect 33376 30200 33382 30252
rect 33428 30240 33456 30280
rect 33502 30268 33508 30320
rect 33560 30308 33566 30320
rect 35250 30308 35256 30320
rect 33560 30280 34284 30308
rect 35211 30280 35256 30308
rect 33560 30268 33566 30280
rect 34146 30240 34152 30252
rect 33428 30212 34152 30240
rect 34146 30200 34152 30212
rect 34204 30200 34210 30252
rect 34256 30184 34284 30280
rect 35250 30268 35256 30280
rect 35308 30268 35314 30320
rect 35894 30268 35900 30320
rect 35952 30268 35958 30320
rect 28813 30175 28871 30181
rect 28813 30172 28825 30175
rect 28460 30144 28825 30172
rect 28813 30141 28825 30144
rect 28859 30141 28871 30175
rect 28813 30135 28871 30141
rect 30101 30175 30159 30181
rect 30101 30141 30113 30175
rect 30147 30172 30159 30175
rect 30558 30172 30564 30184
rect 30147 30144 30564 30172
rect 30147 30141 30159 30144
rect 30101 30135 30159 30141
rect 30558 30132 30564 30144
rect 30616 30132 30622 30184
rect 31294 30132 31300 30184
rect 31352 30172 31358 30184
rect 34057 30175 34115 30181
rect 34057 30172 34069 30175
rect 31352 30144 34069 30172
rect 31352 30132 31358 30144
rect 34057 30141 34069 30144
rect 34103 30141 34115 30175
rect 34057 30135 34115 30141
rect 34238 30132 34244 30184
rect 34296 30172 34302 30184
rect 34977 30175 35035 30181
rect 34977 30172 34989 30175
rect 34296 30144 34989 30172
rect 34296 30132 34302 30144
rect 34977 30141 34989 30144
rect 35023 30141 35035 30175
rect 34977 30135 35035 30141
rect 24118 30104 24124 30116
rect 24079 30076 24124 30104
rect 24118 30064 24124 30076
rect 24176 30064 24182 30116
rect 24780 30104 24808 30132
rect 26421 30107 26479 30113
rect 24780 30076 26372 30104
rect 23753 30039 23811 30045
rect 23753 30036 23765 30039
rect 21284 30008 23765 30036
rect 23753 30005 23765 30008
rect 23799 30005 23811 30039
rect 23753 29999 23811 30005
rect 24854 29996 24860 30048
rect 24912 30036 24918 30048
rect 25501 30039 25559 30045
rect 25501 30036 25513 30039
rect 24912 30008 25513 30036
rect 24912 29996 24918 30008
rect 25501 30005 25513 30008
rect 25547 30005 25559 30039
rect 26344 30036 26372 30076
rect 26421 30073 26433 30107
rect 26467 30104 26479 30107
rect 28534 30104 28540 30116
rect 26467 30076 28540 30104
rect 26467 30073 26479 30076
rect 26421 30067 26479 30073
rect 28534 30064 28540 30076
rect 28592 30064 28598 30116
rect 31110 30064 31116 30116
rect 31168 30104 31174 30116
rect 34790 30104 34796 30116
rect 31168 30076 34796 30104
rect 31168 30064 31174 30076
rect 34790 30064 34796 30076
rect 34848 30064 34854 30116
rect 26602 30036 26608 30048
rect 26344 30008 26608 30036
rect 25501 29999 25559 30005
rect 26602 29996 26608 30008
rect 26660 29996 26666 30048
rect 27614 29996 27620 30048
rect 27672 30036 27678 30048
rect 27893 30039 27951 30045
rect 27893 30036 27905 30039
rect 27672 30008 27905 30036
rect 27672 29996 27678 30008
rect 27893 30005 27905 30008
rect 27939 30005 27951 30039
rect 27893 29999 27951 30005
rect 31386 29996 31392 30048
rect 31444 30036 31450 30048
rect 31573 30039 31631 30045
rect 31573 30036 31585 30039
rect 31444 30008 31585 30036
rect 31444 29996 31450 30008
rect 31573 30005 31585 30008
rect 31619 30005 31631 30039
rect 31573 29999 31631 30005
rect 31662 29996 31668 30048
rect 31720 30036 31726 30048
rect 33505 30039 33563 30045
rect 33505 30036 33517 30039
rect 31720 30008 33517 30036
rect 31720 29996 31726 30008
rect 33505 30005 33517 30008
rect 33551 30005 33563 30039
rect 33505 29999 33563 30005
rect 34146 29996 34152 30048
rect 34204 30036 34210 30048
rect 34422 30036 34428 30048
rect 34204 30008 34428 30036
rect 34204 29996 34210 30008
rect 34422 29996 34428 30008
rect 34480 30036 34486 30048
rect 36725 30039 36783 30045
rect 36725 30036 36737 30039
rect 34480 30008 36737 30036
rect 34480 29996 34486 30008
rect 36725 30005 36737 30008
rect 36771 30005 36783 30039
rect 36725 29999 36783 30005
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 9306 29792 9312 29844
rect 9364 29832 9370 29844
rect 17126 29832 17132 29844
rect 9364 29804 17132 29832
rect 9364 29792 9370 29804
rect 17126 29792 17132 29804
rect 17184 29792 17190 29844
rect 20530 29792 20536 29844
rect 20588 29832 20594 29844
rect 21269 29835 21327 29841
rect 21269 29832 21281 29835
rect 20588 29804 21281 29832
rect 20588 29792 20594 29804
rect 21269 29801 21281 29804
rect 21315 29801 21327 29835
rect 21269 29795 21327 29801
rect 21542 29792 21548 29844
rect 21600 29832 21606 29844
rect 21821 29835 21879 29841
rect 21821 29832 21833 29835
rect 21600 29804 21833 29832
rect 21600 29792 21606 29804
rect 21821 29801 21833 29804
rect 21867 29801 21879 29835
rect 24762 29832 24768 29844
rect 21821 29795 21879 29801
rect 22940 29804 24768 29832
rect 22940 29764 22968 29804
rect 24762 29792 24768 29804
rect 24820 29792 24826 29844
rect 24946 29832 24952 29844
rect 24907 29804 24952 29832
rect 24946 29792 24952 29804
rect 25004 29792 25010 29844
rect 28994 29832 29000 29844
rect 25056 29804 28580 29832
rect 28955 29804 29000 29832
rect 22066 29736 22968 29764
rect 9309 29699 9367 29705
rect 9309 29665 9321 29699
rect 9355 29696 9367 29699
rect 10962 29696 10968 29708
rect 9355 29668 10968 29696
rect 9355 29665 9367 29668
rect 9309 29659 9367 29665
rect 10962 29656 10968 29668
rect 11020 29656 11026 29708
rect 21913 29699 21971 29705
rect 21913 29665 21925 29699
rect 21959 29696 21971 29699
rect 22066 29696 22094 29736
rect 23014 29724 23020 29776
rect 23072 29764 23078 29776
rect 25056 29764 25084 29804
rect 23072 29736 25084 29764
rect 28552 29764 28580 29804
rect 28994 29792 29000 29804
rect 29052 29792 29058 29844
rect 30558 29832 30564 29844
rect 30519 29804 30564 29832
rect 30558 29792 30564 29804
rect 30616 29792 30622 29844
rect 30742 29792 30748 29844
rect 30800 29832 30806 29844
rect 31021 29835 31079 29841
rect 31021 29832 31033 29835
rect 30800 29804 31033 29832
rect 30800 29792 30806 29804
rect 31021 29801 31033 29804
rect 31067 29801 31079 29835
rect 32125 29835 32183 29841
rect 32125 29832 32137 29835
rect 31021 29795 31079 29801
rect 31128 29804 32137 29832
rect 29546 29764 29552 29776
rect 28552 29736 29552 29764
rect 23072 29724 23078 29736
rect 29546 29724 29552 29736
rect 29604 29724 29610 29776
rect 21959 29668 22094 29696
rect 21959 29665 21971 29668
rect 21913 29659 21971 29665
rect 15286 29588 15292 29640
rect 15344 29628 15350 29640
rect 15381 29631 15439 29637
rect 15381 29628 15393 29631
rect 15344 29600 15393 29628
rect 15344 29588 15350 29600
rect 15381 29597 15393 29600
rect 15427 29597 15439 29631
rect 15381 29591 15439 29597
rect 15657 29631 15715 29637
rect 15657 29597 15669 29631
rect 15703 29628 15715 29631
rect 16117 29631 16175 29637
rect 16117 29628 16129 29631
rect 15703 29600 16129 29628
rect 15703 29597 15715 29600
rect 15657 29591 15715 29597
rect 16117 29597 16129 29600
rect 16163 29597 16175 29631
rect 16117 29591 16175 29597
rect 21450 29631 21508 29637
rect 21450 29597 21462 29631
rect 21496 29628 21508 29631
rect 21496 29600 21772 29628
rect 21496 29597 21508 29600
rect 21450 29591 21508 29597
rect 9493 29563 9551 29569
rect 9493 29529 9505 29563
rect 9539 29560 9551 29563
rect 9674 29560 9680 29572
rect 9539 29532 9680 29560
rect 9539 29529 9551 29532
rect 9493 29523 9551 29529
rect 9674 29520 9680 29532
rect 9732 29520 9738 29572
rect 11149 29563 11207 29569
rect 11149 29560 11161 29563
rect 9784 29532 11161 29560
rect 9030 29452 9036 29504
rect 9088 29492 9094 29504
rect 9784 29492 9812 29532
rect 11149 29529 11161 29532
rect 11195 29529 11207 29563
rect 11149 29523 11207 29529
rect 15746 29520 15752 29572
rect 15804 29560 15810 29572
rect 16393 29563 16451 29569
rect 16393 29560 16405 29563
rect 15804 29532 16405 29560
rect 15804 29520 15810 29532
rect 16393 29529 16405 29532
rect 16439 29529 16451 29563
rect 16393 29523 16451 29529
rect 16942 29520 16948 29572
rect 17000 29520 17006 29572
rect 21744 29560 21772 29600
rect 22094 29588 22100 29640
rect 22152 29628 22158 29640
rect 23032 29628 23060 29724
rect 24670 29656 24676 29708
rect 24728 29696 24734 29708
rect 27249 29699 27307 29705
rect 27249 29696 27261 29699
rect 24728 29668 27261 29696
rect 24728 29656 24734 29668
rect 27249 29665 27261 29668
rect 27295 29665 27307 29699
rect 27249 29659 27307 29665
rect 28810 29656 28816 29708
rect 28868 29696 28874 29708
rect 30101 29699 30159 29705
rect 28868 29668 30052 29696
rect 28868 29656 28874 29668
rect 22152 29600 23060 29628
rect 24765 29631 24823 29637
rect 22152 29588 22158 29600
rect 24765 29597 24777 29631
rect 24811 29628 24823 29631
rect 25038 29628 25044 29640
rect 24811 29600 25044 29628
rect 24811 29597 24823 29600
rect 24765 29591 24823 29597
rect 25038 29588 25044 29600
rect 25096 29588 25102 29640
rect 25133 29631 25191 29637
rect 25133 29597 25145 29631
rect 25179 29628 25191 29631
rect 25777 29631 25835 29637
rect 25777 29628 25789 29631
rect 25179 29600 25789 29628
rect 25179 29597 25191 29600
rect 25133 29591 25191 29597
rect 25777 29597 25789 29600
rect 25823 29597 25835 29631
rect 25958 29628 25964 29640
rect 25919 29600 25964 29628
rect 25777 29591 25835 29597
rect 25958 29588 25964 29600
rect 26016 29588 26022 29640
rect 26142 29628 26148 29640
rect 26103 29600 26148 29628
rect 26142 29588 26148 29600
rect 26200 29588 26206 29640
rect 26237 29631 26295 29637
rect 26237 29597 26249 29631
rect 26283 29597 26295 29631
rect 29822 29628 29828 29640
rect 29783 29600 29828 29628
rect 26237 29591 26295 29597
rect 24210 29560 24216 29572
rect 21744 29532 24216 29560
rect 24210 29520 24216 29532
rect 24268 29560 24274 29572
rect 24486 29560 24492 29572
rect 24268 29532 24492 29560
rect 24268 29520 24274 29532
rect 24486 29520 24492 29532
rect 24544 29520 24550 29572
rect 26050 29520 26056 29572
rect 26108 29560 26114 29572
rect 26252 29560 26280 29591
rect 29822 29588 29828 29600
rect 29880 29588 29886 29640
rect 30024 29637 30052 29668
rect 30101 29665 30113 29699
rect 30147 29696 30159 29699
rect 30650 29696 30656 29708
rect 30147 29668 30656 29696
rect 30147 29665 30159 29668
rect 30101 29659 30159 29665
rect 30650 29656 30656 29668
rect 30708 29656 30714 29708
rect 30009 29631 30067 29637
rect 30009 29597 30021 29631
rect 30055 29597 30067 29631
rect 30009 29591 30067 29597
rect 30193 29631 30251 29637
rect 30193 29597 30205 29631
rect 30239 29597 30251 29631
rect 30374 29628 30380 29640
rect 30335 29600 30380 29628
rect 30193 29591 30251 29597
rect 26108 29532 26280 29560
rect 27525 29563 27583 29569
rect 26108 29520 26114 29532
rect 27525 29529 27537 29563
rect 27571 29560 27583 29563
rect 27798 29560 27804 29572
rect 27571 29532 27804 29560
rect 27571 29529 27583 29532
rect 27525 29523 27583 29529
rect 27798 29520 27804 29532
rect 27856 29520 27862 29572
rect 29270 29560 29276 29572
rect 28750 29532 29276 29560
rect 29270 29520 29276 29532
rect 29328 29520 29334 29572
rect 29730 29520 29736 29572
rect 29788 29560 29794 29572
rect 30208 29560 30236 29591
rect 30374 29588 30380 29600
rect 30432 29588 30438 29640
rect 29788 29532 30236 29560
rect 29788 29520 29794 29532
rect 30650 29520 30656 29572
rect 30708 29560 30714 29572
rect 31021 29563 31079 29569
rect 31021 29560 31033 29563
rect 30708 29532 31033 29560
rect 30708 29520 30714 29532
rect 31021 29529 31033 29532
rect 31067 29529 31079 29563
rect 31021 29523 31079 29529
rect 17862 29492 17868 29504
rect 9088 29464 9812 29492
rect 17823 29464 17868 29492
rect 9088 29452 9094 29464
rect 17862 29452 17868 29464
rect 17920 29452 17926 29504
rect 21450 29492 21456 29504
rect 21411 29464 21456 29492
rect 21450 29452 21456 29464
rect 21508 29452 21514 29504
rect 24762 29452 24768 29504
rect 24820 29492 24826 29504
rect 25317 29495 25375 29501
rect 25317 29492 25329 29495
rect 24820 29464 25329 29492
rect 24820 29452 24826 29464
rect 25317 29461 25329 29464
rect 25363 29461 25375 29495
rect 25317 29455 25375 29461
rect 26602 29452 26608 29504
rect 26660 29492 26666 29504
rect 31128 29492 31156 29804
rect 32125 29801 32137 29804
rect 32171 29801 32183 29835
rect 34698 29832 34704 29844
rect 34659 29804 34704 29832
rect 32125 29795 32183 29801
rect 34698 29792 34704 29804
rect 34756 29792 34762 29844
rect 34790 29792 34796 29844
rect 34848 29832 34854 29844
rect 35161 29835 35219 29841
rect 35161 29832 35173 29835
rect 34848 29804 35173 29832
rect 34848 29792 34854 29804
rect 35161 29801 35173 29804
rect 35207 29801 35219 29835
rect 35894 29832 35900 29844
rect 35855 29804 35900 29832
rect 35161 29795 35219 29801
rect 35894 29792 35900 29804
rect 35952 29792 35958 29844
rect 31481 29767 31539 29773
rect 31481 29733 31493 29767
rect 31527 29764 31539 29767
rect 31527 29736 31754 29764
rect 31527 29733 31539 29736
rect 31481 29727 31539 29733
rect 31205 29699 31263 29705
rect 31205 29665 31217 29699
rect 31251 29696 31263 29699
rect 31570 29696 31576 29708
rect 31251 29668 31576 29696
rect 31251 29665 31263 29668
rect 31205 29659 31263 29665
rect 31570 29656 31576 29668
rect 31628 29656 31634 29708
rect 31297 29631 31355 29637
rect 31297 29597 31309 29631
rect 31343 29628 31355 29631
rect 31386 29628 31392 29640
rect 31343 29600 31392 29628
rect 31343 29597 31355 29600
rect 31297 29591 31355 29597
rect 31386 29588 31392 29600
rect 31444 29588 31450 29640
rect 31726 29628 31754 29736
rect 33318 29696 33324 29708
rect 33231 29668 33324 29696
rect 33318 29656 33324 29668
rect 33376 29696 33382 29708
rect 34882 29696 34888 29708
rect 33376 29668 34888 29696
rect 33376 29656 33382 29668
rect 34882 29656 34888 29668
rect 34940 29656 34946 29708
rect 47210 29656 47216 29708
rect 47268 29696 47274 29708
rect 47581 29699 47639 29705
rect 47581 29696 47593 29699
rect 47268 29668 47593 29696
rect 47268 29656 47274 29668
rect 47581 29665 47593 29668
rect 47627 29665 47639 29699
rect 47581 29659 47639 29665
rect 32030 29628 32036 29640
rect 31726 29600 32036 29628
rect 32030 29588 32036 29600
rect 32088 29588 32094 29640
rect 32398 29628 32404 29640
rect 32359 29600 32404 29628
rect 32398 29588 32404 29600
rect 32456 29588 32462 29640
rect 33045 29631 33103 29637
rect 33045 29628 33057 29631
rect 32600 29600 33057 29628
rect 32600 29501 32628 29600
rect 33045 29597 33057 29600
rect 33091 29597 33103 29631
rect 33045 29591 33103 29597
rect 33134 29588 33140 29640
rect 33192 29628 33198 29640
rect 33229 29631 33287 29637
rect 33229 29628 33241 29631
rect 33192 29600 33241 29628
rect 33192 29588 33198 29600
rect 33229 29597 33241 29600
rect 33275 29597 33287 29631
rect 33229 29591 33287 29597
rect 33413 29631 33471 29637
rect 33413 29597 33425 29631
rect 33459 29597 33471 29631
rect 33413 29591 33471 29597
rect 33597 29631 33655 29637
rect 33597 29597 33609 29631
rect 33643 29628 33655 29631
rect 34514 29628 34520 29640
rect 33643 29600 34520 29628
rect 33643 29597 33655 29600
rect 33597 29591 33655 29597
rect 33318 29520 33324 29572
rect 33376 29560 33382 29572
rect 33428 29560 33456 29591
rect 34514 29588 34520 29600
rect 34572 29588 34578 29640
rect 34606 29588 34612 29640
rect 34664 29628 34670 29640
rect 34977 29631 35035 29637
rect 34977 29628 34989 29631
rect 34664 29600 34989 29628
rect 34664 29588 34670 29600
rect 34977 29597 34989 29600
rect 35023 29597 35035 29631
rect 35802 29628 35808 29640
rect 35763 29600 35808 29628
rect 34977 29591 35035 29597
rect 35802 29588 35808 29600
rect 35860 29588 35866 29640
rect 47305 29631 47363 29637
rect 47305 29597 47317 29631
rect 47351 29628 47363 29631
rect 47394 29628 47400 29640
rect 47351 29600 47400 29628
rect 47351 29597 47363 29600
rect 47305 29591 47363 29597
rect 47394 29588 47400 29600
rect 47452 29588 47458 29640
rect 33376 29532 33456 29560
rect 33376 29520 33382 29532
rect 34422 29520 34428 29572
rect 34480 29560 34486 29572
rect 34701 29563 34759 29569
rect 34701 29560 34713 29563
rect 34480 29532 34713 29560
rect 34480 29520 34486 29532
rect 34701 29529 34713 29532
rect 34747 29529 34759 29563
rect 34701 29523 34759 29529
rect 26660 29464 31156 29492
rect 32585 29495 32643 29501
rect 26660 29452 26666 29464
rect 32585 29461 32597 29495
rect 32631 29461 32643 29495
rect 32585 29455 32643 29461
rect 33781 29495 33839 29501
rect 33781 29461 33793 29495
rect 33827 29492 33839 29495
rect 34514 29492 34520 29504
rect 33827 29464 34520 29492
rect 33827 29461 33839 29464
rect 33781 29455 33839 29461
rect 34514 29452 34520 29464
rect 34572 29452 34578 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 9674 29288 9680 29300
rect 9635 29260 9680 29288
rect 9674 29248 9680 29260
rect 9732 29248 9738 29300
rect 16942 29288 16948 29300
rect 16903 29260 16948 29288
rect 16942 29248 16948 29260
rect 17000 29248 17006 29300
rect 25406 29248 25412 29300
rect 25464 29288 25470 29300
rect 29181 29291 29239 29297
rect 29181 29288 29193 29291
rect 25464 29260 29193 29288
rect 25464 29248 25470 29260
rect 29181 29257 29193 29260
rect 29227 29288 29239 29291
rect 32306 29288 32312 29300
rect 29227 29260 31754 29288
rect 32267 29260 32312 29288
rect 29227 29257 29239 29260
rect 29181 29251 29239 29257
rect 13170 29180 13176 29232
rect 13228 29220 13234 29232
rect 13449 29223 13507 29229
rect 13449 29220 13461 29223
rect 13228 29192 13461 29220
rect 13228 29180 13234 29192
rect 13449 29189 13461 29192
rect 13495 29220 13507 29223
rect 14458 29220 14464 29232
rect 13495 29192 14464 29220
rect 13495 29189 13507 29192
rect 13449 29183 13507 29189
rect 14458 29180 14464 29192
rect 14516 29180 14522 29232
rect 21634 29180 21640 29232
rect 21692 29220 21698 29232
rect 21821 29223 21879 29229
rect 21821 29220 21833 29223
rect 21692 29192 21833 29220
rect 21692 29180 21698 29192
rect 21821 29189 21833 29192
rect 21867 29189 21879 29223
rect 21821 29183 21879 29189
rect 25590 29180 25596 29232
rect 25648 29180 25654 29232
rect 31726 29220 31754 29260
rect 32306 29248 32312 29260
rect 32364 29248 32370 29300
rect 32398 29248 32404 29300
rect 32456 29288 32462 29300
rect 33137 29291 33195 29297
rect 33137 29288 33149 29291
rect 32456 29260 33149 29288
rect 32456 29248 32462 29260
rect 33137 29257 33149 29260
rect 33183 29257 33195 29291
rect 34882 29288 34888 29300
rect 33137 29251 33195 29257
rect 33336 29260 34888 29288
rect 32217 29223 32275 29229
rect 32217 29220 32229 29223
rect 31726 29192 32229 29220
rect 32217 29189 32229 29192
rect 32263 29189 32275 29223
rect 32217 29183 32275 29189
rect 9582 29152 9588 29164
rect 9543 29124 9588 29152
rect 9582 29112 9588 29124
rect 9640 29112 9646 29164
rect 13538 29112 13544 29164
rect 13596 29152 13602 29164
rect 14093 29155 14151 29161
rect 14093 29152 14105 29155
rect 13596 29124 14105 29152
rect 13596 29112 13602 29124
rect 14093 29121 14105 29124
rect 14139 29121 14151 29155
rect 14093 29115 14151 29121
rect 15194 29112 15200 29164
rect 15252 29152 15258 29164
rect 15381 29155 15439 29161
rect 15381 29152 15393 29155
rect 15252 29124 15393 29152
rect 15252 29112 15258 29124
rect 15381 29121 15393 29124
rect 15427 29152 15439 29155
rect 15654 29152 15660 29164
rect 15427 29124 15660 29152
rect 15427 29121 15439 29124
rect 15381 29115 15439 29121
rect 15654 29112 15660 29124
rect 15712 29112 15718 29164
rect 16850 29152 16856 29164
rect 16811 29124 16856 29152
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 22005 29155 22063 29161
rect 22005 29121 22017 29155
rect 22051 29152 22063 29155
rect 22462 29152 22468 29164
rect 22051 29124 22468 29152
rect 22051 29121 22063 29124
rect 22005 29115 22063 29121
rect 22462 29112 22468 29124
rect 22520 29152 22526 29164
rect 23290 29152 23296 29164
rect 22520 29124 23296 29152
rect 22520 29112 22526 29124
rect 23290 29112 23296 29124
rect 23348 29112 23354 29164
rect 24305 29155 24363 29161
rect 24305 29121 24317 29155
rect 24351 29121 24363 29155
rect 27890 29152 27896 29164
rect 27851 29124 27896 29152
rect 24305 29115 24363 29121
rect 15470 29084 15476 29096
rect 15431 29056 15476 29084
rect 15470 29044 15476 29056
rect 15528 29044 15534 29096
rect 15746 29084 15752 29096
rect 15707 29056 15752 29084
rect 15746 29044 15752 29056
rect 15804 29044 15810 29096
rect 13630 29016 13636 29028
rect 13591 28988 13636 29016
rect 13630 28976 13636 28988
rect 13688 28976 13694 29028
rect 14277 29019 14335 29025
rect 14277 28985 14289 29019
rect 14323 29016 14335 29019
rect 16868 29016 16896 29112
rect 24320 29084 24348 29115
rect 27890 29112 27896 29124
rect 27948 29112 27954 29164
rect 30650 29152 30656 29164
rect 30611 29124 30656 29152
rect 30650 29112 30656 29124
rect 30708 29112 30714 29164
rect 30837 29155 30895 29161
rect 30837 29121 30849 29155
rect 30883 29152 30895 29155
rect 31386 29152 31392 29164
rect 30883 29124 31392 29152
rect 30883 29121 30895 29124
rect 30837 29115 30895 29121
rect 31386 29112 31392 29124
rect 31444 29112 31450 29164
rect 33336 29161 33364 29260
rect 34882 29248 34888 29260
rect 34940 29288 34946 29300
rect 35989 29291 36047 29297
rect 35989 29288 36001 29291
rect 34940 29260 36001 29288
rect 34940 29248 34946 29260
rect 35989 29257 36001 29260
rect 36035 29257 36047 29291
rect 35989 29251 36047 29257
rect 34514 29220 34520 29232
rect 34475 29192 34520 29220
rect 34514 29180 34520 29192
rect 34572 29180 34578 29232
rect 35526 29180 35532 29232
rect 35584 29180 35590 29232
rect 33321 29155 33379 29161
rect 33321 29121 33333 29155
rect 33367 29121 33379 29155
rect 34238 29152 34244 29164
rect 34199 29124 34244 29152
rect 33321 29115 33379 29121
rect 34238 29112 34244 29124
rect 34296 29112 34302 29164
rect 24946 29084 24952 29096
rect 24320 29056 24952 29084
rect 24946 29044 24952 29056
rect 25004 29044 25010 29096
rect 30374 29044 30380 29096
rect 30432 29084 30438 29096
rect 33505 29087 33563 29093
rect 33505 29084 33517 29087
rect 30432 29056 30880 29084
rect 30432 29044 30438 29056
rect 21818 29016 21824 29028
rect 14323 28988 16896 29016
rect 21008 28988 21824 29016
rect 14323 28985 14335 28988
rect 14277 28979 14335 28985
rect 10134 28908 10140 28960
rect 10192 28948 10198 28960
rect 10686 28948 10692 28960
rect 10192 28920 10692 28948
rect 10192 28908 10198 28920
rect 10686 28908 10692 28920
rect 10744 28948 10750 28960
rect 12710 28948 12716 28960
rect 10744 28920 12716 28948
rect 10744 28908 10750 28920
rect 12710 28908 12716 28920
rect 12768 28908 12774 28960
rect 14734 28908 14740 28960
rect 14792 28948 14798 28960
rect 21008 28948 21036 28988
rect 21818 28976 21824 28988
rect 21876 28976 21882 29028
rect 26050 29016 26056 29028
rect 26011 28988 26056 29016
rect 26050 28976 26056 28988
rect 26108 28976 26114 29028
rect 27522 28976 27528 29028
rect 27580 29016 27586 29028
rect 30558 29016 30564 29028
rect 27580 28988 30564 29016
rect 27580 28976 27586 28988
rect 30558 28976 30564 28988
rect 30616 29016 30622 29028
rect 30742 29016 30748 29028
rect 30616 28988 30748 29016
rect 30616 28976 30622 28988
rect 14792 28920 21036 28948
rect 14792 28908 14798 28920
rect 21082 28908 21088 28960
rect 21140 28948 21146 28960
rect 22189 28951 22247 28957
rect 22189 28948 22201 28951
rect 21140 28920 22201 28948
rect 21140 28908 21146 28920
rect 22189 28917 22201 28920
rect 22235 28948 22247 28951
rect 22554 28948 22560 28960
rect 22235 28920 22560 28948
rect 22235 28917 22247 28920
rect 22189 28911 22247 28917
rect 22554 28908 22560 28920
rect 22612 28908 22618 28960
rect 24568 28951 24626 28957
rect 24568 28917 24580 28951
rect 24614 28948 24626 28951
rect 25314 28948 25320 28960
rect 24614 28920 25320 28948
rect 24614 28917 24626 28920
rect 24568 28911 24626 28917
rect 25314 28908 25320 28920
rect 25372 28908 25378 28960
rect 30668 28957 30696 28988
rect 30742 28976 30748 28988
rect 30800 28976 30806 29028
rect 30653 28951 30711 28957
rect 30653 28917 30665 28951
rect 30699 28917 30711 28951
rect 30852 28948 30880 29056
rect 31726 29056 33517 29084
rect 31018 29016 31024 29028
rect 30979 28988 31024 29016
rect 31018 28976 31024 28988
rect 31076 29016 31082 29028
rect 31726 29016 31754 29056
rect 33505 29053 33517 29056
rect 33551 29053 33563 29087
rect 33505 29047 33563 29053
rect 33597 29087 33655 29093
rect 33597 29053 33609 29087
rect 33643 29084 33655 29087
rect 34146 29084 34152 29096
rect 33643 29056 34152 29084
rect 33643 29053 33655 29056
rect 33597 29047 33655 29053
rect 34146 29044 34152 29056
rect 34204 29044 34210 29096
rect 31076 28988 31754 29016
rect 31076 28976 31082 28988
rect 33502 28948 33508 28960
rect 30852 28920 33508 28948
rect 30653 28911 30711 28917
rect 33502 28908 33508 28920
rect 33560 28908 33566 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 14458 28744 14464 28756
rect 14419 28716 14464 28744
rect 14458 28704 14464 28716
rect 14516 28704 14522 28756
rect 25869 28747 25927 28753
rect 14568 28716 22048 28744
rect 10594 28676 10600 28688
rect 10244 28648 10600 28676
rect 10244 28617 10272 28648
rect 10594 28636 10600 28648
rect 10652 28676 10658 28688
rect 10870 28676 10876 28688
rect 10652 28648 10876 28676
rect 10652 28636 10658 28648
rect 10870 28636 10876 28648
rect 10928 28636 10934 28688
rect 14090 28636 14096 28688
rect 14148 28676 14154 28688
rect 14568 28676 14596 28716
rect 14148 28648 14596 28676
rect 14148 28636 14154 28648
rect 10229 28611 10287 28617
rect 10229 28577 10241 28611
rect 10275 28577 10287 28611
rect 10229 28571 10287 28577
rect 10505 28611 10563 28617
rect 10505 28577 10517 28611
rect 10551 28608 10563 28611
rect 11241 28611 11299 28617
rect 11241 28608 11253 28611
rect 10551 28580 11253 28608
rect 10551 28577 10563 28580
rect 10505 28571 10563 28577
rect 11241 28577 11253 28580
rect 11287 28577 11299 28611
rect 11241 28571 11299 28577
rect 12710 28568 12716 28620
rect 12768 28608 12774 28620
rect 12989 28611 13047 28617
rect 12989 28608 13001 28611
rect 12768 28580 13001 28608
rect 12768 28568 12774 28580
rect 12989 28577 13001 28580
rect 13035 28577 13047 28611
rect 12989 28571 13047 28577
rect 14182 28568 14188 28620
rect 14240 28608 14246 28620
rect 16025 28611 16083 28617
rect 14240 28580 15332 28608
rect 14240 28568 14246 28580
rect 10134 28540 10140 28552
rect 10095 28512 10140 28540
rect 10134 28500 10140 28512
rect 10192 28500 10198 28552
rect 10962 28540 10968 28552
rect 10923 28512 10968 28540
rect 10962 28500 10968 28512
rect 11020 28500 11026 28552
rect 14093 28543 14151 28549
rect 14093 28509 14105 28543
rect 14139 28509 14151 28543
rect 14093 28503 14151 28509
rect 14277 28543 14335 28549
rect 14277 28509 14289 28543
rect 14323 28540 14335 28543
rect 14734 28540 14740 28552
rect 14323 28512 14740 28540
rect 14323 28509 14335 28512
rect 14277 28503 14335 28509
rect 11974 28432 11980 28484
rect 12032 28432 12038 28484
rect 14108 28472 14136 28503
rect 14734 28500 14740 28512
rect 14792 28500 14798 28552
rect 15105 28543 15163 28549
rect 15105 28509 15117 28543
rect 15151 28540 15163 28543
rect 15194 28540 15200 28552
rect 15151 28512 15200 28540
rect 15151 28509 15163 28512
rect 15105 28503 15163 28509
rect 15194 28500 15200 28512
rect 15252 28500 15258 28552
rect 15304 28549 15332 28580
rect 16025 28577 16037 28611
rect 16071 28608 16083 28611
rect 16666 28608 16672 28620
rect 16071 28580 16672 28608
rect 16071 28577 16083 28580
rect 16025 28571 16083 28577
rect 16666 28568 16672 28580
rect 16724 28568 16730 28620
rect 19521 28611 19579 28617
rect 19521 28577 19533 28611
rect 19567 28608 19579 28611
rect 21634 28608 21640 28620
rect 19567 28580 21640 28608
rect 19567 28577 19579 28580
rect 19521 28571 19579 28577
rect 21634 28568 21640 28580
rect 21692 28568 21698 28620
rect 22020 28608 22048 28716
rect 25869 28713 25881 28747
rect 25915 28744 25927 28747
rect 26234 28744 26240 28756
rect 25915 28716 26240 28744
rect 25915 28713 25927 28716
rect 25869 28707 25927 28713
rect 26234 28704 26240 28716
rect 26292 28704 26298 28756
rect 27798 28704 27804 28756
rect 27856 28744 27862 28756
rect 27985 28747 28043 28753
rect 27985 28744 27997 28747
rect 27856 28716 27997 28744
rect 27856 28704 27862 28716
rect 27985 28713 27997 28716
rect 28031 28713 28043 28747
rect 27985 28707 28043 28713
rect 28721 28747 28779 28753
rect 28721 28713 28733 28747
rect 28767 28744 28779 28747
rect 28810 28744 28816 28756
rect 28767 28716 28816 28744
rect 28767 28713 28779 28716
rect 28721 28707 28779 28713
rect 28810 28704 28816 28716
rect 28868 28704 28874 28756
rect 29822 28704 29828 28756
rect 29880 28744 29886 28756
rect 30101 28747 30159 28753
rect 30101 28744 30113 28747
rect 29880 28716 30113 28744
rect 29880 28704 29886 28716
rect 30101 28713 30113 28716
rect 30147 28713 30159 28747
rect 30101 28707 30159 28713
rect 30466 28704 30472 28756
rect 30524 28744 30530 28756
rect 30745 28747 30803 28753
rect 30745 28744 30757 28747
rect 30524 28716 30757 28744
rect 30524 28704 30530 28716
rect 30745 28713 30757 28716
rect 30791 28713 30803 28747
rect 30745 28707 30803 28713
rect 31478 28704 31484 28756
rect 31536 28744 31542 28756
rect 32309 28747 32367 28753
rect 32309 28744 32321 28747
rect 31536 28716 32321 28744
rect 31536 28704 31542 28716
rect 32309 28713 32321 28716
rect 32355 28713 32367 28747
rect 33502 28744 33508 28756
rect 33463 28716 33508 28744
rect 32309 28707 32367 28713
rect 33502 28704 33508 28716
rect 33560 28744 33566 28756
rect 33962 28744 33968 28756
rect 33560 28716 33968 28744
rect 33560 28704 33566 28716
rect 33962 28704 33968 28716
rect 34020 28704 34026 28756
rect 34885 28747 34943 28753
rect 34885 28713 34897 28747
rect 34931 28744 34943 28747
rect 35342 28744 35348 28756
rect 34931 28716 35348 28744
rect 34931 28713 34943 28716
rect 34885 28707 34943 28713
rect 35342 28704 35348 28716
rect 35400 28704 35406 28756
rect 35526 28744 35532 28756
rect 35487 28716 35532 28744
rect 35526 28704 35532 28716
rect 35584 28704 35590 28756
rect 22738 28636 22744 28688
rect 22796 28676 22802 28688
rect 22922 28676 22928 28688
rect 22796 28648 22928 28676
rect 22796 28636 22802 28648
rect 22922 28636 22928 28648
rect 22980 28676 22986 28688
rect 22980 28648 27660 28676
rect 22980 28636 22986 28648
rect 24765 28611 24823 28617
rect 24765 28608 24777 28611
rect 22020 28580 24777 28608
rect 24765 28577 24777 28580
rect 24811 28577 24823 28611
rect 26050 28608 26056 28620
rect 24765 28571 24823 28577
rect 24872 28580 26056 28608
rect 15289 28543 15347 28549
rect 15289 28509 15301 28543
rect 15335 28509 15347 28543
rect 15289 28503 15347 28509
rect 15473 28543 15531 28549
rect 15473 28509 15485 28543
rect 15519 28540 15531 28543
rect 15930 28540 15936 28552
rect 15519 28512 15936 28540
rect 15519 28509 15531 28512
rect 15473 28503 15531 28509
rect 15930 28500 15936 28512
rect 15988 28500 15994 28552
rect 17770 28500 17776 28552
rect 17828 28540 17834 28552
rect 18233 28543 18291 28549
rect 18233 28540 18245 28543
rect 17828 28512 18245 28540
rect 17828 28500 17834 28512
rect 18233 28509 18245 28512
rect 18279 28509 18291 28543
rect 18233 28503 18291 28509
rect 19245 28543 19303 28549
rect 19245 28509 19257 28543
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 14550 28472 14556 28484
rect 14108 28444 14556 28472
rect 14550 28432 14556 28444
rect 14608 28432 14614 28484
rect 14921 28475 14979 28481
rect 14921 28441 14933 28475
rect 14967 28472 14979 28475
rect 15562 28472 15568 28484
rect 14967 28444 15568 28472
rect 14967 28441 14979 28444
rect 14921 28435 14979 28441
rect 15562 28432 15568 28444
rect 15620 28432 15626 28484
rect 16298 28472 16304 28484
rect 16259 28444 16304 28472
rect 16298 28432 16304 28444
rect 16356 28432 16362 28484
rect 17310 28432 17316 28484
rect 17368 28432 17374 28484
rect 19260 28472 19288 28503
rect 20990 28500 20996 28552
rect 21048 28540 21054 28552
rect 21453 28543 21511 28549
rect 21453 28540 21465 28543
rect 21048 28512 21465 28540
rect 21048 28500 21054 28512
rect 21453 28509 21465 28512
rect 21499 28509 21511 28543
rect 21453 28503 21511 28509
rect 21818 28500 21824 28552
rect 21876 28540 21882 28552
rect 22649 28543 22707 28549
rect 21876 28512 21921 28540
rect 21876 28500 21882 28512
rect 22649 28509 22661 28543
rect 22695 28540 22707 28543
rect 22738 28540 22744 28552
rect 22695 28512 22744 28540
rect 22695 28509 22707 28512
rect 22649 28503 22707 28509
rect 22738 28500 22744 28512
rect 22796 28500 22802 28552
rect 22925 28543 22983 28549
rect 22925 28509 22937 28543
rect 22971 28509 22983 28543
rect 22925 28503 22983 28509
rect 24397 28543 24455 28549
rect 24397 28509 24409 28543
rect 24443 28509 24455 28543
rect 24578 28540 24584 28552
rect 24539 28512 24584 28540
rect 24397 28503 24455 28509
rect 19426 28472 19432 28484
rect 19260 28444 19432 28472
rect 19426 28432 19432 28444
rect 19484 28432 19490 28484
rect 20530 28432 20536 28484
rect 20588 28432 20594 28484
rect 21174 28432 21180 28484
rect 21232 28472 21238 28484
rect 21637 28475 21695 28481
rect 21637 28472 21649 28475
rect 21232 28444 21649 28472
rect 21232 28432 21238 28444
rect 21637 28441 21649 28444
rect 21683 28441 21695 28475
rect 21637 28435 21695 28441
rect 21726 28432 21732 28484
rect 21784 28472 21790 28484
rect 21784 28444 21829 28472
rect 21784 28432 21790 28444
rect 22554 28432 22560 28484
rect 22612 28472 22618 28484
rect 22940 28472 22968 28503
rect 22612 28444 22968 28472
rect 24412 28472 24440 28503
rect 24578 28500 24584 28512
rect 24636 28500 24642 28552
rect 24673 28543 24731 28549
rect 24673 28509 24685 28543
rect 24719 28540 24731 28543
rect 24872 28540 24900 28580
rect 26050 28568 26056 28580
rect 26108 28568 26114 28620
rect 24719 28512 24900 28540
rect 24949 28543 25007 28549
rect 24719 28509 24731 28512
rect 24673 28503 24731 28509
rect 24949 28509 24961 28543
rect 24995 28509 25007 28543
rect 24949 28503 25007 28509
rect 25685 28543 25743 28549
rect 25685 28509 25697 28543
rect 25731 28509 25743 28543
rect 25685 28503 25743 28509
rect 24762 28472 24768 28484
rect 24412 28444 24768 28472
rect 22612 28432 22618 28444
rect 24762 28432 24768 28444
rect 24820 28432 24826 28484
rect 24964 28472 24992 28503
rect 24872 28444 24992 28472
rect 25133 28475 25191 28481
rect 14366 28364 14372 28416
rect 14424 28404 14430 28416
rect 15197 28407 15255 28413
rect 15197 28404 15209 28407
rect 14424 28376 15209 28404
rect 14424 28364 14430 28376
rect 15197 28373 15209 28376
rect 15243 28373 15255 28407
rect 15580 28404 15608 28432
rect 17773 28407 17831 28413
rect 17773 28404 17785 28407
rect 15580 28376 17785 28404
rect 15197 28367 15255 28373
rect 17773 28373 17785 28376
rect 17819 28404 17831 28407
rect 18046 28404 18052 28416
rect 17819 28376 18052 28404
rect 17819 28373 17831 28376
rect 17773 28367 17831 28373
rect 18046 28364 18052 28376
rect 18104 28364 18110 28416
rect 18230 28364 18236 28416
rect 18288 28404 18294 28416
rect 18325 28407 18383 28413
rect 18325 28404 18337 28407
rect 18288 28376 18337 28404
rect 18288 28364 18294 28376
rect 18325 28373 18337 28376
rect 18371 28373 18383 28407
rect 18325 28367 18383 28373
rect 20993 28407 21051 28413
rect 20993 28373 21005 28407
rect 21039 28404 21051 28407
rect 21358 28404 21364 28416
rect 21039 28376 21364 28404
rect 21039 28373 21051 28376
rect 20993 28367 21051 28373
rect 21358 28364 21364 28376
rect 21416 28364 21422 28416
rect 22002 28404 22008 28416
rect 21963 28376 22008 28404
rect 22002 28364 22008 28376
rect 22060 28364 22066 28416
rect 22278 28364 22284 28416
rect 22336 28404 22342 28416
rect 22465 28407 22523 28413
rect 22465 28404 22477 28407
rect 22336 28376 22477 28404
rect 22336 28364 22342 28376
rect 22465 28373 22477 28376
rect 22511 28373 22523 28407
rect 22465 28367 22523 28373
rect 22833 28407 22891 28413
rect 22833 28373 22845 28407
rect 22879 28404 22891 28407
rect 24872 28404 24900 28444
rect 25133 28441 25145 28475
rect 25179 28472 25191 28475
rect 25314 28472 25320 28484
rect 25179 28444 25320 28472
rect 25179 28441 25191 28444
rect 25133 28435 25191 28441
rect 25314 28432 25320 28444
rect 25372 28432 25378 28484
rect 25406 28432 25412 28484
rect 25464 28472 25470 28484
rect 25700 28472 25728 28503
rect 26326 28500 26332 28552
rect 26384 28540 26390 28552
rect 27522 28549 27528 28552
rect 27341 28543 27399 28549
rect 27341 28540 27353 28543
rect 26384 28512 27353 28540
rect 26384 28500 26390 28512
rect 27341 28509 27353 28512
rect 27387 28509 27399 28543
rect 27341 28503 27399 28509
rect 27489 28543 27528 28549
rect 27489 28509 27501 28543
rect 27489 28503 27528 28509
rect 27522 28500 27528 28503
rect 27580 28500 27586 28552
rect 26970 28472 26976 28484
rect 25464 28444 26976 28472
rect 25464 28432 25470 28444
rect 26970 28432 26976 28444
rect 27028 28432 27034 28484
rect 27632 28481 27660 28648
rect 27706 28636 27712 28688
rect 27764 28636 27770 28688
rect 28166 28636 28172 28688
rect 28224 28676 28230 28688
rect 28905 28679 28963 28685
rect 28905 28676 28917 28679
rect 28224 28648 28917 28676
rect 28224 28636 28230 28648
rect 28905 28645 28917 28648
rect 28951 28676 28963 28679
rect 30650 28676 30656 28688
rect 28951 28648 30656 28676
rect 28951 28645 28963 28648
rect 28905 28639 28963 28645
rect 30650 28636 30656 28648
rect 30708 28636 30714 28688
rect 27724 28549 27752 28636
rect 27982 28568 27988 28620
rect 28040 28608 28046 28620
rect 28626 28608 28632 28620
rect 28040 28580 28396 28608
rect 28587 28580 28632 28608
rect 28040 28568 28046 28580
rect 27709 28543 27767 28549
rect 27709 28509 27721 28543
rect 27755 28509 27767 28543
rect 27709 28503 27767 28509
rect 27798 28500 27804 28552
rect 27856 28549 27862 28552
rect 27856 28540 27864 28549
rect 28166 28540 28172 28552
rect 27856 28512 27901 28540
rect 28000 28512 28172 28540
rect 27856 28503 27864 28512
rect 27856 28500 27862 28503
rect 27617 28475 27675 28481
rect 27617 28441 27629 28475
rect 27663 28472 27675 28475
rect 28000 28472 28028 28512
rect 28166 28500 28172 28512
rect 28224 28500 28230 28552
rect 27663 28444 28028 28472
rect 28368 28472 28396 28580
rect 28626 28568 28632 28580
rect 28684 28568 28690 28620
rect 30837 28611 30895 28617
rect 30837 28608 30849 28611
rect 29932 28580 30849 28608
rect 28534 28540 28540 28552
rect 28495 28512 28540 28540
rect 28534 28500 28540 28512
rect 28592 28500 28598 28552
rect 28718 28500 28724 28552
rect 28776 28540 28782 28552
rect 29932 28549 29960 28580
rect 30837 28577 30849 28580
rect 30883 28608 30895 28611
rect 31386 28608 31392 28620
rect 30883 28580 31392 28608
rect 30883 28577 30895 28580
rect 30837 28571 30895 28577
rect 31386 28568 31392 28580
rect 31444 28568 31450 28620
rect 31588 28580 32536 28608
rect 31588 28552 31616 28580
rect 29917 28543 29975 28549
rect 28776 28512 29868 28540
rect 28776 28500 28782 28512
rect 29733 28475 29791 28481
rect 29733 28472 29745 28475
rect 28368 28444 29745 28472
rect 27663 28441 27675 28444
rect 27617 28435 27675 28441
rect 29733 28441 29745 28444
rect 29779 28441 29791 28475
rect 29840 28472 29868 28512
rect 29917 28509 29929 28543
rect 29963 28509 29975 28543
rect 30558 28540 30564 28552
rect 30519 28512 30564 28540
rect 29917 28503 29975 28509
rect 30558 28500 30564 28512
rect 30616 28500 30622 28552
rect 31570 28540 31576 28552
rect 31531 28512 31576 28540
rect 31570 28500 31576 28512
rect 31628 28500 31634 28552
rect 31665 28543 31723 28549
rect 31665 28509 31677 28543
rect 31711 28540 31723 28543
rect 32030 28540 32036 28552
rect 31711 28512 32036 28540
rect 31711 28509 31723 28512
rect 31665 28503 31723 28509
rect 32030 28500 32036 28512
rect 32088 28540 32094 28552
rect 32508 28549 32536 28580
rect 32309 28543 32367 28549
rect 32309 28540 32321 28543
rect 32088 28512 32321 28540
rect 32088 28500 32094 28512
rect 32309 28509 32321 28512
rect 32355 28509 32367 28543
rect 32309 28503 32367 28509
rect 32493 28543 32551 28549
rect 32493 28509 32505 28543
rect 32539 28540 32551 28543
rect 34606 28540 34612 28552
rect 32539 28512 34612 28540
rect 32539 28509 32551 28512
rect 32493 28503 32551 28509
rect 34606 28500 34612 28512
rect 34664 28500 34670 28552
rect 34701 28543 34759 28549
rect 34701 28509 34713 28543
rect 34747 28509 34759 28543
rect 34701 28503 34759 28509
rect 33410 28472 33416 28484
rect 29840 28444 33416 28472
rect 29733 28435 29791 28441
rect 33410 28432 33416 28444
rect 33468 28432 33474 28484
rect 33502 28432 33508 28484
rect 33560 28472 33566 28484
rect 34716 28472 34744 28503
rect 35342 28500 35348 28552
rect 35400 28540 35406 28552
rect 35437 28543 35495 28549
rect 35437 28540 35449 28543
rect 35400 28512 35449 28540
rect 35400 28500 35406 28512
rect 35437 28509 35449 28512
rect 35483 28509 35495 28543
rect 35437 28503 35495 28509
rect 46934 28500 46940 28552
rect 46992 28540 46998 28552
rect 47673 28543 47731 28549
rect 47673 28540 47685 28543
rect 46992 28512 47685 28540
rect 46992 28500 46998 28512
rect 47673 28509 47685 28512
rect 47719 28509 47731 28543
rect 47673 28503 47731 28509
rect 33560 28444 34744 28472
rect 33560 28432 33566 28444
rect 30374 28404 30380 28416
rect 22879 28376 30380 28404
rect 22879 28373 22891 28376
rect 22833 28367 22891 28373
rect 30374 28364 30380 28376
rect 30432 28364 30438 28416
rect 31386 28364 31392 28416
rect 31444 28404 31450 28416
rect 31849 28407 31907 28413
rect 31849 28404 31861 28407
rect 31444 28376 31861 28404
rect 31444 28364 31450 28376
rect 31849 28373 31861 28376
rect 31895 28373 31907 28407
rect 31849 28367 31907 28373
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 1762 28160 1768 28212
rect 1820 28200 1826 28212
rect 14090 28200 14096 28212
rect 1820 28172 14096 28200
rect 1820 28160 1826 28172
rect 14090 28160 14096 28172
rect 14148 28160 14154 28212
rect 14182 28160 14188 28212
rect 14240 28200 14246 28212
rect 14645 28203 14703 28209
rect 14645 28200 14657 28203
rect 14240 28172 14657 28200
rect 14240 28160 14246 28172
rect 14645 28169 14657 28172
rect 14691 28169 14703 28203
rect 14645 28163 14703 28169
rect 16298 28160 16304 28212
rect 16356 28200 16362 28212
rect 16945 28203 17003 28209
rect 16945 28200 16957 28203
rect 16356 28172 16957 28200
rect 16356 28160 16362 28172
rect 16945 28169 16957 28172
rect 16991 28169 17003 28203
rect 20530 28200 20536 28212
rect 20491 28172 20536 28200
rect 16945 28163 17003 28169
rect 20530 28160 20536 28172
rect 20588 28160 20594 28212
rect 21174 28200 21180 28212
rect 21135 28172 21180 28200
rect 21174 28160 21180 28172
rect 21232 28160 21238 28212
rect 21358 28160 21364 28212
rect 21416 28200 21422 28212
rect 22189 28203 22247 28209
rect 22189 28200 22201 28203
rect 21416 28172 22201 28200
rect 21416 28160 21422 28172
rect 22189 28169 22201 28172
rect 22235 28200 22247 28203
rect 22370 28200 22376 28212
rect 22235 28172 22376 28200
rect 22235 28169 22247 28172
rect 22189 28163 22247 28169
rect 22370 28160 22376 28172
rect 22428 28160 22434 28212
rect 24857 28203 24915 28209
rect 24857 28169 24869 28203
rect 24903 28200 24915 28203
rect 25406 28200 25412 28212
rect 24903 28172 25412 28200
rect 24903 28169 24915 28172
rect 24857 28163 24915 28169
rect 25406 28160 25412 28172
rect 25464 28160 25470 28212
rect 25590 28200 25596 28212
rect 25551 28172 25596 28200
rect 25590 28160 25596 28172
rect 25648 28160 25654 28212
rect 26326 28200 26332 28212
rect 26287 28172 26332 28200
rect 26326 28160 26332 28172
rect 26384 28160 26390 28212
rect 27154 28200 27160 28212
rect 27115 28172 27160 28200
rect 27154 28160 27160 28172
rect 27212 28160 27218 28212
rect 27430 28160 27436 28212
rect 27488 28200 27494 28212
rect 27893 28203 27951 28209
rect 27893 28200 27905 28203
rect 27488 28172 27905 28200
rect 27488 28160 27494 28172
rect 27893 28169 27905 28172
rect 27939 28200 27951 28203
rect 28718 28200 28724 28212
rect 27939 28172 28724 28200
rect 27939 28169 27951 28172
rect 27893 28163 27951 28169
rect 28718 28160 28724 28172
rect 28776 28160 28782 28212
rect 29288 28172 41414 28200
rect 9140 28104 10916 28132
rect 9140 28073 9168 28104
rect 9125 28067 9183 28073
rect 9125 28033 9137 28067
rect 9171 28033 9183 28067
rect 10888 28064 10916 28104
rect 10962 28092 10968 28144
rect 11020 28132 11026 28144
rect 11793 28135 11851 28141
rect 11793 28132 11805 28135
rect 11020 28104 11805 28132
rect 11020 28092 11026 28104
rect 11793 28101 11805 28104
rect 11839 28101 11851 28135
rect 11793 28095 11851 28101
rect 14921 28135 14979 28141
rect 14921 28101 14933 28135
rect 14967 28132 14979 28135
rect 15470 28132 15476 28144
rect 14967 28104 15476 28132
rect 14967 28101 14979 28104
rect 14921 28095 14979 28101
rect 15470 28092 15476 28104
rect 15528 28132 15534 28144
rect 15528 28104 15884 28132
rect 15528 28092 15534 28104
rect 11330 28064 11336 28076
rect 10888 28036 11336 28064
rect 9125 28027 9183 28033
rect 11330 28024 11336 28036
rect 11388 28024 11394 28076
rect 11517 28067 11575 28073
rect 11517 28033 11529 28067
rect 11563 28033 11575 28067
rect 11517 28027 11575 28033
rect 13541 28067 13599 28073
rect 13541 28033 13553 28067
rect 13587 28033 13599 28067
rect 14550 28064 14556 28076
rect 14511 28036 14556 28064
rect 13541 28027 13599 28033
rect 9309 27999 9367 28005
rect 9309 27965 9321 27999
rect 9355 27996 9367 27999
rect 9674 27996 9680 28008
rect 9355 27968 9680 27996
rect 9355 27965 9367 27968
rect 9309 27959 9367 27965
rect 9674 27956 9680 27968
rect 9732 27956 9738 28008
rect 9769 27999 9827 28005
rect 9769 27965 9781 27999
rect 9815 27965 9827 27999
rect 9769 27959 9827 27965
rect 7558 27888 7564 27940
rect 7616 27928 7622 27940
rect 9784 27928 9812 27959
rect 10778 27956 10784 28008
rect 10836 27996 10842 28008
rect 11532 27996 11560 28027
rect 10836 27968 11560 27996
rect 13556 27996 13584 28027
rect 14550 28024 14556 28036
rect 14608 28024 14614 28076
rect 14734 28024 14740 28076
rect 14792 28064 14798 28076
rect 15562 28064 15568 28076
rect 14792 28036 14837 28064
rect 15523 28036 15568 28064
rect 14792 28024 14798 28036
rect 15562 28024 15568 28036
rect 15620 28024 15626 28076
rect 15746 28064 15752 28076
rect 15707 28036 15752 28064
rect 15746 28024 15752 28036
rect 15804 28024 15810 28076
rect 15856 28073 15884 28104
rect 15930 28092 15936 28144
rect 15988 28132 15994 28144
rect 17037 28135 17095 28141
rect 17037 28132 17049 28135
rect 15988 28104 17049 28132
rect 15988 28092 15994 28104
rect 17037 28101 17049 28104
rect 17083 28101 17095 28135
rect 18230 28132 18236 28144
rect 18191 28104 18236 28132
rect 17037 28095 17095 28101
rect 18230 28092 18236 28104
rect 18288 28092 18294 28144
rect 21634 28092 21640 28144
rect 21692 28132 21698 28144
rect 21821 28135 21879 28141
rect 21821 28132 21833 28135
rect 21692 28104 21833 28132
rect 21692 28092 21698 28104
rect 21821 28101 21833 28104
rect 21867 28101 21879 28135
rect 27614 28132 27620 28144
rect 21821 28095 21879 28101
rect 21928 28104 22968 28132
rect 15841 28067 15899 28073
rect 15841 28033 15853 28067
rect 15887 28033 15899 28067
rect 15841 28027 15899 28033
rect 16482 28024 16488 28076
rect 16540 28064 16546 28076
rect 17129 28067 17187 28073
rect 17129 28064 17141 28067
rect 16540 28036 17141 28064
rect 16540 28024 16546 28036
rect 17129 28033 17141 28036
rect 17175 28033 17187 28067
rect 18046 28064 18052 28076
rect 18007 28036 18052 28064
rect 17129 28027 17187 28033
rect 18046 28024 18052 28036
rect 18104 28024 18110 28076
rect 20254 28064 20260 28076
rect 19812 28036 20260 28064
rect 15381 27999 15439 28005
rect 13556 27968 15332 27996
rect 10836 27956 10842 27968
rect 14366 27928 14372 27940
rect 7616 27900 9812 27928
rect 14327 27900 14372 27928
rect 7616 27888 7622 27900
rect 14366 27888 14372 27900
rect 14424 27888 14430 27940
rect 15304 27928 15332 27968
rect 15381 27965 15393 27999
rect 15427 27996 15439 27999
rect 16669 27999 16727 28005
rect 16669 27996 16681 27999
rect 15427 27968 16681 27996
rect 15427 27965 15439 27968
rect 15381 27959 15439 27965
rect 16669 27965 16681 27968
rect 16715 27965 16727 27999
rect 16669 27959 16727 27965
rect 19812 27928 19840 28036
rect 20254 28024 20260 28036
rect 20312 28064 20318 28076
rect 20441 28067 20499 28073
rect 20312 28036 20392 28064
rect 20312 28024 20318 28036
rect 19889 27999 19947 28005
rect 19889 27965 19901 27999
rect 19935 27965 19947 27999
rect 20364 27996 20392 28036
rect 20441 28033 20453 28067
rect 20487 28064 20499 28067
rect 20622 28064 20628 28076
rect 20487 28036 20628 28064
rect 20487 28033 20499 28036
rect 20441 28027 20499 28033
rect 20622 28024 20628 28036
rect 20680 28024 20686 28076
rect 21082 28064 21088 28076
rect 21043 28036 21088 28064
rect 21082 28024 21088 28036
rect 21140 28024 21146 28076
rect 21269 28067 21327 28073
rect 21269 28033 21281 28067
rect 21315 28064 21327 28067
rect 21358 28064 21364 28076
rect 21315 28036 21364 28064
rect 21315 28033 21327 28036
rect 21269 28027 21327 28033
rect 21358 28024 21364 28036
rect 21416 28024 21422 28076
rect 21928 27996 21956 28104
rect 22002 28024 22008 28076
rect 22060 28073 22066 28076
rect 22060 28067 22109 28073
rect 22060 28033 22063 28067
rect 22097 28033 22109 28067
rect 22060 28027 22109 28033
rect 22060 28024 22066 28027
rect 22278 28024 22284 28076
rect 22336 28064 22342 28076
rect 22940 28073 22968 28104
rect 26252 28104 27620 28132
rect 26252 28073 26280 28104
rect 27614 28092 27620 28104
rect 27672 28092 27678 28144
rect 27798 28132 27804 28144
rect 27724 28104 27804 28132
rect 22925 28067 22983 28073
rect 22336 28036 22381 28064
rect 22336 28024 22342 28036
rect 22925 28033 22937 28067
rect 22971 28064 22983 28067
rect 24673 28067 24731 28073
rect 24673 28064 24685 28067
rect 22971 28036 24685 28064
rect 22971 28033 22983 28036
rect 22925 28027 22983 28033
rect 24673 28033 24685 28036
rect 24719 28033 24731 28067
rect 24673 28027 24731 28033
rect 25501 28067 25559 28073
rect 25501 28033 25513 28067
rect 25547 28033 25559 28067
rect 25501 28027 25559 28033
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28033 26295 28067
rect 26418 28064 26424 28076
rect 26379 28036 26424 28064
rect 26237 28027 26295 28033
rect 20364 27968 21956 27996
rect 25516 27996 25544 28027
rect 26418 28024 26424 28036
rect 26476 28024 26482 28076
rect 27065 28067 27123 28073
rect 27065 28033 27077 28067
rect 27111 28064 27123 28067
rect 27430 28064 27436 28076
rect 27111 28036 27436 28064
rect 27111 28033 27123 28036
rect 27065 28027 27123 28033
rect 27430 28024 27436 28036
rect 27488 28024 27494 28076
rect 27724 28073 27752 28104
rect 27798 28092 27804 28104
rect 27856 28132 27862 28144
rect 29181 28135 29239 28141
rect 29181 28132 29193 28135
rect 27856 28104 29193 28132
rect 27856 28092 27862 28104
rect 29181 28101 29193 28104
rect 29227 28101 29239 28135
rect 29181 28095 29239 28101
rect 27709 28067 27767 28073
rect 27709 28033 27721 28067
rect 27755 28033 27767 28067
rect 27709 28027 27767 28033
rect 28074 28024 28080 28076
rect 28132 28064 28138 28076
rect 28445 28067 28503 28073
rect 28445 28064 28457 28067
rect 28132 28036 28457 28064
rect 28132 28024 28138 28036
rect 28445 28033 28457 28036
rect 28491 28033 28503 28067
rect 29086 28064 29092 28076
rect 29047 28036 29092 28064
rect 28445 28027 28503 28033
rect 29086 28024 29092 28036
rect 29144 28024 29150 28076
rect 26326 27996 26332 28008
rect 25516 27968 26332 27996
rect 19889 27959 19947 27965
rect 15304 27900 19840 27928
rect 19904 27928 19932 27959
rect 26326 27956 26332 27968
rect 26384 27956 26390 28008
rect 27154 27956 27160 28008
rect 27212 27996 27218 28008
rect 28537 27999 28595 28005
rect 28537 27996 28549 27999
rect 27212 27968 28549 27996
rect 27212 27956 27218 27968
rect 28537 27965 28549 27968
rect 28583 27965 28595 27999
rect 28537 27959 28595 27965
rect 29288 27928 29316 28172
rect 30377 28135 30435 28141
rect 30377 28101 30389 28135
rect 30423 28132 30435 28135
rect 32306 28132 32312 28144
rect 30423 28104 32312 28132
rect 30423 28101 30435 28104
rect 30377 28095 30435 28101
rect 32306 28092 32312 28104
rect 32364 28092 32370 28144
rect 35253 28135 35311 28141
rect 35253 28132 35265 28135
rect 34454 28104 35265 28132
rect 35253 28101 35265 28104
rect 35299 28101 35311 28135
rect 35253 28095 35311 28101
rect 31202 28064 31208 28076
rect 31163 28036 31208 28064
rect 31202 28024 31208 28036
rect 31260 28024 31266 28076
rect 31386 28064 31392 28076
rect 31347 28036 31392 28064
rect 31386 28024 31392 28036
rect 31444 28024 31450 28076
rect 31478 28024 31484 28076
rect 31536 28064 31542 28076
rect 35161 28067 35219 28073
rect 31536 28036 31581 28064
rect 31536 28024 31542 28036
rect 35161 28033 35173 28067
rect 35207 28064 35219 28067
rect 35342 28064 35348 28076
rect 35207 28036 35348 28064
rect 35207 28033 35219 28036
rect 35161 28027 35219 28033
rect 35342 28024 35348 28036
rect 35400 28024 35406 28076
rect 32953 27999 33011 28005
rect 32953 27996 32965 27999
rect 31726 27968 32965 27996
rect 19904 27900 21956 27928
rect 13538 27820 13544 27872
rect 13596 27860 13602 27872
rect 13633 27863 13691 27869
rect 13633 27860 13645 27863
rect 13596 27832 13645 27860
rect 13596 27820 13602 27832
rect 13633 27829 13645 27832
rect 13679 27829 13691 27863
rect 21928 27860 21956 27900
rect 23032 27900 29316 27928
rect 30561 27931 30619 27937
rect 23032 27860 23060 27900
rect 30561 27897 30573 27931
rect 30607 27928 30619 27931
rect 31478 27928 31484 27940
rect 30607 27900 31484 27928
rect 30607 27897 30619 27900
rect 30561 27891 30619 27897
rect 31478 27888 31484 27900
rect 31536 27928 31542 27940
rect 31726 27928 31754 27968
rect 32953 27965 32965 27968
rect 32999 27965 33011 27999
rect 33226 27996 33232 28008
rect 33187 27968 33232 27996
rect 32953 27959 33011 27965
rect 33226 27956 33232 27968
rect 33284 27956 33290 28008
rect 34698 27996 34704 28008
rect 34659 27968 34704 27996
rect 34698 27956 34704 27968
rect 34756 27956 34762 28008
rect 41386 27996 41414 28172
rect 47578 28064 47584 28076
rect 47539 28036 47584 28064
rect 47578 28024 47584 28036
rect 47636 28024 47642 28076
rect 46382 27996 46388 28008
rect 41386 27968 46388 27996
rect 46382 27956 46388 27968
rect 46440 27956 46446 28008
rect 31536 27900 31754 27928
rect 31536 27888 31542 27900
rect 21928 27832 23060 27860
rect 13633 27823 13691 27829
rect 23106 27820 23112 27872
rect 23164 27860 23170 27872
rect 23164 27832 23209 27860
rect 23164 27820 23170 27832
rect 25682 27820 25688 27872
rect 25740 27860 25746 27872
rect 27062 27860 27068 27872
rect 25740 27832 27068 27860
rect 25740 27820 25746 27832
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 28166 27820 28172 27872
rect 28224 27860 28230 27872
rect 30742 27860 30748 27872
rect 28224 27832 30748 27860
rect 28224 27820 28230 27832
rect 30742 27820 30748 27832
rect 30800 27820 30806 27872
rect 31018 27860 31024 27872
rect 30979 27832 31024 27860
rect 31018 27820 31024 27832
rect 31076 27820 31082 27872
rect 47670 27860 47676 27872
rect 47631 27832 47676 27860
rect 47670 27820 47676 27832
rect 47728 27820 47734 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 3970 27616 3976 27668
rect 4028 27656 4034 27668
rect 21174 27656 21180 27668
rect 4028 27628 14596 27656
rect 4028 27616 4034 27628
rect 9674 27588 9680 27600
rect 9635 27560 9680 27588
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 11974 27548 11980 27600
rect 12032 27588 12038 27600
rect 12069 27591 12127 27597
rect 12069 27588 12081 27591
rect 12032 27560 12081 27588
rect 12032 27548 12038 27560
rect 12069 27557 12081 27560
rect 12115 27557 12127 27591
rect 12069 27551 12127 27557
rect 14568 27529 14596 27628
rect 20732 27628 21180 27656
rect 15746 27548 15752 27600
rect 15804 27588 15810 27600
rect 17862 27588 17868 27600
rect 15804 27560 17868 27588
rect 15804 27548 15810 27560
rect 17862 27548 17868 27560
rect 17920 27548 17926 27600
rect 20533 27591 20591 27597
rect 20533 27557 20545 27591
rect 20579 27588 20591 27591
rect 20732 27588 20760 27628
rect 21174 27616 21180 27628
rect 21232 27616 21238 27668
rect 21542 27656 21548 27668
rect 21503 27628 21548 27656
rect 21542 27616 21548 27628
rect 21600 27656 21606 27668
rect 23201 27659 23259 27665
rect 23201 27656 23213 27659
rect 21600 27628 23213 27656
rect 21600 27616 21606 27628
rect 23201 27625 23213 27628
rect 23247 27625 23259 27659
rect 23201 27619 23259 27625
rect 26418 27616 26424 27668
rect 26476 27656 26482 27668
rect 28442 27656 28448 27668
rect 26476 27628 28448 27656
rect 26476 27616 26482 27628
rect 28442 27616 28448 27628
rect 28500 27616 28506 27668
rect 28534 27616 28540 27668
rect 28592 27656 28598 27668
rect 33502 27656 33508 27668
rect 28592 27628 33508 27656
rect 28592 27616 28598 27628
rect 33502 27616 33508 27628
rect 33560 27656 33566 27668
rect 33870 27656 33876 27668
rect 33560 27628 33876 27656
rect 33560 27616 33566 27628
rect 33870 27616 33876 27628
rect 33928 27616 33934 27668
rect 23569 27591 23627 27597
rect 23569 27588 23581 27591
rect 20579 27560 20760 27588
rect 20824 27560 23581 27588
rect 20579 27557 20591 27560
rect 20533 27551 20591 27557
rect 14553 27523 14611 27529
rect 14553 27489 14565 27523
rect 14599 27489 14611 27523
rect 16666 27520 16672 27532
rect 16627 27492 16672 27520
rect 14553 27483 14611 27489
rect 16666 27480 16672 27492
rect 16724 27480 16730 27532
rect 20824 27529 20852 27560
rect 23569 27557 23581 27560
rect 23615 27588 23627 27591
rect 24210 27588 24216 27600
rect 23615 27560 24216 27588
rect 23615 27557 23627 27560
rect 23569 27551 23627 27557
rect 24210 27548 24216 27560
rect 24268 27548 24274 27600
rect 27065 27591 27123 27597
rect 27065 27557 27077 27591
rect 27111 27588 27123 27591
rect 27246 27588 27252 27600
rect 27111 27560 27252 27588
rect 27111 27557 27123 27560
rect 27065 27551 27123 27557
rect 27246 27548 27252 27560
rect 27304 27548 27310 27600
rect 29086 27588 29092 27600
rect 27540 27560 29092 27588
rect 20809 27523 20867 27529
rect 20809 27489 20821 27523
rect 20855 27489 20867 27523
rect 20809 27483 20867 27489
rect 20990 27480 20996 27532
rect 21048 27520 21054 27532
rect 21453 27523 21511 27529
rect 21453 27520 21465 27523
rect 21048 27492 21465 27520
rect 21048 27480 21054 27492
rect 21453 27489 21465 27492
rect 21499 27520 21511 27523
rect 22741 27523 22799 27529
rect 22741 27520 22753 27523
rect 21499 27492 22753 27520
rect 21499 27489 21511 27492
rect 21453 27483 21511 27489
rect 22741 27489 22753 27492
rect 22787 27489 22799 27523
rect 23290 27520 23296 27532
rect 23251 27492 23296 27520
rect 22741 27483 22799 27489
rect 9582 27452 9588 27464
rect 9543 27424 9588 27452
rect 9582 27412 9588 27424
rect 9640 27412 9646 27464
rect 10873 27455 10931 27461
rect 10873 27421 10885 27455
rect 10919 27421 10931 27455
rect 10873 27415 10931 27421
rect 10888 27384 10916 27415
rect 10962 27412 10968 27464
rect 11020 27452 11026 27464
rect 11057 27455 11115 27461
rect 11057 27452 11069 27455
rect 11020 27424 11069 27452
rect 11020 27412 11026 27424
rect 11057 27421 11069 27424
rect 11103 27421 11115 27455
rect 11057 27415 11115 27421
rect 11977 27455 12035 27461
rect 11977 27421 11989 27455
rect 12023 27452 12035 27455
rect 12618 27452 12624 27464
rect 12023 27424 12624 27452
rect 12023 27421 12035 27424
rect 11977 27415 12035 27421
rect 12618 27412 12624 27424
rect 12676 27412 12682 27464
rect 13354 27452 13360 27464
rect 13315 27424 13360 27452
rect 13354 27412 13360 27424
rect 13412 27412 13418 27464
rect 14090 27452 14096 27464
rect 14051 27424 14096 27452
rect 14090 27412 14096 27424
rect 14148 27412 14154 27464
rect 16390 27452 16396 27464
rect 16351 27424 16396 27452
rect 16390 27412 16396 27424
rect 16448 27412 16454 27464
rect 17770 27412 17776 27464
rect 17828 27452 17834 27464
rect 17865 27455 17923 27461
rect 17865 27452 17877 27455
rect 17828 27424 17877 27452
rect 17828 27412 17834 27424
rect 17865 27421 17877 27424
rect 17911 27421 17923 27455
rect 17865 27415 17923 27421
rect 20441 27455 20499 27461
rect 20441 27421 20453 27455
rect 20487 27421 20499 27455
rect 20441 27415 20499 27421
rect 20717 27455 20775 27461
rect 20717 27421 20729 27455
rect 20763 27452 20775 27455
rect 21082 27452 21088 27464
rect 20763 27424 21088 27452
rect 20763 27421 20775 27424
rect 20717 27415 20775 27421
rect 11514 27384 11520 27396
rect 10888 27356 11520 27384
rect 11514 27344 11520 27356
rect 11572 27344 11578 27396
rect 13449 27387 13507 27393
rect 13449 27353 13461 27387
rect 13495 27384 13507 27387
rect 14277 27387 14335 27393
rect 14277 27384 14289 27387
rect 13495 27356 14289 27384
rect 13495 27353 13507 27356
rect 13449 27347 13507 27353
rect 14277 27353 14289 27356
rect 14323 27353 14335 27387
rect 20456 27384 20484 27415
rect 21082 27412 21088 27424
rect 21140 27412 21146 27464
rect 21266 27412 21272 27464
rect 21324 27452 21330 27464
rect 21637 27455 21695 27461
rect 21637 27452 21649 27455
rect 21324 27424 21649 27452
rect 21324 27412 21330 27424
rect 21637 27421 21649 27424
rect 21683 27421 21695 27455
rect 22370 27452 22376 27464
rect 22331 27424 22376 27452
rect 21637 27415 21695 27421
rect 22370 27412 22376 27424
rect 22428 27412 22434 27464
rect 22756 27452 22784 27483
rect 23290 27480 23296 27492
rect 23348 27480 23354 27532
rect 23201 27455 23259 27461
rect 23201 27452 23213 27455
rect 22480 27424 22692 27452
rect 22756 27424 23213 27452
rect 20456 27356 21312 27384
rect 14277 27347 14335 27353
rect 10870 27276 10876 27328
rect 10928 27316 10934 27328
rect 10965 27319 11023 27325
rect 10965 27316 10977 27319
rect 10928 27288 10977 27316
rect 10928 27276 10934 27288
rect 10965 27285 10977 27288
rect 11011 27285 11023 27319
rect 10965 27279 11023 27285
rect 13630 27276 13636 27328
rect 13688 27316 13694 27328
rect 15378 27316 15384 27328
rect 13688 27288 15384 27316
rect 13688 27276 13694 27288
rect 15378 27276 15384 27288
rect 15436 27316 15442 27328
rect 16482 27316 16488 27328
rect 15436 27288 16488 27316
rect 15436 27276 15442 27288
rect 16482 27276 16488 27288
rect 16540 27276 16546 27328
rect 17957 27319 18015 27325
rect 17957 27285 17969 27319
rect 18003 27316 18015 27319
rect 18046 27316 18052 27328
rect 18003 27288 18052 27316
rect 18003 27285 18015 27288
rect 17957 27279 18015 27285
rect 18046 27276 18052 27288
rect 18104 27276 18110 27328
rect 20898 27316 20904 27328
rect 20859 27288 20904 27316
rect 20898 27276 20904 27288
rect 20956 27276 20962 27328
rect 21284 27316 21312 27356
rect 21358 27344 21364 27396
rect 21416 27384 21422 27396
rect 22480 27384 22508 27424
rect 21416 27356 21461 27384
rect 21836 27356 22508 27384
rect 22557 27387 22615 27393
rect 21416 27344 21422 27356
rect 21836 27328 21864 27356
rect 22557 27353 22569 27387
rect 22603 27353 22615 27387
rect 22664 27384 22692 27424
rect 23201 27421 23213 27424
rect 23247 27421 23259 27455
rect 24854 27452 24860 27464
rect 24815 27424 24860 27452
rect 23201 27415 23259 27421
rect 24854 27412 24860 27424
rect 24912 27412 24918 27464
rect 26142 27452 26148 27464
rect 26103 27424 26148 27452
rect 26142 27412 26148 27424
rect 26200 27412 26206 27464
rect 27062 27412 27068 27464
rect 27120 27452 27126 27464
rect 27540 27452 27568 27560
rect 29086 27548 29092 27560
rect 29144 27588 29150 27600
rect 30742 27588 30748 27600
rect 29144 27560 29868 27588
rect 30703 27560 30748 27588
rect 29144 27548 29150 27560
rect 27614 27480 27620 27532
rect 27672 27520 27678 27532
rect 27672 27492 29776 27520
rect 27672 27480 27678 27492
rect 28276 27464 28304 27492
rect 27893 27455 27951 27461
rect 27893 27452 27905 27455
rect 27120 27424 27905 27452
rect 27120 27412 27126 27424
rect 27893 27421 27905 27424
rect 27939 27421 27951 27455
rect 27893 27415 27951 27421
rect 28077 27455 28135 27461
rect 28077 27421 28089 27455
rect 28123 27452 28135 27455
rect 28258 27452 28264 27464
rect 28123 27424 28264 27452
rect 28123 27421 28135 27424
rect 28077 27415 28135 27421
rect 28258 27412 28264 27424
rect 28316 27412 28322 27464
rect 28534 27412 28540 27464
rect 28592 27452 28598 27464
rect 29748 27461 29776 27492
rect 29840 27464 29868 27560
rect 30742 27548 30748 27560
rect 30800 27548 30806 27600
rect 32125 27591 32183 27597
rect 32125 27557 32137 27591
rect 32171 27588 32183 27591
rect 33226 27588 33232 27600
rect 32171 27560 33232 27588
rect 32171 27557 32183 27560
rect 32125 27551 32183 27557
rect 33226 27548 33232 27560
rect 33284 27548 33290 27600
rect 46934 27588 46940 27600
rect 46308 27560 46940 27588
rect 31110 27520 31116 27532
rect 30208 27492 31116 27520
rect 29549 27455 29607 27461
rect 29549 27452 29561 27455
rect 28592 27424 29561 27452
rect 28592 27412 28598 27424
rect 29549 27421 29561 27424
rect 29595 27421 29607 27455
rect 29549 27415 29607 27421
rect 29733 27455 29791 27461
rect 29733 27421 29745 27455
rect 29779 27421 29791 27455
rect 29733 27415 29791 27421
rect 29822 27412 29828 27464
rect 29880 27452 29886 27464
rect 30101 27455 30159 27461
rect 30101 27452 30113 27455
rect 29880 27424 30113 27452
rect 29880 27412 29886 27424
rect 30101 27421 30113 27424
rect 30147 27421 30159 27455
rect 30101 27415 30159 27421
rect 22664 27356 24900 27384
rect 22557 27347 22615 27353
rect 21634 27316 21640 27328
rect 21284 27288 21640 27316
rect 21634 27276 21640 27288
rect 21692 27276 21698 27328
rect 21818 27316 21824 27328
rect 21779 27288 21824 27316
rect 21818 27276 21824 27288
rect 21876 27276 21882 27328
rect 22094 27276 22100 27328
rect 22152 27316 22158 27328
rect 22572 27316 22600 27347
rect 22152 27288 22600 27316
rect 24872 27316 24900 27356
rect 24946 27344 24952 27396
rect 25004 27384 25010 27396
rect 25041 27387 25099 27393
rect 25041 27384 25053 27387
rect 25004 27356 25053 27384
rect 25004 27344 25010 27356
rect 25041 27353 25053 27356
rect 25087 27384 25099 27387
rect 25130 27384 25136 27396
rect 25087 27356 25136 27384
rect 25087 27353 25099 27356
rect 25041 27347 25099 27353
rect 25130 27344 25136 27356
rect 25188 27344 25194 27396
rect 26694 27384 26700 27396
rect 25240 27356 26700 27384
rect 25240 27316 25268 27356
rect 26694 27344 26700 27356
rect 26752 27384 26758 27396
rect 26881 27387 26939 27393
rect 26881 27384 26893 27387
rect 26752 27356 26893 27384
rect 26752 27344 26758 27356
rect 26881 27353 26893 27356
rect 26927 27353 26939 27387
rect 26881 27347 26939 27353
rect 27709 27387 27767 27393
rect 27709 27353 27721 27387
rect 27755 27384 27767 27387
rect 27982 27384 27988 27396
rect 27755 27356 27988 27384
rect 27755 27353 27767 27356
rect 27709 27347 27767 27353
rect 27982 27344 27988 27356
rect 28040 27344 28046 27396
rect 28166 27384 28172 27396
rect 28127 27356 28172 27384
rect 28166 27344 28172 27356
rect 28224 27344 28230 27396
rect 28718 27384 28724 27396
rect 28679 27356 28724 27384
rect 28718 27344 28724 27356
rect 28776 27344 28782 27396
rect 28905 27387 28963 27393
rect 28905 27353 28917 27387
rect 28951 27384 28963 27387
rect 30208 27384 30236 27492
rect 31110 27480 31116 27492
rect 31168 27480 31174 27532
rect 46308 27529 46336 27560
rect 46934 27548 46940 27560
rect 46992 27548 46998 27600
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27489 46351 27523
rect 46293 27483 46351 27489
rect 46477 27523 46535 27529
rect 46477 27489 46489 27523
rect 46523 27520 46535 27523
rect 47670 27520 47676 27532
rect 46523 27492 47676 27520
rect 46523 27489 46535 27492
rect 46477 27483 46535 27489
rect 47670 27480 47676 27492
rect 47728 27480 47734 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 30561 27455 30619 27461
rect 30561 27421 30573 27455
rect 30607 27421 30619 27455
rect 30561 27415 30619 27421
rect 28951 27356 30236 27384
rect 28951 27353 28963 27356
rect 28905 27347 28963 27353
rect 26234 27316 26240 27328
rect 24872 27288 25268 27316
rect 26195 27288 26240 27316
rect 22152 27276 22158 27288
rect 26234 27276 26240 27288
rect 26292 27276 26298 27328
rect 28442 27276 28448 27328
rect 28500 27316 28506 27328
rect 28920 27316 28948 27347
rect 28500 27288 28948 27316
rect 30009 27319 30067 27325
rect 28500 27276 28506 27288
rect 30009 27285 30021 27319
rect 30055 27316 30067 27319
rect 30576 27316 30604 27415
rect 31018 27412 31024 27464
rect 31076 27452 31082 27464
rect 31662 27461 31668 27464
rect 31481 27455 31539 27461
rect 31481 27452 31493 27455
rect 31076 27424 31493 27452
rect 31076 27412 31082 27424
rect 31481 27421 31493 27424
rect 31527 27421 31539 27455
rect 31481 27415 31539 27421
rect 31629 27455 31668 27461
rect 31629 27421 31641 27455
rect 31629 27415 31668 27421
rect 31662 27412 31668 27415
rect 31720 27412 31726 27464
rect 31938 27452 31944 27464
rect 31996 27461 32002 27464
rect 31904 27424 31944 27452
rect 31938 27412 31944 27424
rect 31996 27415 32004 27461
rect 31996 27412 32002 27415
rect 30742 27344 30748 27396
rect 30800 27384 30806 27396
rect 31294 27384 31300 27396
rect 30800 27356 31300 27384
rect 30800 27344 30806 27356
rect 31294 27344 31300 27356
rect 31352 27384 31358 27396
rect 31757 27387 31815 27393
rect 31757 27384 31769 27387
rect 31352 27356 31769 27384
rect 31352 27344 31358 27356
rect 31757 27353 31769 27356
rect 31803 27353 31815 27387
rect 31757 27347 31815 27353
rect 31846 27344 31852 27396
rect 31904 27384 31910 27396
rect 31904 27356 31949 27384
rect 31904 27344 31910 27356
rect 30650 27316 30656 27328
rect 30055 27288 30656 27316
rect 30055 27285 30067 27288
rect 30009 27279 30067 27285
rect 30650 27276 30656 27288
rect 30708 27276 30714 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 10962 27072 10968 27124
rect 11020 27112 11026 27124
rect 13630 27112 13636 27124
rect 11020 27084 13636 27112
rect 11020 27072 11026 27084
rect 13630 27072 13636 27084
rect 13688 27072 13694 27124
rect 15286 27112 15292 27124
rect 15199 27084 15292 27112
rect 15286 27072 15292 27084
rect 15344 27112 15350 27124
rect 15930 27112 15936 27124
rect 15344 27084 15936 27112
rect 15344 27072 15350 27084
rect 15930 27072 15936 27084
rect 15988 27072 15994 27124
rect 17221 27115 17279 27121
rect 17221 27081 17233 27115
rect 17267 27112 17279 27115
rect 17310 27112 17316 27124
rect 17267 27084 17316 27112
rect 17267 27081 17279 27084
rect 17221 27075 17279 27081
rect 17310 27072 17316 27084
rect 17368 27072 17374 27124
rect 19242 27072 19248 27124
rect 19300 27112 19306 27124
rect 21818 27112 21824 27124
rect 19300 27084 21824 27112
rect 19300 27072 19306 27084
rect 21818 27072 21824 27084
rect 21876 27072 21882 27124
rect 24486 27072 24492 27124
rect 24544 27112 24550 27124
rect 26142 27112 26148 27124
rect 24544 27084 26148 27112
rect 24544 27072 24550 27084
rect 26142 27072 26148 27084
rect 26200 27072 26206 27124
rect 27246 27072 27252 27124
rect 27304 27112 27310 27124
rect 27817 27115 27875 27121
rect 27817 27112 27829 27115
rect 27304 27084 27829 27112
rect 27304 27072 27310 27084
rect 27817 27081 27829 27084
rect 27863 27112 27875 27115
rect 28534 27112 28540 27124
rect 27863 27084 28540 27112
rect 27863 27081 27875 27084
rect 27817 27075 27875 27081
rect 28534 27072 28540 27084
rect 28592 27072 28598 27124
rect 28629 27115 28687 27121
rect 28629 27081 28641 27115
rect 28675 27112 28687 27115
rect 28718 27112 28724 27124
rect 28675 27084 28724 27112
rect 28675 27081 28687 27084
rect 28629 27075 28687 27081
rect 28718 27072 28724 27084
rect 28776 27072 28782 27124
rect 29270 27112 29276 27124
rect 29231 27084 29276 27112
rect 29270 27072 29276 27084
rect 29328 27072 29334 27124
rect 30837 27115 30895 27121
rect 30837 27081 30849 27115
rect 30883 27112 30895 27115
rect 31294 27112 31300 27124
rect 30883 27084 31300 27112
rect 30883 27081 30895 27084
rect 30837 27075 30895 27081
rect 31294 27072 31300 27084
rect 31352 27112 31358 27124
rect 31352 27084 32352 27112
rect 31352 27072 31358 27084
rect 7466 27004 7472 27056
rect 7524 27044 7530 27056
rect 18046 27044 18052 27056
rect 7524 27016 17264 27044
rect 18007 27016 18052 27044
rect 7524 27004 7530 27016
rect 10689 26979 10747 26985
rect 10689 26945 10701 26979
rect 10735 26976 10747 26979
rect 10778 26976 10784 26988
rect 10735 26948 10784 26976
rect 10735 26945 10747 26948
rect 10689 26939 10747 26945
rect 10778 26936 10784 26948
rect 10836 26976 10842 26988
rect 10962 26976 10968 26988
rect 10836 26948 10968 26976
rect 10836 26936 10842 26948
rect 10962 26936 10968 26948
rect 11020 26936 11026 26988
rect 11609 26979 11667 26985
rect 11609 26945 11621 26979
rect 11655 26976 11667 26979
rect 12618 26976 12624 26988
rect 11655 26948 12624 26976
rect 11655 26945 11667 26948
rect 11609 26939 11667 26945
rect 12618 26936 12624 26948
rect 12676 26936 12682 26988
rect 13906 26976 13912 26988
rect 13867 26948 13912 26976
rect 13906 26936 13912 26948
rect 13964 26936 13970 26988
rect 14090 26936 14096 26988
rect 14148 26976 14154 26988
rect 14918 26976 14924 26988
rect 14148 26948 14924 26976
rect 14148 26936 14154 26948
rect 14918 26936 14924 26948
rect 14976 26976 14982 26988
rect 15105 26979 15163 26985
rect 15105 26976 15117 26979
rect 14976 26948 15117 26976
rect 14976 26936 14982 26948
rect 15105 26945 15117 26948
rect 15151 26945 15163 26979
rect 15378 26976 15384 26988
rect 15339 26948 15384 26976
rect 15105 26939 15163 26945
rect 15378 26936 15384 26948
rect 15436 26936 15442 26988
rect 15841 26979 15899 26985
rect 15841 26945 15853 26979
rect 15887 26976 15899 26979
rect 16390 26976 16396 26988
rect 15887 26948 16396 26976
rect 15887 26945 15899 26948
rect 15841 26939 15899 26945
rect 15194 26868 15200 26920
rect 15252 26908 15258 26920
rect 15856 26908 15884 26939
rect 16390 26936 16396 26948
rect 16448 26936 16454 26988
rect 16666 26936 16672 26988
rect 16724 26976 16730 26988
rect 17129 26979 17187 26985
rect 17129 26976 17141 26979
rect 16724 26948 17141 26976
rect 16724 26936 16730 26948
rect 17129 26945 17141 26948
rect 17175 26945 17187 26979
rect 17129 26939 17187 26945
rect 15252 26880 15884 26908
rect 17236 26908 17264 27016
rect 18046 27004 18052 27016
rect 18104 27004 18110 27056
rect 20622 27004 20628 27056
rect 20680 27044 20686 27056
rect 23106 27044 23112 27056
rect 20680 27016 23112 27044
rect 20680 27004 20686 27016
rect 17862 26976 17868 26988
rect 17823 26948 17868 26976
rect 17862 26936 17868 26948
rect 17920 26936 17926 26988
rect 20732 26985 20760 27016
rect 23106 27004 23112 27016
rect 23164 27004 23170 27056
rect 27614 27044 27620 27056
rect 23952 27016 25912 27044
rect 27575 27016 27620 27044
rect 20717 26979 20775 26985
rect 19260 26948 20668 26976
rect 19260 26908 19288 26948
rect 17236 26880 19288 26908
rect 19705 26911 19763 26917
rect 15252 26868 15258 26880
rect 19705 26877 19717 26911
rect 19751 26908 19763 26911
rect 20070 26908 20076 26920
rect 19751 26880 20076 26908
rect 19751 26877 19763 26880
rect 19705 26871 19763 26877
rect 20070 26868 20076 26880
rect 20128 26868 20134 26920
rect 20640 26908 20668 26948
rect 20717 26945 20729 26979
rect 20763 26945 20775 26979
rect 20717 26939 20775 26945
rect 20898 26936 20904 26988
rect 20956 26976 20962 26988
rect 21821 26979 21879 26985
rect 21821 26976 21833 26979
rect 20956 26948 21833 26976
rect 20956 26936 20962 26948
rect 21821 26945 21833 26948
rect 21867 26945 21879 26979
rect 22002 26976 22008 26988
rect 21963 26948 22008 26976
rect 21821 26939 21879 26945
rect 22002 26936 22008 26948
rect 22060 26936 22066 26988
rect 22094 26936 22100 26988
rect 22152 26976 22158 26988
rect 22373 26979 22431 26985
rect 22152 26948 22197 26976
rect 22152 26936 22158 26948
rect 22373 26945 22385 26979
rect 22419 26976 22431 26979
rect 22646 26976 22652 26988
rect 22419 26948 22652 26976
rect 22419 26945 22431 26948
rect 22373 26939 22431 26945
rect 22646 26936 22652 26948
rect 22704 26976 22710 26988
rect 23952 26976 23980 27016
rect 22704 26948 23980 26976
rect 24029 26979 24087 26985
rect 22704 26936 22710 26948
rect 24029 26945 24041 26979
rect 24075 26945 24087 26979
rect 24302 26976 24308 26988
rect 24263 26948 24308 26976
rect 24029 26939 24087 26945
rect 22189 26911 22247 26917
rect 22189 26908 22201 26911
rect 20640 26880 22201 26908
rect 22189 26877 22201 26880
rect 22235 26877 22247 26911
rect 24044 26908 24072 26939
rect 24302 26936 24308 26948
rect 24360 26936 24366 26988
rect 25682 26976 25688 26988
rect 25643 26948 25688 26976
rect 25682 26936 25688 26948
rect 25740 26936 25746 26988
rect 24854 26908 24860 26920
rect 24044 26880 24860 26908
rect 22189 26871 22247 26877
rect 24854 26868 24860 26880
rect 24912 26868 24918 26920
rect 9582 26800 9588 26852
rect 9640 26840 9646 26852
rect 9640 26812 12434 26840
rect 9640 26800 9646 26812
rect 10594 26732 10600 26784
rect 10652 26772 10658 26784
rect 10689 26775 10747 26781
rect 10689 26772 10701 26775
rect 10652 26744 10701 26772
rect 10652 26732 10658 26744
rect 10689 26741 10701 26744
rect 10735 26741 10747 26775
rect 10689 26735 10747 26741
rect 11606 26732 11612 26784
rect 11664 26772 11670 26784
rect 11701 26775 11759 26781
rect 11701 26772 11713 26775
rect 11664 26744 11713 26772
rect 11664 26732 11670 26744
rect 11701 26741 11713 26744
rect 11747 26741 11759 26775
rect 12406 26772 12434 26812
rect 14550 26800 14556 26852
rect 14608 26840 14614 26852
rect 24121 26843 24179 26849
rect 14608 26812 15976 26840
rect 14608 26800 14614 26812
rect 14093 26775 14151 26781
rect 14093 26772 14105 26775
rect 12406 26744 14105 26772
rect 11701 26735 11759 26741
rect 14093 26741 14105 26744
rect 14139 26741 14151 26775
rect 14093 26735 14151 26741
rect 15105 26775 15163 26781
rect 15105 26741 15117 26775
rect 15151 26772 15163 26775
rect 15654 26772 15660 26784
rect 15151 26744 15660 26772
rect 15151 26741 15163 26744
rect 15105 26735 15163 26741
rect 15654 26732 15660 26744
rect 15712 26732 15718 26784
rect 15838 26772 15844 26784
rect 15799 26744 15844 26772
rect 15838 26732 15844 26744
rect 15896 26732 15902 26784
rect 15948 26772 15976 26812
rect 24121 26809 24133 26843
rect 24167 26809 24179 26843
rect 24121 26803 24179 26809
rect 20622 26772 20628 26784
rect 15948 26744 20628 26772
rect 20622 26732 20628 26744
rect 20680 26732 20686 26784
rect 20806 26772 20812 26784
rect 20767 26744 20812 26772
rect 20806 26732 20812 26744
rect 20864 26732 20870 26784
rect 22554 26772 22560 26784
rect 22515 26744 22560 26772
rect 22554 26732 22560 26744
rect 22612 26732 22618 26784
rect 23842 26772 23848 26784
rect 23803 26744 23848 26772
rect 23842 26732 23848 26744
rect 23900 26732 23906 26784
rect 24136 26772 24164 26803
rect 24210 26800 24216 26852
rect 24268 26840 24274 26852
rect 24670 26840 24676 26852
rect 24268 26812 24676 26840
rect 24268 26800 24274 26812
rect 24670 26800 24676 26812
rect 24728 26800 24734 26852
rect 24578 26772 24584 26784
rect 24136 26744 24584 26772
rect 24578 26732 24584 26744
rect 24636 26732 24642 26784
rect 25884 26781 25912 27016
rect 27614 27004 27620 27016
rect 27672 27004 27678 27056
rect 27982 27004 27988 27056
rect 28040 27044 28046 27056
rect 31018 27044 31024 27056
rect 28040 27016 31024 27044
rect 28040 27004 28046 27016
rect 31018 27004 31024 27016
rect 31076 27004 31082 27056
rect 31110 27004 31116 27056
rect 31168 27044 31174 27056
rect 31168 27016 31754 27044
rect 31168 27004 31174 27016
rect 28537 26979 28595 26985
rect 28537 26976 28549 26979
rect 27908 26948 28549 26976
rect 27246 26868 27252 26920
rect 27304 26908 27310 26920
rect 27908 26908 27936 26948
rect 28537 26945 28549 26948
rect 28583 26945 28595 26979
rect 29178 26976 29184 26988
rect 29139 26948 29184 26976
rect 28537 26939 28595 26945
rect 29178 26936 29184 26948
rect 29236 26936 29242 26988
rect 30834 26979 30892 26985
rect 30834 26976 30846 26979
rect 29288 26948 30846 26976
rect 27304 26880 27936 26908
rect 27304 26868 27310 26880
rect 27982 26868 27988 26920
rect 28040 26908 28046 26920
rect 28626 26908 28632 26920
rect 28040 26880 28632 26908
rect 28040 26868 28046 26880
rect 28626 26868 28632 26880
rect 28684 26908 28690 26920
rect 29288 26908 29316 26948
rect 30834 26945 30846 26948
rect 30880 26976 30892 26979
rect 31202 26976 31208 26988
rect 30880 26948 31208 26976
rect 30880 26945 30892 26948
rect 30834 26939 30892 26945
rect 31202 26936 31208 26948
rect 31260 26936 31266 26988
rect 28684 26880 29316 26908
rect 31297 26911 31355 26917
rect 28684 26868 28690 26880
rect 31297 26877 31309 26911
rect 31343 26908 31355 26911
rect 31570 26908 31576 26920
rect 31343 26880 31576 26908
rect 31343 26877 31355 26880
rect 31297 26871 31355 26877
rect 31570 26868 31576 26880
rect 31628 26868 31634 26920
rect 31726 26908 31754 27016
rect 32324 26985 32352 27084
rect 33134 27004 33140 27056
rect 33192 27044 33198 27056
rect 33502 27044 33508 27056
rect 33192 27016 33508 27044
rect 33192 27004 33198 27016
rect 33502 27004 33508 27016
rect 33560 27044 33566 27056
rect 33560 27016 33640 27044
rect 33560 27004 33566 27016
rect 32309 26979 32367 26985
rect 32309 26945 32321 26979
rect 32355 26945 32367 26979
rect 32309 26939 32367 26945
rect 32401 26979 32459 26985
rect 32401 26945 32413 26979
rect 32447 26976 32459 26979
rect 32490 26976 32496 26988
rect 32447 26948 32496 26976
rect 32447 26945 32459 26948
rect 32401 26939 32459 26945
rect 32490 26936 32496 26948
rect 32548 26936 32554 26988
rect 32585 26979 32643 26985
rect 32585 26945 32597 26979
rect 32631 26945 32643 26979
rect 32585 26939 32643 26945
rect 32677 26979 32735 26985
rect 32677 26945 32689 26979
rect 32723 26945 32735 26979
rect 33410 26976 33416 26988
rect 33371 26948 33416 26976
rect 32677 26939 32735 26945
rect 32600 26908 32628 26939
rect 31726 26880 32628 26908
rect 26234 26800 26240 26852
rect 26292 26840 26298 26852
rect 32692 26840 32720 26939
rect 33410 26936 33416 26948
rect 33468 26936 33474 26988
rect 33612 26985 33640 27016
rect 33597 26979 33655 26985
rect 33597 26945 33609 26979
rect 33643 26945 33655 26979
rect 33962 26976 33968 26988
rect 33923 26948 33968 26976
rect 33597 26939 33655 26945
rect 33962 26936 33968 26948
rect 34020 26936 34026 26988
rect 32950 26868 32956 26920
rect 33008 26908 33014 26920
rect 33689 26911 33747 26917
rect 33689 26908 33701 26911
rect 33008 26880 33701 26908
rect 33008 26868 33014 26880
rect 33689 26877 33701 26880
rect 33735 26877 33747 26911
rect 33689 26871 33747 26877
rect 33781 26911 33839 26917
rect 33781 26877 33793 26911
rect 33827 26908 33839 26911
rect 40402 26908 40408 26920
rect 33827 26880 40408 26908
rect 33827 26877 33839 26880
rect 33781 26871 33839 26877
rect 40402 26868 40408 26880
rect 40460 26868 40466 26920
rect 26292 26812 32720 26840
rect 26292 26800 26298 26812
rect 25869 26775 25927 26781
rect 25869 26741 25881 26775
rect 25915 26772 25927 26775
rect 27338 26772 27344 26784
rect 25915 26744 27344 26772
rect 25915 26741 25927 26744
rect 25869 26735 25927 26741
rect 27338 26732 27344 26744
rect 27396 26732 27402 26784
rect 27798 26772 27804 26784
rect 27759 26744 27804 26772
rect 27798 26732 27804 26744
rect 27856 26732 27862 26784
rect 27982 26772 27988 26784
rect 27943 26744 27988 26772
rect 27982 26732 27988 26744
rect 28040 26732 28046 26784
rect 29914 26732 29920 26784
rect 29972 26772 29978 26784
rect 30653 26775 30711 26781
rect 30653 26772 30665 26775
rect 29972 26744 30665 26772
rect 29972 26732 29978 26744
rect 30653 26741 30665 26744
rect 30699 26741 30711 26775
rect 30653 26735 30711 26741
rect 31018 26732 31024 26784
rect 31076 26772 31082 26784
rect 31205 26775 31263 26781
rect 31205 26772 31217 26775
rect 31076 26744 31217 26772
rect 31076 26732 31082 26744
rect 31205 26741 31217 26744
rect 31251 26741 31263 26775
rect 31205 26735 31263 26741
rect 32125 26775 32183 26781
rect 32125 26741 32137 26775
rect 32171 26772 32183 26775
rect 33318 26772 33324 26784
rect 32171 26744 33324 26772
rect 32171 26741 32183 26744
rect 32125 26735 32183 26741
rect 33318 26732 33324 26744
rect 33376 26732 33382 26784
rect 34149 26775 34207 26781
rect 34149 26741 34161 26775
rect 34195 26772 34207 26775
rect 34698 26772 34704 26784
rect 34195 26744 34704 26772
rect 34195 26741 34207 26744
rect 34149 26735 34207 26741
rect 34698 26732 34704 26744
rect 34756 26732 34762 26784
rect 46290 26732 46296 26784
rect 46348 26772 46354 26784
rect 47765 26775 47823 26781
rect 47765 26772 47777 26775
rect 46348 26744 47777 26772
rect 46348 26732 46354 26744
rect 47765 26741 47777 26744
rect 47811 26741 47823 26775
rect 47765 26735 47823 26741
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 11330 26528 11336 26580
rect 11388 26568 11394 26580
rect 12342 26568 12348 26580
rect 11388 26540 12348 26568
rect 11388 26528 11394 26540
rect 12342 26528 12348 26540
rect 12400 26528 12406 26580
rect 14553 26571 14611 26577
rect 14553 26537 14565 26571
rect 14599 26568 14611 26571
rect 14734 26568 14740 26580
rect 14599 26540 14740 26568
rect 14599 26537 14611 26540
rect 14553 26531 14611 26537
rect 14734 26528 14740 26540
rect 14792 26528 14798 26580
rect 14918 26528 14924 26580
rect 14976 26568 14982 26580
rect 16853 26571 16911 26577
rect 16853 26568 16865 26571
rect 14976 26540 16865 26568
rect 14976 26528 14982 26540
rect 16853 26537 16865 26540
rect 16899 26537 16911 26571
rect 16853 26531 16911 26537
rect 19784 26571 19842 26577
rect 19784 26537 19796 26571
rect 19830 26568 19842 26571
rect 22554 26568 22560 26580
rect 19830 26540 22560 26568
rect 19830 26537 19842 26540
rect 19784 26531 19842 26537
rect 22554 26528 22560 26540
rect 22612 26528 22618 26580
rect 24765 26571 24823 26577
rect 24765 26537 24777 26571
rect 24811 26537 24823 26571
rect 27062 26568 27068 26580
rect 27023 26540 27068 26568
rect 24765 26531 24823 26537
rect 22278 26500 22284 26512
rect 20824 26472 22284 26500
rect 10594 26432 10600 26444
rect 10555 26404 10600 26432
rect 10594 26392 10600 26404
rect 10652 26392 10658 26444
rect 10870 26432 10876 26444
rect 10831 26404 10876 26432
rect 10870 26392 10876 26404
rect 10928 26392 10934 26444
rect 15105 26435 15163 26441
rect 15105 26401 15117 26435
rect 15151 26432 15163 26435
rect 15838 26432 15844 26444
rect 15151 26404 15844 26432
rect 15151 26401 15163 26404
rect 15105 26395 15163 26401
rect 15838 26392 15844 26404
rect 15896 26392 15902 26444
rect 19426 26392 19432 26444
rect 19484 26432 19490 26444
rect 19521 26435 19579 26441
rect 19521 26432 19533 26435
rect 19484 26404 19533 26432
rect 19484 26392 19490 26404
rect 19521 26401 19533 26404
rect 19567 26432 19579 26435
rect 20824 26432 20852 26472
rect 22278 26460 22284 26472
rect 22336 26460 22342 26512
rect 24578 26460 24584 26512
rect 24636 26500 24642 26512
rect 24780 26500 24808 26531
rect 27062 26528 27068 26540
rect 27120 26528 27126 26580
rect 27246 26568 27252 26580
rect 27207 26540 27252 26568
rect 27246 26528 27252 26540
rect 27304 26528 27310 26580
rect 27982 26528 27988 26580
rect 28040 26568 28046 26580
rect 28261 26571 28319 26577
rect 28261 26568 28273 26571
rect 28040 26540 28273 26568
rect 28040 26528 28046 26540
rect 28261 26537 28273 26540
rect 28307 26537 28319 26571
rect 28261 26531 28319 26537
rect 28721 26571 28779 26577
rect 28721 26537 28733 26571
rect 28767 26568 28779 26571
rect 31386 26568 31392 26580
rect 28767 26540 31392 26568
rect 28767 26537 28779 26540
rect 28721 26531 28779 26537
rect 31386 26528 31392 26540
rect 31444 26528 31450 26580
rect 31570 26528 31576 26580
rect 31628 26568 31634 26580
rect 32401 26571 32459 26577
rect 32401 26568 32413 26571
rect 31628 26540 32413 26568
rect 31628 26528 31634 26540
rect 32401 26537 32413 26540
rect 32447 26537 32459 26571
rect 32401 26531 32459 26537
rect 27154 26500 27160 26512
rect 24636 26472 27160 26500
rect 24636 26460 24642 26472
rect 27154 26460 27160 26472
rect 27212 26460 27218 26512
rect 27338 26460 27344 26512
rect 27396 26500 27402 26512
rect 30101 26503 30159 26509
rect 27396 26472 28994 26500
rect 27396 26460 27402 26472
rect 19567 26404 20852 26432
rect 21269 26435 21327 26441
rect 19567 26401 19579 26404
rect 19521 26395 19579 26401
rect 21269 26401 21281 26435
rect 21315 26401 21327 26435
rect 21269 26395 21327 26401
rect 14182 26364 14188 26376
rect 14143 26336 14188 26364
rect 14182 26324 14188 26336
rect 14240 26324 14246 26376
rect 14369 26367 14427 26373
rect 14369 26333 14381 26367
rect 14415 26364 14427 26367
rect 14734 26364 14740 26376
rect 14415 26336 14740 26364
rect 14415 26333 14427 26336
rect 14369 26327 14427 26333
rect 14734 26324 14740 26336
rect 14792 26324 14798 26376
rect 21284 26364 21312 26395
rect 21634 26392 21640 26444
rect 21692 26432 21698 26444
rect 21821 26435 21879 26441
rect 21821 26432 21833 26435
rect 21692 26404 21833 26432
rect 21692 26392 21698 26404
rect 21821 26401 21833 26404
rect 21867 26401 21879 26435
rect 21821 26395 21879 26401
rect 21910 26392 21916 26444
rect 21968 26432 21974 26444
rect 23845 26435 23903 26441
rect 23845 26432 23857 26435
rect 21968 26404 23857 26432
rect 21968 26392 21974 26404
rect 23845 26401 23857 26404
rect 23891 26401 23903 26435
rect 28534 26432 28540 26444
rect 23845 26395 23903 26401
rect 24320 26404 24900 26432
rect 21729 26367 21787 26373
rect 21729 26364 21741 26367
rect 21284 26336 21741 26364
rect 21729 26333 21741 26336
rect 21775 26364 21787 26367
rect 22002 26364 22008 26376
rect 21775 26336 22008 26364
rect 21775 26333 21787 26336
rect 21729 26327 21787 26333
rect 22002 26324 22008 26336
rect 22060 26324 22066 26376
rect 23477 26367 23535 26373
rect 23477 26333 23489 26367
rect 23523 26364 23535 26367
rect 24320 26364 24348 26404
rect 24872 26376 24900 26404
rect 28194 26404 28540 26432
rect 24670 26364 24676 26376
rect 23523 26336 24348 26364
rect 24631 26336 24676 26364
rect 23523 26333 23535 26336
rect 23477 26327 23535 26333
rect 24670 26324 24676 26336
rect 24728 26324 24734 26376
rect 24854 26364 24860 26376
rect 24815 26336 24860 26364
rect 24854 26324 24860 26336
rect 24912 26324 24918 26376
rect 26694 26364 26700 26376
rect 26655 26336 26700 26364
rect 26694 26324 26700 26336
rect 26752 26324 26758 26376
rect 27065 26367 27123 26373
rect 27065 26333 27077 26367
rect 27111 26364 27123 26367
rect 27154 26364 27160 26376
rect 27111 26336 27160 26364
rect 27111 26333 27123 26336
rect 27065 26327 27123 26333
rect 27154 26324 27160 26336
rect 27212 26324 27218 26376
rect 28194 26373 28222 26404
rect 28534 26392 28540 26404
rect 28592 26392 28598 26444
rect 28169 26367 28227 26373
rect 28169 26333 28181 26367
rect 28215 26333 28227 26367
rect 28169 26327 28227 26333
rect 28445 26367 28503 26373
rect 28445 26333 28457 26367
rect 28491 26364 28503 26367
rect 28718 26364 28724 26376
rect 28491 26336 28724 26364
rect 28491 26333 28503 26336
rect 28445 26327 28503 26333
rect 28718 26324 28724 26336
rect 28776 26324 28782 26376
rect 28966 26364 28994 26472
rect 30101 26469 30113 26503
rect 30147 26500 30159 26503
rect 30374 26500 30380 26512
rect 30147 26472 30380 26500
rect 30147 26469 30159 26472
rect 30101 26463 30159 26469
rect 30374 26460 30380 26472
rect 30432 26460 30438 26512
rect 32490 26460 32496 26512
rect 32548 26500 32554 26512
rect 32548 26472 33640 26500
rect 32548 26460 32554 26472
rect 29638 26392 29644 26444
rect 29696 26432 29702 26444
rect 30653 26435 30711 26441
rect 29696 26404 29868 26432
rect 29696 26392 29702 26404
rect 29840 26373 29868 26404
rect 30653 26401 30665 26435
rect 30699 26432 30711 26435
rect 31018 26432 31024 26444
rect 30699 26404 31024 26432
rect 30699 26401 30711 26404
rect 30653 26395 30711 26401
rect 31018 26392 31024 26404
rect 31076 26392 31082 26444
rect 31386 26392 31392 26444
rect 31444 26432 31450 26444
rect 33410 26432 33416 26444
rect 31444 26404 33416 26432
rect 31444 26392 31450 26404
rect 33410 26392 33416 26404
rect 33468 26392 33474 26444
rect 33612 26376 33640 26472
rect 33686 26392 33692 26444
rect 33744 26432 33750 26444
rect 46290 26432 46296 26444
rect 33744 26404 33789 26432
rect 46251 26404 46296 26432
rect 33744 26392 33750 26404
rect 46290 26392 46296 26404
rect 46348 26392 46354 26444
rect 29825 26367 29883 26373
rect 28966 26336 29592 26364
rect 11606 26256 11612 26308
rect 11664 26256 11670 26308
rect 15378 26296 15384 26308
rect 15339 26268 15384 26296
rect 15378 26256 15384 26268
rect 15436 26256 15442 26308
rect 16022 26256 16028 26308
rect 16080 26256 16086 26308
rect 20806 26256 20812 26308
rect 20864 26256 20870 26308
rect 21082 26256 21088 26308
rect 21140 26296 21146 26308
rect 21140 26268 21312 26296
rect 21140 26256 21146 26268
rect 13354 26188 13360 26240
rect 13412 26228 13418 26240
rect 17770 26228 17776 26240
rect 13412 26200 17776 26228
rect 13412 26188 13418 26200
rect 17770 26188 17776 26200
rect 17828 26188 17834 26240
rect 21284 26228 21312 26268
rect 21358 26256 21364 26308
rect 21416 26296 21422 26308
rect 21910 26296 21916 26308
rect 21416 26268 21916 26296
rect 21416 26256 21422 26268
rect 21910 26256 21916 26268
rect 21968 26256 21974 26308
rect 23658 26296 23664 26308
rect 22020 26268 23520 26296
rect 23619 26268 23664 26296
rect 22020 26228 22048 26268
rect 21284 26200 22048 26228
rect 23492 26228 23520 26268
rect 23658 26256 23664 26268
rect 23716 26296 23722 26308
rect 24302 26296 24308 26308
rect 23716 26268 24308 26296
rect 23716 26256 23722 26268
rect 24302 26256 24308 26268
rect 24360 26296 24366 26308
rect 24397 26299 24455 26305
rect 24397 26296 24409 26299
rect 24360 26268 24409 26296
rect 24360 26256 24366 26268
rect 24397 26265 24409 26268
rect 24443 26265 24455 26299
rect 25498 26296 25504 26308
rect 24397 26259 24455 26265
rect 24504 26268 25504 26296
rect 24504 26228 24532 26268
rect 25498 26256 25504 26268
rect 25556 26256 25562 26308
rect 26326 26256 26332 26308
rect 26384 26296 26390 26308
rect 29178 26296 29184 26308
rect 26384 26268 29184 26296
rect 26384 26256 26390 26268
rect 29178 26256 29184 26268
rect 29236 26256 29242 26308
rect 25038 26228 25044 26240
rect 23492 26200 24532 26228
rect 24999 26200 25044 26228
rect 25038 26188 25044 26200
rect 25096 26188 25102 26240
rect 29564 26228 29592 26336
rect 29825 26333 29837 26367
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 29914 26324 29920 26376
rect 29972 26364 29978 26376
rect 30190 26373 30196 26376
rect 30175 26367 30196 26373
rect 29972 26336 30017 26364
rect 29972 26324 29978 26336
rect 30175 26333 30187 26367
rect 30175 26327 30196 26333
rect 30190 26324 30196 26327
rect 30248 26324 30254 26376
rect 33318 26364 33324 26376
rect 33279 26336 33324 26364
rect 33318 26324 33324 26336
rect 33376 26324 33382 26376
rect 33502 26364 33508 26376
rect 33463 26336 33508 26364
rect 33502 26324 33508 26336
rect 33560 26324 33566 26376
rect 33594 26324 33600 26376
rect 33652 26364 33658 26376
rect 33873 26367 33931 26373
rect 33652 26336 33697 26364
rect 33652 26324 33658 26336
rect 33873 26333 33885 26367
rect 33919 26364 33931 26367
rect 33962 26364 33968 26376
rect 33919 26336 33968 26364
rect 33919 26333 33931 26336
rect 33873 26327 33931 26333
rect 33962 26324 33968 26336
rect 34020 26324 34026 26376
rect 29641 26299 29699 26305
rect 29641 26265 29653 26299
rect 29687 26296 29699 26299
rect 30929 26299 30987 26305
rect 30929 26296 30941 26299
rect 29687 26268 30941 26296
rect 29687 26265 29699 26268
rect 29641 26259 29699 26265
rect 30929 26265 30941 26268
rect 30975 26265 30987 26299
rect 32582 26296 32588 26308
rect 32154 26268 32588 26296
rect 30929 26259 30987 26265
rect 32582 26256 32588 26268
rect 32640 26256 32646 26308
rect 46477 26299 46535 26305
rect 46477 26265 46489 26299
rect 46523 26296 46535 26299
rect 46842 26296 46848 26308
rect 46523 26268 46848 26296
rect 46523 26265 46535 26268
rect 46477 26259 46535 26265
rect 46842 26256 46848 26268
rect 46900 26256 46906 26308
rect 48133 26299 48191 26305
rect 48133 26265 48145 26299
rect 48179 26296 48191 26299
rect 48222 26296 48228 26308
rect 48179 26268 48228 26296
rect 48179 26265 48191 26268
rect 48133 26259 48191 26265
rect 48222 26256 48228 26268
rect 48280 26256 48286 26308
rect 30190 26228 30196 26240
rect 29564 26200 30196 26228
rect 30190 26188 30196 26200
rect 30248 26188 30254 26240
rect 34054 26228 34060 26240
rect 34015 26200 34060 26228
rect 34054 26188 34060 26200
rect 34112 26188 34118 26240
rect 46382 26188 46388 26240
rect 46440 26228 46446 26240
rect 46750 26228 46756 26240
rect 46440 26200 46756 26228
rect 46440 26188 46446 26200
rect 46750 26188 46756 26200
rect 46808 26188 46814 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 13265 26027 13323 26033
rect 13265 25993 13277 26027
rect 13311 26024 13323 26027
rect 14182 26024 14188 26036
rect 13311 25996 14188 26024
rect 13311 25993 13323 25996
rect 13265 25987 13323 25993
rect 14182 25984 14188 25996
rect 14240 26024 14246 26036
rect 15105 26027 15163 26033
rect 15105 26024 15117 26027
rect 14240 25996 15117 26024
rect 14240 25984 14246 25996
rect 15105 25993 15117 25996
rect 15151 25993 15163 26027
rect 15286 26024 15292 26036
rect 15247 25996 15292 26024
rect 15105 25987 15163 25993
rect 15286 25984 15292 25996
rect 15344 25984 15350 26036
rect 16022 26024 16028 26036
rect 15983 25996 16028 26024
rect 16022 25984 16028 25996
rect 16080 25984 16086 26036
rect 17405 26027 17463 26033
rect 17405 25993 17417 26027
rect 17451 26024 17463 26027
rect 17770 26024 17776 26036
rect 17451 25996 17776 26024
rect 17451 25993 17463 25996
rect 17405 25987 17463 25993
rect 17770 25984 17776 25996
rect 17828 25984 17834 26036
rect 23842 26024 23848 26036
rect 23803 25996 23848 26024
rect 23842 25984 23848 25996
rect 23900 25984 23906 26036
rect 25498 25984 25504 26036
rect 25556 26024 25562 26036
rect 28813 26027 28871 26033
rect 28813 26024 28825 26027
rect 25556 25996 28825 26024
rect 25556 25984 25562 25996
rect 28813 25993 28825 25996
rect 28859 25993 28871 26027
rect 28813 25987 28871 25993
rect 29638 25984 29644 26036
rect 29696 26024 29702 26036
rect 30469 26027 30527 26033
rect 30469 26024 30481 26027
rect 29696 25996 30481 26024
rect 29696 25984 29702 25996
rect 30469 25993 30481 25996
rect 30515 25993 30527 26027
rect 31294 26024 31300 26036
rect 31255 25996 31300 26024
rect 30469 25987 30527 25993
rect 31294 25984 31300 25996
rect 31352 25984 31358 26036
rect 32582 26024 32588 26036
rect 32543 25996 32588 26024
rect 32582 25984 32588 25996
rect 32640 25984 32646 26036
rect 33594 25984 33600 26036
rect 33652 26024 33658 26036
rect 35621 26027 35679 26033
rect 35621 26024 35633 26027
rect 33652 25996 35633 26024
rect 33652 25984 33658 25996
rect 35621 25993 35633 25996
rect 35667 25993 35679 26027
rect 35621 25987 35679 25993
rect 46109 26027 46167 26033
rect 46109 25993 46121 26027
rect 46155 26024 46167 26027
rect 47762 26024 47768 26036
rect 46155 25996 47768 26024
rect 46155 25993 46167 25996
rect 46109 25987 46167 25993
rect 47762 25984 47768 25996
rect 47820 25984 47826 26036
rect 11422 25916 11428 25968
rect 11480 25956 11486 25968
rect 11701 25959 11759 25965
rect 11701 25956 11713 25959
rect 11480 25928 11713 25956
rect 11480 25916 11486 25928
rect 11701 25925 11713 25928
rect 11747 25925 11759 25959
rect 11701 25919 11759 25925
rect 12342 25916 12348 25968
rect 12400 25956 12406 25968
rect 12897 25959 12955 25965
rect 12897 25956 12909 25959
rect 12400 25928 12909 25956
rect 12400 25916 12406 25928
rect 12897 25925 12909 25928
rect 12943 25925 12955 25959
rect 12897 25919 12955 25925
rect 13113 25959 13171 25965
rect 13113 25925 13125 25959
rect 13159 25956 13171 25959
rect 14274 25956 14280 25968
rect 13159 25928 14280 25956
rect 13159 25925 13171 25928
rect 13113 25919 13171 25925
rect 14274 25916 14280 25928
rect 14332 25916 14338 25968
rect 14918 25956 14924 25968
rect 14879 25928 14924 25956
rect 14918 25916 14924 25928
rect 14976 25916 14982 25968
rect 18049 25959 18107 25965
rect 18049 25925 18061 25959
rect 18095 25956 18107 25959
rect 30929 25959 30987 25965
rect 18095 25928 26924 25956
rect 18095 25925 18107 25928
rect 18049 25919 18107 25925
rect 9953 25891 10011 25897
rect 9953 25857 9965 25891
rect 9999 25888 10011 25891
rect 10962 25888 10968 25900
rect 9999 25860 10968 25888
rect 9999 25857 10011 25860
rect 9953 25851 10011 25857
rect 10962 25848 10968 25860
rect 11020 25848 11026 25900
rect 11330 25848 11336 25900
rect 11388 25888 11394 25900
rect 11517 25891 11575 25897
rect 11517 25888 11529 25891
rect 11388 25860 11529 25888
rect 11388 25848 11394 25860
rect 11517 25857 11529 25860
rect 11563 25857 11575 25891
rect 11517 25851 11575 25857
rect 11793 25891 11851 25897
rect 11793 25857 11805 25891
rect 11839 25888 11851 25891
rect 11882 25888 11888 25900
rect 11839 25860 11888 25888
rect 11839 25857 11851 25860
rect 11793 25851 11851 25857
rect 11882 25848 11888 25860
rect 11940 25848 11946 25900
rect 14182 25888 14188 25900
rect 14143 25860 14188 25888
rect 14182 25848 14188 25860
rect 14240 25848 14246 25900
rect 14734 25848 14740 25900
rect 14792 25888 14798 25900
rect 15197 25891 15255 25897
rect 15197 25888 15209 25891
rect 14792 25860 15209 25888
rect 14792 25848 14798 25860
rect 15197 25857 15209 25860
rect 15243 25857 15255 25891
rect 15197 25851 15255 25857
rect 15933 25891 15991 25897
rect 15933 25857 15945 25891
rect 15979 25888 15991 25891
rect 16666 25888 16672 25900
rect 15979 25860 16672 25888
rect 15979 25857 15991 25860
rect 15933 25851 15991 25857
rect 16666 25848 16672 25860
rect 16724 25848 16730 25900
rect 17218 25888 17224 25900
rect 17179 25860 17224 25888
rect 17218 25848 17224 25860
rect 17276 25888 17282 25900
rect 18233 25891 18291 25897
rect 18233 25888 18245 25891
rect 17276 25860 18245 25888
rect 17276 25848 17282 25860
rect 18233 25857 18245 25860
rect 18279 25857 18291 25891
rect 18233 25851 18291 25857
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25857 20867 25891
rect 20990 25888 20996 25900
rect 20951 25860 20996 25888
rect 20809 25851 20867 25857
rect 15473 25823 15531 25829
rect 15473 25789 15485 25823
rect 15519 25820 15531 25823
rect 20824 25820 20852 25851
rect 20990 25848 20996 25860
rect 21048 25848 21054 25900
rect 21266 25888 21272 25900
rect 21227 25860 21272 25888
rect 21266 25848 21272 25860
rect 21324 25848 21330 25900
rect 22925 25891 22983 25897
rect 22925 25857 22937 25891
rect 22971 25888 22983 25891
rect 23753 25891 23811 25897
rect 22971 25860 23428 25888
rect 22971 25857 22983 25860
rect 22925 25851 22983 25857
rect 15519 25792 20852 25820
rect 20901 25823 20959 25829
rect 15519 25789 15531 25792
rect 15473 25783 15531 25789
rect 20901 25789 20913 25823
rect 20947 25820 20959 25823
rect 21358 25820 21364 25832
rect 20947 25792 21364 25820
rect 20947 25789 20959 25792
rect 20901 25783 20959 25789
rect 21358 25780 21364 25792
rect 21416 25780 21422 25832
rect 11514 25752 11520 25764
rect 11475 25724 11520 25752
rect 11514 25712 11520 25724
rect 11572 25712 11578 25764
rect 14182 25712 14188 25764
rect 14240 25752 14246 25764
rect 19242 25752 19248 25764
rect 14240 25724 19248 25752
rect 14240 25712 14246 25724
rect 19242 25712 19248 25724
rect 19300 25712 19306 25764
rect 21085 25755 21143 25761
rect 21085 25721 21097 25755
rect 21131 25752 21143 25755
rect 21542 25752 21548 25764
rect 21131 25724 21548 25752
rect 21131 25721 21143 25724
rect 21085 25715 21143 25721
rect 21542 25712 21548 25724
rect 21600 25712 21606 25764
rect 23400 25761 23428 25860
rect 23753 25857 23765 25891
rect 23799 25888 23811 25891
rect 24210 25888 24216 25900
rect 23799 25860 24216 25888
rect 23799 25857 23811 25860
rect 23753 25851 23811 25857
rect 24210 25848 24216 25860
rect 24268 25848 24274 25900
rect 24578 25888 24584 25900
rect 24539 25860 24584 25888
rect 24578 25848 24584 25860
rect 24636 25848 24642 25900
rect 24670 25848 24676 25900
rect 24728 25888 24734 25900
rect 24728 25860 24773 25888
rect 24728 25848 24734 25860
rect 24029 25823 24087 25829
rect 24029 25789 24041 25823
rect 24075 25789 24087 25823
rect 24854 25820 24860 25832
rect 24815 25792 24860 25820
rect 24029 25783 24087 25789
rect 23385 25755 23443 25761
rect 23385 25721 23397 25755
rect 23431 25721 23443 25755
rect 24044 25752 24072 25783
rect 24854 25780 24860 25792
rect 24912 25780 24918 25832
rect 25682 25752 25688 25764
rect 24044 25724 25688 25752
rect 23385 25715 23443 25721
rect 25682 25712 25688 25724
rect 25740 25712 25746 25764
rect 26896 25752 26924 25928
rect 30929 25925 30941 25959
rect 30975 25956 30987 25959
rect 31386 25956 31392 25968
rect 30975 25928 31392 25956
rect 30975 25925 30987 25928
rect 30929 25919 30987 25925
rect 26973 25891 27031 25897
rect 26973 25857 26985 25891
rect 27019 25888 27031 25891
rect 27246 25888 27252 25900
rect 27019 25860 27252 25888
rect 27019 25857 27031 25860
rect 26973 25851 27031 25857
rect 27246 25848 27252 25860
rect 27304 25848 27310 25900
rect 28626 25888 28632 25900
rect 28587 25860 28632 25888
rect 28626 25848 28632 25860
rect 28684 25848 28690 25900
rect 30285 25891 30343 25897
rect 30285 25857 30297 25891
rect 30331 25888 30343 25891
rect 30944 25888 30972 25919
rect 31386 25916 31392 25928
rect 31444 25916 31450 25968
rect 34054 25916 34060 25968
rect 34112 25956 34118 25968
rect 34149 25959 34207 25965
rect 34149 25956 34161 25959
rect 34112 25928 34161 25956
rect 34112 25916 34118 25928
rect 34149 25925 34161 25928
rect 34195 25925 34207 25959
rect 34149 25919 34207 25925
rect 34606 25916 34612 25968
rect 34664 25916 34670 25968
rect 31113 25891 31171 25897
rect 31113 25888 31125 25891
rect 30331 25860 30972 25888
rect 31036 25860 31125 25888
rect 30331 25857 30343 25860
rect 30285 25851 30343 25857
rect 30101 25823 30159 25829
rect 30101 25789 30113 25823
rect 30147 25820 30159 25823
rect 31036 25820 31064 25860
rect 31113 25857 31125 25860
rect 31159 25888 31171 25891
rect 31570 25888 31576 25900
rect 31159 25860 31576 25888
rect 31159 25857 31171 25860
rect 31113 25851 31171 25857
rect 31570 25848 31576 25860
rect 31628 25848 31634 25900
rect 32493 25891 32551 25897
rect 32493 25857 32505 25891
rect 32539 25888 32551 25891
rect 33778 25888 33784 25900
rect 32539 25860 33784 25888
rect 32539 25857 32551 25860
rect 32493 25851 32551 25857
rect 33778 25848 33784 25860
rect 33836 25848 33842 25900
rect 46293 25891 46351 25897
rect 46293 25857 46305 25891
rect 46339 25888 46351 25891
rect 46658 25888 46664 25900
rect 46339 25860 46664 25888
rect 46339 25857 46351 25860
rect 46293 25851 46351 25857
rect 46658 25848 46664 25860
rect 46716 25848 46722 25900
rect 46753 25891 46811 25897
rect 46753 25857 46765 25891
rect 46799 25857 46811 25891
rect 46753 25851 46811 25857
rect 30147 25792 31064 25820
rect 30147 25789 30159 25792
rect 30101 25783 30159 25789
rect 31478 25780 31484 25832
rect 31536 25820 31542 25832
rect 33870 25820 33876 25832
rect 31536 25792 33876 25820
rect 31536 25780 31542 25792
rect 33870 25780 33876 25792
rect 33928 25780 33934 25832
rect 45830 25780 45836 25832
rect 45888 25820 45894 25832
rect 46382 25820 46388 25832
rect 45888 25792 46388 25820
rect 45888 25780 45894 25792
rect 46382 25780 46388 25792
rect 46440 25820 46446 25832
rect 46768 25820 46796 25851
rect 46440 25792 46796 25820
rect 46440 25780 46446 25792
rect 33042 25752 33048 25764
rect 26896 25724 33048 25752
rect 33042 25712 33048 25724
rect 33100 25712 33106 25764
rect 46290 25712 46296 25764
rect 46348 25752 46354 25764
rect 47765 25755 47823 25761
rect 47765 25752 47777 25755
rect 46348 25724 47777 25752
rect 46348 25712 46354 25724
rect 47765 25721 47777 25724
rect 47811 25721 47823 25755
rect 47765 25715 47823 25721
rect 9674 25644 9680 25696
rect 9732 25684 9738 25696
rect 10045 25687 10103 25693
rect 10045 25684 10057 25687
rect 9732 25656 10057 25684
rect 9732 25644 9738 25656
rect 10045 25653 10057 25656
rect 10091 25653 10103 25687
rect 10045 25647 10103 25653
rect 11422 25644 11428 25696
rect 11480 25684 11486 25696
rect 13081 25687 13139 25693
rect 13081 25684 13093 25687
rect 11480 25656 13093 25684
rect 11480 25644 11486 25656
rect 13081 25653 13093 25656
rect 13127 25653 13139 25687
rect 13081 25647 13139 25653
rect 14369 25687 14427 25693
rect 14369 25653 14381 25687
rect 14415 25684 14427 25687
rect 14550 25684 14556 25696
rect 14415 25656 14556 25684
rect 14415 25653 14427 25656
rect 14369 25647 14427 25653
rect 14550 25644 14556 25656
rect 14608 25644 14614 25696
rect 20530 25684 20536 25696
rect 20491 25656 20536 25684
rect 20530 25644 20536 25656
rect 20588 25644 20594 25696
rect 22370 25644 22376 25696
rect 22428 25684 22434 25696
rect 22741 25687 22799 25693
rect 22741 25684 22753 25687
rect 22428 25656 22753 25684
rect 22428 25644 22434 25656
rect 22741 25653 22753 25656
rect 22787 25653 22799 25687
rect 22741 25647 22799 25653
rect 24762 25644 24768 25696
rect 24820 25684 24826 25696
rect 24820 25656 24865 25684
rect 24820 25644 24826 25656
rect 26602 25644 26608 25696
rect 26660 25684 26666 25696
rect 27154 25684 27160 25696
rect 26660 25656 27160 25684
rect 26660 25644 26666 25656
rect 27154 25644 27160 25656
rect 27212 25644 27218 25696
rect 31018 25644 31024 25696
rect 31076 25684 31082 25696
rect 31478 25684 31484 25696
rect 31076 25656 31484 25684
rect 31076 25644 31082 25656
rect 31478 25644 31484 25656
rect 31536 25644 31542 25696
rect 46474 25644 46480 25696
rect 46532 25684 46538 25696
rect 46845 25687 46903 25693
rect 46845 25684 46857 25687
rect 46532 25656 46857 25684
rect 46532 25644 46538 25656
rect 46845 25653 46857 25656
rect 46891 25653 46903 25687
rect 46845 25647 46903 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 14274 25480 14280 25492
rect 2746 25452 12434 25480
rect 14235 25452 14280 25480
rect 2314 25304 2320 25356
rect 2372 25344 2378 25356
rect 2746 25344 2774 25452
rect 10962 25372 10968 25424
rect 11020 25412 11026 25424
rect 12069 25415 12127 25421
rect 12069 25412 12081 25415
rect 11020 25384 12081 25412
rect 11020 25372 11026 25384
rect 12069 25381 12081 25384
rect 12115 25381 12127 25415
rect 12406 25412 12434 25452
rect 14274 25440 14280 25452
rect 14332 25440 14338 25492
rect 15105 25483 15163 25489
rect 15105 25449 15117 25483
rect 15151 25480 15163 25483
rect 15194 25480 15200 25492
rect 15151 25452 15200 25480
rect 15151 25449 15163 25452
rect 15105 25443 15163 25449
rect 15194 25440 15200 25452
rect 15252 25440 15258 25492
rect 15378 25440 15384 25492
rect 15436 25480 15442 25492
rect 15657 25483 15715 25489
rect 15657 25480 15669 25483
rect 15436 25452 15669 25480
rect 15436 25440 15442 25452
rect 15657 25449 15669 25452
rect 15703 25449 15715 25483
rect 25682 25480 25688 25492
rect 15657 25443 15715 25449
rect 19306 25452 25688 25480
rect 19306 25412 19334 25452
rect 25682 25440 25688 25452
rect 25740 25440 25746 25492
rect 27430 25440 27436 25492
rect 27488 25480 27494 25492
rect 28813 25483 28871 25489
rect 28813 25480 28825 25483
rect 27488 25452 28825 25480
rect 27488 25440 27494 25452
rect 28813 25449 28825 25452
rect 28859 25449 28871 25483
rect 31570 25480 31576 25492
rect 31531 25452 31576 25480
rect 28813 25443 28871 25449
rect 31570 25440 31576 25452
rect 31628 25440 31634 25492
rect 34238 25440 34244 25492
rect 34296 25480 34302 25492
rect 43346 25480 43352 25492
rect 34296 25452 43352 25480
rect 34296 25440 34302 25452
rect 43346 25440 43352 25452
rect 43404 25440 43410 25492
rect 12406 25384 19334 25412
rect 12069 25375 12127 25381
rect 23658 25372 23664 25424
rect 23716 25412 23722 25424
rect 23845 25415 23903 25421
rect 23845 25412 23857 25415
rect 23716 25384 23857 25412
rect 23716 25372 23722 25384
rect 23845 25381 23857 25384
rect 23891 25381 23903 25415
rect 23845 25375 23903 25381
rect 24397 25415 24455 25421
rect 24397 25381 24409 25415
rect 24443 25412 24455 25415
rect 24670 25412 24676 25424
rect 24443 25384 24676 25412
rect 24443 25381 24455 25384
rect 24397 25375 24455 25381
rect 24670 25372 24676 25384
rect 24728 25372 24734 25424
rect 26697 25415 26755 25421
rect 26697 25412 26709 25415
rect 25608 25384 26709 25412
rect 9674 25344 9680 25356
rect 2372 25316 2774 25344
rect 9635 25316 9680 25344
rect 2372 25304 2378 25316
rect 9674 25304 9680 25316
rect 9732 25304 9738 25356
rect 12342 25344 12348 25356
rect 11900 25316 12348 25344
rect 1854 25276 1860 25288
rect 1815 25248 1860 25276
rect 1854 25236 1860 25248
rect 1912 25236 1918 25288
rect 11900 25285 11928 25316
rect 12342 25304 12348 25316
rect 12400 25344 12406 25356
rect 20530 25344 20536 25356
rect 12400 25316 14964 25344
rect 12400 25304 12406 25316
rect 11885 25279 11943 25285
rect 11885 25245 11897 25279
rect 11931 25245 11943 25279
rect 12618 25276 12624 25288
rect 12531 25248 12624 25276
rect 11885 25239 11943 25245
rect 12618 25236 12624 25248
rect 12676 25276 12682 25288
rect 13262 25276 13268 25288
rect 12676 25248 13268 25276
rect 12676 25236 12682 25248
rect 13262 25236 13268 25248
rect 13320 25236 13326 25288
rect 13357 25279 13415 25285
rect 13357 25245 13369 25279
rect 13403 25276 13415 25279
rect 13446 25276 13452 25288
rect 13403 25248 13452 25276
rect 13403 25245 13415 25248
rect 13357 25239 13415 25245
rect 13446 25236 13452 25248
rect 13504 25236 13510 25288
rect 13538 25236 13544 25288
rect 13596 25276 13602 25288
rect 14936 25285 14964 25316
rect 15856 25316 20536 25344
rect 15856 25288 15884 25316
rect 20530 25304 20536 25316
rect 20588 25304 20594 25356
rect 22370 25344 22376 25356
rect 22331 25316 22376 25344
rect 22370 25304 22376 25316
rect 22428 25304 22434 25356
rect 24762 25344 24768 25356
rect 24596 25316 24768 25344
rect 14921 25279 14979 25285
rect 13596 25248 14872 25276
rect 13596 25236 13602 25248
rect 9950 25208 9956 25220
rect 9911 25180 9956 25208
rect 9950 25168 9956 25180
rect 10008 25168 10014 25220
rect 12713 25211 12771 25217
rect 12713 25208 12725 25211
rect 11178 25180 12725 25208
rect 12713 25177 12725 25180
rect 12759 25177 12771 25211
rect 12713 25171 12771 25177
rect 14093 25211 14151 25217
rect 14093 25177 14105 25211
rect 14139 25208 14151 25211
rect 14182 25208 14188 25220
rect 14139 25180 14188 25208
rect 14139 25177 14151 25180
rect 14093 25171 14151 25177
rect 14182 25168 14188 25180
rect 14240 25168 14246 25220
rect 14309 25211 14367 25217
rect 14309 25177 14321 25211
rect 14355 25208 14367 25211
rect 14734 25208 14740 25220
rect 14355 25180 14740 25208
rect 14355 25177 14367 25180
rect 14309 25171 14367 25177
rect 14734 25168 14740 25180
rect 14792 25168 14798 25220
rect 14844 25208 14872 25248
rect 14921 25245 14933 25279
rect 14967 25245 14979 25279
rect 15654 25276 15660 25288
rect 15615 25248 15660 25276
rect 14921 25239 14979 25245
rect 15654 25236 15660 25248
rect 15712 25236 15718 25288
rect 15838 25236 15844 25288
rect 15896 25276 15902 25288
rect 16485 25279 16543 25285
rect 15896 25248 15989 25276
rect 15896 25236 15902 25248
rect 16485 25245 16497 25279
rect 16531 25245 16543 25279
rect 17681 25279 17739 25285
rect 17681 25276 17693 25279
rect 16485 25239 16543 25245
rect 16684 25248 17693 25276
rect 16500 25208 16528 25239
rect 14844 25180 16528 25208
rect 16684 25152 16712 25248
rect 17681 25245 17693 25248
rect 17727 25245 17739 25279
rect 17681 25239 17739 25245
rect 22097 25279 22155 25285
rect 22097 25245 22109 25279
rect 22143 25245 22155 25279
rect 22097 25239 22155 25245
rect 22112 25208 22140 25239
rect 23474 25236 23480 25288
rect 23532 25236 23538 25288
rect 24596 25285 24624 25316
rect 24762 25304 24768 25316
rect 24820 25304 24826 25356
rect 24581 25279 24639 25285
rect 24581 25245 24593 25279
rect 24627 25245 24639 25279
rect 24581 25239 24639 25245
rect 24673 25279 24731 25285
rect 24673 25245 24685 25279
rect 24719 25276 24731 25279
rect 25038 25276 25044 25288
rect 24719 25248 25044 25276
rect 24719 25245 24731 25248
rect 24673 25239 24731 25245
rect 25038 25236 25044 25248
rect 25096 25236 25102 25288
rect 25608 25285 25636 25384
rect 26697 25381 26709 25384
rect 26743 25381 26755 25415
rect 34057 25415 34115 25421
rect 26697 25375 26755 25381
rect 27172 25384 30129 25412
rect 25774 25304 25780 25356
rect 25832 25344 25838 25356
rect 27172 25353 27200 25384
rect 27157 25347 27215 25353
rect 27157 25344 27169 25347
rect 25832 25316 27169 25344
rect 25832 25304 25838 25316
rect 27157 25313 27169 25316
rect 27203 25313 27215 25347
rect 27157 25307 27215 25313
rect 27341 25347 27399 25353
rect 27341 25313 27353 25347
rect 27387 25344 27399 25347
rect 28166 25344 28172 25356
rect 27387 25316 28172 25344
rect 27387 25313 27399 25316
rect 27341 25307 27399 25313
rect 28166 25304 28172 25316
rect 28224 25304 28230 25356
rect 30101 25344 30129 25384
rect 34057 25381 34069 25415
rect 34103 25412 34115 25415
rect 34606 25412 34612 25424
rect 34103 25384 34612 25412
rect 34103 25381 34115 25384
rect 34057 25375 34115 25381
rect 34606 25372 34612 25384
rect 34664 25372 34670 25424
rect 30929 25347 30987 25353
rect 30929 25344 30941 25347
rect 30101 25316 30941 25344
rect 25593 25279 25651 25285
rect 25593 25245 25605 25279
rect 25639 25245 25651 25279
rect 25593 25239 25651 25245
rect 25682 25236 25688 25288
rect 25740 25276 25746 25288
rect 25869 25279 25927 25285
rect 25869 25276 25881 25279
rect 25740 25248 25881 25276
rect 25740 25236 25746 25248
rect 25869 25245 25881 25248
rect 25915 25245 25927 25279
rect 25869 25239 25927 25245
rect 27065 25279 27123 25285
rect 27065 25245 27077 25279
rect 27111 25276 27123 25279
rect 28534 25276 28540 25288
rect 27111 25248 28540 25276
rect 27111 25245 27123 25248
rect 27065 25239 27123 25245
rect 28534 25236 28540 25248
rect 28592 25236 28598 25288
rect 28629 25279 28687 25285
rect 28629 25245 28641 25279
rect 28675 25276 28687 25279
rect 29270 25276 29276 25288
rect 28675 25248 29276 25276
rect 28675 25245 28687 25248
rect 28629 25239 28687 25245
rect 29270 25236 29276 25248
rect 29328 25236 29334 25288
rect 29638 25236 29644 25288
rect 29696 25254 29702 25288
rect 29817 25257 29875 25263
rect 29817 25254 29829 25257
rect 29696 25236 29829 25254
rect 29656 25226 29829 25236
rect 29817 25223 29829 25226
rect 29863 25223 29875 25257
rect 29914 25236 29920 25288
rect 29972 25276 29978 25288
rect 30101 25285 30129 25316
rect 30929 25313 30941 25316
rect 30975 25313 30987 25347
rect 30929 25307 30987 25313
rect 31202 25304 31208 25356
rect 31260 25344 31266 25356
rect 31481 25347 31539 25353
rect 31481 25344 31493 25347
rect 31260 25316 31493 25344
rect 31260 25304 31266 25316
rect 31481 25313 31493 25316
rect 31527 25313 31539 25347
rect 31481 25307 31539 25313
rect 33870 25304 33876 25356
rect 33928 25344 33934 25356
rect 34701 25347 34759 25353
rect 34701 25344 34713 25347
rect 33928 25316 34713 25344
rect 33928 25304 33934 25316
rect 34701 25313 34713 25316
rect 34747 25313 34759 25347
rect 46474 25344 46480 25356
rect 46435 25316 46480 25344
rect 34701 25307 34759 25313
rect 46474 25304 46480 25316
rect 46532 25304 46538 25356
rect 48130 25344 48136 25356
rect 48091 25316 48136 25344
rect 48130 25304 48136 25316
rect 48188 25304 48194 25356
rect 30060 25279 30129 25285
rect 29972 25248 30017 25276
rect 29972 25236 29978 25248
rect 30060 25245 30072 25279
rect 30106 25248 30129 25279
rect 30183 25279 30241 25285
rect 30106 25245 30118 25248
rect 30060 25239 30118 25245
rect 30183 25245 30195 25279
rect 30229 25276 30241 25279
rect 30282 25278 30288 25288
rect 30277 25276 30288 25278
rect 30229 25248 30288 25276
rect 30229 25245 30241 25248
rect 30183 25239 30241 25245
rect 30282 25236 30288 25248
rect 30340 25236 30346 25288
rect 31665 25279 31723 25285
rect 31665 25245 31677 25279
rect 31711 25276 31723 25279
rect 32490 25276 32496 25288
rect 31711 25248 32496 25276
rect 31711 25245 31723 25248
rect 31665 25239 31723 25245
rect 32490 25236 32496 25248
rect 32548 25236 32554 25288
rect 33778 25236 33784 25288
rect 33836 25276 33842 25288
rect 33965 25279 34023 25285
rect 33965 25276 33977 25279
rect 33836 25248 33977 25276
rect 33836 25236 33842 25248
rect 33965 25245 33977 25248
rect 34011 25245 34023 25279
rect 45462 25276 45468 25288
rect 45423 25248 45468 25276
rect 33965 25239 34023 25245
rect 45462 25236 45468 25248
rect 45520 25236 45526 25288
rect 46293 25279 46351 25285
rect 46293 25245 46305 25279
rect 46339 25245 46351 25279
rect 46293 25239 46351 25245
rect 22278 25208 22284 25220
rect 22112 25180 22284 25208
rect 22278 25168 22284 25180
rect 22336 25168 22342 25220
rect 24397 25211 24455 25217
rect 24397 25177 24409 25211
rect 24443 25177 24455 25211
rect 24397 25171 24455 25177
rect 1854 25100 1860 25152
rect 1912 25140 1918 25152
rect 1949 25143 2007 25149
rect 1949 25140 1961 25143
rect 1912 25112 1961 25140
rect 1912 25100 1918 25112
rect 1949 25109 1961 25112
rect 1995 25109 2007 25143
rect 1949 25103 2007 25109
rect 10870 25100 10876 25152
rect 10928 25140 10934 25152
rect 11425 25143 11483 25149
rect 11425 25140 11437 25143
rect 10928 25112 11437 25140
rect 10928 25100 10934 25112
rect 11425 25109 11437 25112
rect 11471 25109 11483 25143
rect 11425 25103 11483 25109
rect 13449 25143 13507 25149
rect 13449 25109 13461 25143
rect 13495 25140 13507 25143
rect 13630 25140 13636 25152
rect 13495 25112 13636 25140
rect 13495 25109 13507 25112
rect 13449 25103 13507 25109
rect 13630 25100 13636 25112
rect 13688 25100 13694 25152
rect 14458 25140 14464 25152
rect 14419 25112 14464 25140
rect 14458 25100 14464 25112
rect 14516 25100 14522 25152
rect 16666 25140 16672 25152
rect 16627 25112 16672 25140
rect 16666 25100 16672 25112
rect 16724 25100 16730 25152
rect 17773 25143 17831 25149
rect 17773 25109 17785 25143
rect 17819 25140 17831 25143
rect 17954 25140 17960 25152
rect 17819 25112 17960 25140
rect 17819 25109 17831 25112
rect 17773 25103 17831 25109
rect 17954 25100 17960 25112
rect 18012 25100 18018 25152
rect 21726 25100 21732 25152
rect 21784 25140 21790 25152
rect 24412 25140 24440 25171
rect 28810 25168 28816 25220
rect 28868 25208 28874 25220
rect 29362 25208 29368 25220
rect 28868 25180 29368 25208
rect 28868 25168 28874 25180
rect 29362 25168 29368 25180
rect 29420 25168 29426 25220
rect 29817 25217 29875 25223
rect 30650 25168 30656 25220
rect 30708 25208 30714 25220
rect 30745 25211 30803 25217
rect 30745 25208 30757 25211
rect 30708 25180 30757 25208
rect 30708 25168 30714 25180
rect 30745 25177 30757 25180
rect 30791 25177 30803 25211
rect 30745 25171 30803 25177
rect 31389 25211 31447 25217
rect 31389 25177 31401 25211
rect 31435 25208 31447 25211
rect 31570 25208 31576 25220
rect 31435 25180 31576 25208
rect 31435 25177 31447 25180
rect 31389 25171 31447 25177
rect 31570 25168 31576 25180
rect 31628 25168 31634 25220
rect 34698 25168 34704 25220
rect 34756 25208 34762 25220
rect 34977 25211 35035 25217
rect 34977 25208 34989 25211
rect 34756 25180 34989 25208
rect 34756 25168 34762 25180
rect 34977 25177 34989 25180
rect 35023 25177 35035 25211
rect 34977 25171 35035 25177
rect 35986 25168 35992 25220
rect 36044 25168 36050 25220
rect 46308 25208 46336 25239
rect 46474 25208 46480 25220
rect 46308 25180 46480 25208
rect 46474 25168 46480 25180
rect 46532 25168 46538 25220
rect 25406 25140 25412 25152
rect 21784 25112 24440 25140
rect 25367 25112 25412 25140
rect 21784 25100 21790 25112
rect 25406 25100 25412 25112
rect 25464 25100 25470 25152
rect 25777 25143 25835 25149
rect 25777 25109 25789 25143
rect 25823 25140 25835 25143
rect 25866 25140 25872 25152
rect 25823 25112 25872 25140
rect 25823 25109 25835 25112
rect 25777 25103 25835 25109
rect 25866 25100 25872 25112
rect 25924 25100 25930 25152
rect 29638 25140 29644 25152
rect 29599 25112 29644 25140
rect 29638 25100 29644 25112
rect 29696 25100 29702 25152
rect 31846 25140 31852 25152
rect 31807 25112 31852 25140
rect 31846 25100 31852 25112
rect 31904 25100 31910 25152
rect 32950 25100 32956 25152
rect 33008 25140 33014 25152
rect 36449 25143 36507 25149
rect 36449 25140 36461 25143
rect 33008 25112 36461 25140
rect 33008 25100 33014 25112
rect 36449 25109 36461 25112
rect 36495 25109 36507 25143
rect 36449 25103 36507 25109
rect 45554 25100 45560 25152
rect 45612 25140 45618 25152
rect 45612 25112 45657 25140
rect 45612 25100 45618 25112
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 24857 24939 24915 24945
rect 24857 24905 24869 24939
rect 24903 24936 24915 24939
rect 25866 24936 25872 24948
rect 24903 24908 25872 24936
rect 24903 24905 24915 24908
rect 24857 24899 24915 24905
rect 25866 24896 25872 24908
rect 25924 24896 25930 24948
rect 29914 24936 29920 24948
rect 29472 24908 29920 24936
rect 10870 24828 10876 24880
rect 10928 24868 10934 24880
rect 11517 24871 11575 24877
rect 11517 24868 11529 24871
rect 10928 24840 11529 24868
rect 10928 24828 10934 24840
rect 11517 24837 11529 24840
rect 11563 24837 11575 24871
rect 11717 24871 11775 24877
rect 11717 24868 11729 24871
rect 11517 24831 11575 24837
rect 11716 24837 11729 24868
rect 11763 24837 11775 24871
rect 13630 24868 13636 24880
rect 13591 24840 13636 24868
rect 11716 24831 11775 24837
rect 11716 24800 11744 24831
rect 13630 24828 13636 24840
rect 13688 24828 13694 24880
rect 17954 24828 17960 24880
rect 18012 24828 18018 24880
rect 21266 24868 21272 24880
rect 21227 24840 21272 24868
rect 21266 24828 21272 24840
rect 21324 24828 21330 24880
rect 25774 24828 25780 24880
rect 25832 24868 25838 24880
rect 26053 24871 26111 24877
rect 26053 24868 26065 24871
rect 25832 24840 26065 24868
rect 25832 24828 25838 24840
rect 26053 24837 26065 24840
rect 26099 24837 26111 24871
rect 26053 24831 26111 24837
rect 26142 24828 26148 24880
rect 26200 24868 26206 24880
rect 29472 24877 29500 24908
rect 29914 24896 29920 24908
rect 29972 24896 29978 24948
rect 30006 24896 30012 24948
rect 30064 24936 30070 24948
rect 30282 24936 30288 24948
rect 30064 24908 30288 24936
rect 30064 24896 30070 24908
rect 30282 24896 30288 24908
rect 30340 24896 30346 24948
rect 32950 24936 32956 24948
rect 30392 24908 32956 24936
rect 29457 24871 29515 24877
rect 29457 24868 29469 24871
rect 26200 24840 29469 24868
rect 26200 24828 26206 24840
rect 12437 24803 12495 24809
rect 11716 24772 11836 24800
rect 11808 24744 11836 24772
rect 12437 24769 12449 24803
rect 12483 24769 12495 24803
rect 23014 24800 23020 24812
rect 22975 24772 23020 24800
rect 12437 24763 12495 24769
rect 8386 24732 8392 24744
rect 8347 24704 8392 24732
rect 8386 24692 8392 24704
rect 8444 24692 8450 24744
rect 8573 24735 8631 24741
rect 8573 24701 8585 24735
rect 8619 24732 8631 24735
rect 8754 24732 8760 24744
rect 8619 24704 8760 24732
rect 8619 24701 8631 24704
rect 8573 24695 8631 24701
rect 8754 24692 8760 24704
rect 8812 24692 8818 24744
rect 8849 24735 8907 24741
rect 8849 24701 8861 24735
rect 8895 24701 8907 24735
rect 8849 24695 8907 24701
rect 3602 24556 3608 24608
rect 3660 24596 3666 24608
rect 8864 24596 8892 24695
rect 11790 24692 11796 24744
rect 11848 24692 11854 24744
rect 11422 24624 11428 24676
rect 11480 24664 11486 24676
rect 11885 24667 11943 24673
rect 11885 24664 11897 24667
rect 11480 24636 11897 24664
rect 11480 24624 11486 24636
rect 11885 24633 11897 24636
rect 11931 24633 11943 24667
rect 12452 24664 12480 24763
rect 23014 24760 23020 24772
rect 23072 24760 23078 24812
rect 23109 24803 23167 24809
rect 23109 24769 23121 24803
rect 23155 24800 23167 24803
rect 23474 24800 23480 24812
rect 23155 24772 23480 24800
rect 23155 24769 23167 24772
rect 23109 24763 23167 24769
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 24670 24800 24676 24812
rect 24631 24772 24676 24800
rect 24670 24760 24676 24772
rect 24728 24760 24734 24812
rect 24946 24760 24952 24812
rect 25004 24800 25010 24812
rect 25004 24772 25049 24800
rect 25004 24760 25010 24772
rect 25682 24760 25688 24812
rect 25740 24800 25746 24812
rect 25869 24803 25927 24809
rect 25869 24800 25881 24803
rect 25740 24772 25881 24800
rect 25740 24760 25746 24772
rect 25869 24769 25881 24772
rect 25915 24769 25927 24803
rect 25869 24763 25927 24769
rect 26237 24803 26295 24809
rect 26237 24769 26249 24803
rect 26283 24800 26295 24803
rect 26418 24800 26424 24812
rect 26283 24772 26424 24800
rect 26283 24769 26295 24772
rect 26237 24763 26295 24769
rect 26418 24760 26424 24772
rect 26476 24760 26482 24812
rect 26988 24809 27016 24840
rect 29457 24837 29469 24840
rect 29503 24837 29515 24871
rect 29457 24831 29515 24837
rect 29638 24828 29644 24880
rect 29696 24868 29702 24880
rect 29696 24840 30328 24868
rect 29696 24828 29702 24840
rect 26973 24803 27031 24809
rect 26973 24769 26985 24803
rect 27019 24769 27031 24803
rect 27982 24800 27988 24812
rect 27943 24772 27988 24800
rect 26973 24763 27031 24769
rect 27982 24760 27988 24772
rect 28040 24760 28046 24812
rect 28169 24803 28227 24809
rect 28169 24769 28181 24803
rect 28215 24800 28227 24803
rect 28534 24800 28540 24812
rect 28215 24772 28540 24800
rect 28215 24769 28227 24772
rect 28169 24763 28227 24769
rect 28534 24760 28540 24772
rect 28592 24800 28598 24812
rect 28592 24772 28994 24800
rect 28592 24760 28598 24772
rect 13449 24735 13507 24741
rect 13449 24701 13461 24735
rect 13495 24732 13507 24735
rect 14366 24732 14372 24744
rect 13495 24704 14372 24732
rect 13495 24701 13507 24704
rect 13449 24695 13507 24701
rect 14366 24692 14372 24704
rect 14424 24692 14430 24744
rect 14550 24732 14556 24744
rect 14511 24704 14556 24732
rect 14550 24692 14556 24704
rect 14608 24692 14614 24744
rect 17034 24692 17040 24744
rect 17092 24732 17098 24744
rect 17221 24735 17279 24741
rect 17221 24732 17233 24735
rect 17092 24704 17233 24732
rect 17092 24692 17098 24704
rect 17221 24701 17233 24704
rect 17267 24701 17279 24735
rect 17221 24695 17279 24701
rect 17497 24735 17555 24741
rect 17497 24701 17509 24735
rect 17543 24732 17555 24735
rect 18046 24732 18052 24744
rect 17543 24704 18052 24732
rect 17543 24701 17555 24704
rect 17497 24695 17555 24701
rect 18046 24692 18052 24704
rect 18104 24692 18110 24744
rect 18966 24732 18972 24744
rect 18879 24704 18972 24732
rect 18966 24692 18972 24704
rect 19024 24732 19030 24744
rect 19429 24735 19487 24741
rect 19429 24732 19441 24735
rect 19024 24704 19441 24732
rect 19024 24692 19030 24704
rect 19429 24701 19441 24704
rect 19475 24701 19487 24735
rect 19610 24732 19616 24744
rect 19571 24704 19616 24732
rect 19429 24695 19487 24701
rect 19610 24692 19616 24704
rect 19668 24692 19674 24744
rect 28258 24692 28264 24744
rect 28316 24732 28322 24744
rect 28445 24735 28503 24741
rect 28445 24732 28457 24735
rect 28316 24704 28457 24732
rect 28316 24692 28322 24704
rect 28445 24701 28457 24704
rect 28491 24701 28503 24735
rect 28966 24732 28994 24772
rect 29270 24760 29276 24812
rect 29328 24800 29334 24812
rect 29914 24800 29920 24812
rect 29328 24772 29920 24800
rect 29328 24760 29334 24772
rect 29914 24760 29920 24772
rect 29972 24760 29978 24812
rect 30300 24809 30328 24840
rect 30285 24803 30343 24809
rect 30285 24769 30297 24803
rect 30331 24769 30343 24803
rect 30285 24763 30343 24769
rect 30392 24732 30420 24908
rect 32950 24896 32956 24908
rect 33008 24896 33014 24948
rect 30558 24828 30564 24880
rect 30616 24868 30622 24880
rect 31202 24868 31208 24880
rect 30616 24840 31208 24868
rect 30616 24828 30622 24840
rect 31202 24828 31208 24840
rect 31260 24828 31266 24880
rect 35710 24868 35716 24880
rect 35623 24840 35716 24868
rect 35710 24828 35716 24840
rect 35768 24868 35774 24880
rect 45462 24868 45468 24880
rect 35768 24840 36124 24868
rect 35768 24828 35774 24840
rect 31021 24803 31079 24809
rect 31021 24769 31033 24803
rect 31067 24800 31079 24803
rect 31294 24800 31300 24812
rect 31067 24772 31300 24800
rect 31067 24769 31079 24772
rect 31021 24763 31079 24769
rect 31294 24760 31300 24772
rect 31352 24760 31358 24812
rect 33778 24760 33784 24812
rect 33836 24800 33842 24812
rect 34701 24803 34759 24809
rect 34701 24800 34713 24803
rect 33836 24772 34713 24800
rect 33836 24760 33842 24772
rect 34701 24769 34713 24772
rect 34747 24769 34759 24803
rect 34701 24763 34759 24769
rect 34793 24803 34851 24809
rect 34793 24769 34805 24803
rect 34839 24800 34851 24803
rect 35986 24800 35992 24812
rect 34839 24772 35992 24800
rect 34839 24769 34851 24772
rect 34793 24763 34851 24769
rect 35986 24760 35992 24772
rect 36044 24760 36050 24812
rect 36096 24809 36124 24840
rect 40052 24840 41460 24868
rect 36081 24803 36139 24809
rect 36081 24769 36093 24803
rect 36127 24800 36139 24803
rect 40052 24800 40080 24840
rect 36127 24772 40080 24800
rect 36127 24769 36139 24772
rect 36081 24763 36139 24769
rect 30558 24732 30564 24744
rect 28966 24704 30420 24732
rect 30519 24704 30564 24732
rect 28445 24695 28503 24701
rect 30558 24692 30564 24704
rect 30616 24692 30622 24744
rect 40034 24732 40040 24744
rect 30852 24704 36032 24732
rect 39995 24704 40040 24732
rect 12618 24664 12624 24676
rect 12452 24636 12624 24664
rect 11885 24627 11943 24633
rect 12618 24624 12624 24636
rect 12676 24664 12682 24676
rect 14458 24664 14464 24676
rect 12676 24636 14464 24664
rect 12676 24624 12682 24636
rect 14458 24624 14464 24636
rect 14516 24624 14522 24676
rect 25866 24624 25872 24676
rect 25924 24664 25930 24676
rect 27157 24667 27215 24673
rect 27157 24664 27169 24667
rect 25924 24636 27169 24664
rect 25924 24624 25930 24636
rect 27157 24633 27169 24636
rect 27203 24633 27215 24667
rect 27157 24627 27215 24633
rect 27890 24624 27896 24676
rect 27948 24664 27954 24676
rect 27948 24636 30696 24664
rect 27948 24624 27954 24636
rect 3660 24568 8892 24596
rect 3660 24556 3666 24568
rect 11606 24556 11612 24608
rect 11664 24596 11670 24608
rect 11701 24599 11759 24605
rect 11701 24596 11713 24599
rect 11664 24568 11713 24596
rect 11664 24556 11670 24568
rect 11701 24565 11713 24568
rect 11747 24565 11759 24599
rect 11701 24559 11759 24565
rect 11974 24556 11980 24608
rect 12032 24596 12038 24608
rect 12529 24599 12587 24605
rect 12529 24596 12541 24599
rect 12032 24568 12541 24596
rect 12032 24556 12038 24568
rect 12529 24565 12541 24568
rect 12575 24565 12587 24599
rect 12529 24559 12587 24565
rect 23014 24556 23020 24608
rect 23072 24596 23078 24608
rect 24489 24599 24547 24605
rect 24489 24596 24501 24599
rect 23072 24568 24501 24596
rect 23072 24556 23078 24568
rect 24489 24565 24501 24568
rect 24535 24565 24547 24599
rect 24489 24559 24547 24565
rect 25958 24556 25964 24608
rect 26016 24596 26022 24608
rect 26421 24599 26479 24605
rect 26421 24596 26433 24599
rect 26016 24568 26433 24596
rect 26016 24556 26022 24568
rect 26421 24565 26433 24568
rect 26467 24565 26479 24599
rect 26421 24559 26479 24565
rect 28074 24556 28080 24608
rect 28132 24596 28138 24608
rect 28353 24599 28411 24605
rect 28353 24596 28365 24599
rect 28132 24568 28365 24596
rect 28132 24556 28138 24568
rect 28353 24565 28365 24568
rect 28399 24565 28411 24599
rect 28353 24559 28411 24565
rect 30101 24599 30159 24605
rect 30101 24565 30113 24599
rect 30147 24596 30159 24599
rect 30374 24596 30380 24608
rect 30147 24568 30380 24596
rect 30147 24565 30159 24568
rect 30101 24559 30159 24565
rect 30374 24556 30380 24568
rect 30432 24556 30438 24608
rect 30466 24556 30472 24608
rect 30524 24596 30530 24608
rect 30668 24596 30696 24636
rect 30852 24596 30880 24704
rect 33042 24624 33048 24676
rect 33100 24664 33106 24676
rect 35710 24664 35716 24676
rect 33100 24636 35716 24664
rect 33100 24624 33106 24636
rect 35710 24624 35716 24636
rect 35768 24624 35774 24676
rect 36004 24664 36032 24704
rect 40034 24692 40040 24704
rect 40092 24692 40098 24744
rect 40221 24735 40279 24741
rect 40221 24701 40233 24735
rect 40267 24732 40279 24735
rect 40310 24732 40316 24744
rect 40267 24704 40316 24732
rect 40267 24701 40279 24704
rect 40221 24695 40279 24701
rect 40310 24692 40316 24704
rect 40368 24692 40374 24744
rect 40402 24692 40408 24744
rect 40460 24732 40466 24744
rect 40497 24735 40555 24741
rect 40497 24732 40509 24735
rect 40460 24704 40509 24732
rect 40460 24692 40466 24704
rect 40497 24701 40509 24704
rect 40543 24701 40555 24735
rect 41432 24732 41460 24840
rect 44192 24840 45468 24868
rect 42886 24760 42892 24812
rect 42944 24800 42950 24812
rect 43441 24803 43499 24809
rect 43441 24800 43453 24803
rect 42944 24772 43453 24800
rect 42944 24760 42950 24772
rect 43441 24769 43453 24772
rect 43487 24769 43499 24803
rect 43622 24800 43628 24812
rect 43583 24772 43628 24800
rect 43441 24763 43499 24769
rect 43622 24760 43628 24772
rect 43680 24760 43686 24812
rect 44192 24732 44220 24840
rect 45462 24828 45468 24840
rect 45520 24828 45526 24880
rect 46768 24840 46980 24868
rect 44542 24760 44548 24812
rect 44600 24800 44606 24812
rect 44637 24803 44695 24809
rect 44637 24800 44649 24803
rect 44600 24772 44649 24800
rect 44600 24760 44606 24772
rect 44637 24769 44649 24772
rect 44683 24769 44695 24803
rect 44637 24763 44695 24769
rect 45281 24803 45339 24809
rect 45281 24769 45293 24803
rect 45327 24800 45339 24803
rect 45554 24800 45560 24812
rect 45327 24772 45560 24800
rect 45327 24769 45339 24772
rect 45281 24763 45339 24769
rect 45554 24760 45560 24772
rect 45612 24760 45618 24812
rect 41432 24704 44220 24732
rect 40497 24695 40555 24701
rect 44266 24692 44272 24744
rect 44324 24732 44330 24744
rect 46768 24732 46796 24840
rect 46842 24760 46848 24812
rect 46900 24760 46906 24812
rect 46952 24800 46980 24840
rect 47118 24800 47124 24812
rect 46952 24772 47124 24800
rect 47118 24760 47124 24772
rect 47176 24800 47182 24812
rect 47581 24803 47639 24809
rect 47581 24800 47593 24803
rect 47176 24772 47593 24800
rect 47176 24760 47182 24772
rect 47581 24769 47593 24772
rect 47627 24769 47639 24803
rect 47581 24763 47639 24769
rect 44324 24704 46796 24732
rect 46860 24732 46888 24760
rect 47673 24735 47731 24741
rect 47673 24732 47685 24735
rect 46860 24704 47685 24732
rect 44324 24692 44330 24704
rect 47673 24701 47685 24704
rect 47719 24701 47731 24735
rect 47673 24695 47731 24701
rect 46842 24664 46848 24676
rect 36004 24636 46848 24664
rect 46842 24624 46848 24636
rect 46900 24624 46906 24676
rect 31386 24596 31392 24608
rect 30524 24568 30569 24596
rect 30668 24568 30880 24596
rect 31347 24568 31392 24596
rect 30524 24556 30530 24568
rect 31386 24556 31392 24568
rect 31444 24556 31450 24608
rect 36354 24596 36360 24608
rect 36315 24568 36360 24596
rect 36354 24556 36360 24568
rect 36412 24556 36418 24608
rect 43533 24599 43591 24605
rect 43533 24565 43545 24599
rect 43579 24596 43591 24599
rect 43898 24596 43904 24608
rect 43579 24568 43904 24596
rect 43579 24565 43591 24568
rect 43533 24559 43591 24565
rect 43898 24556 43904 24568
rect 43956 24556 43962 24608
rect 44729 24599 44787 24605
rect 44729 24565 44741 24599
rect 44775 24596 44787 24599
rect 46382 24596 46388 24608
rect 44775 24568 46388 24596
rect 44775 24565 44787 24568
rect 44729 24559 44787 24565
rect 46382 24556 46388 24568
rect 46440 24556 46446 24608
rect 46566 24596 46572 24608
rect 46527 24568 46572 24596
rect 46566 24556 46572 24568
rect 46624 24556 46630 24608
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 9950 24352 9956 24404
rect 10008 24392 10014 24404
rect 10321 24395 10379 24401
rect 10321 24392 10333 24395
rect 10008 24364 10333 24392
rect 10008 24352 10014 24364
rect 10321 24361 10333 24364
rect 10367 24361 10379 24395
rect 10321 24355 10379 24361
rect 11790 24352 11796 24404
rect 11848 24392 11854 24404
rect 12529 24395 12587 24401
rect 12529 24392 12541 24395
rect 11848 24364 12541 24392
rect 11848 24352 11854 24364
rect 12529 24361 12541 24364
rect 12575 24361 12587 24395
rect 17034 24392 17040 24404
rect 16995 24364 17040 24392
rect 12529 24355 12587 24361
rect 17034 24352 17040 24364
rect 17092 24352 17098 24404
rect 18509 24395 18567 24401
rect 18509 24392 18521 24395
rect 17788 24364 18521 24392
rect 12713 24327 12771 24333
rect 12713 24324 12725 24327
rect 12406 24296 12725 24324
rect 12406 24268 12434 24296
rect 12713 24293 12725 24296
rect 12759 24293 12771 24327
rect 15838 24324 15844 24336
rect 12713 24287 12771 24293
rect 14844 24296 15844 24324
rect 8386 24216 8392 24268
rect 8444 24256 8450 24268
rect 10870 24256 10876 24268
rect 8444 24228 10876 24256
rect 8444 24216 8450 24228
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 10965 24259 11023 24265
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 12406 24256 12440 24268
rect 11011 24228 12440 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 12434 24216 12440 24228
rect 12492 24216 12498 24268
rect 14844 24265 14872 24296
rect 15838 24284 15844 24296
rect 15896 24284 15902 24336
rect 14829 24259 14887 24265
rect 14829 24225 14841 24259
rect 14875 24225 14887 24259
rect 14829 24219 14887 24225
rect 15105 24259 15163 24265
rect 15105 24225 15117 24259
rect 15151 24256 15163 24259
rect 15378 24256 15384 24268
rect 15151 24228 15384 24256
rect 15151 24225 15163 24228
rect 15105 24219 15163 24225
rect 15378 24216 15384 24228
rect 15436 24216 15442 24268
rect 10502 24191 10560 24197
rect 10502 24157 10514 24191
rect 10548 24188 10560 24191
rect 11422 24188 11428 24200
rect 10548 24160 11428 24188
rect 10548 24157 10560 24160
rect 10502 24151 10560 24157
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 11606 24188 11612 24200
rect 11567 24160 11612 24188
rect 11606 24148 11612 24160
rect 11664 24148 11670 24200
rect 11882 24188 11888 24200
rect 11843 24160 11888 24188
rect 11882 24148 11888 24160
rect 11940 24148 11946 24200
rect 13078 24188 13084 24200
rect 12176 24160 13084 24188
rect 11624 24120 11652 24148
rect 12176 24120 12204 24160
rect 13078 24148 13084 24160
rect 13136 24148 13142 24200
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24188 13231 24191
rect 13538 24188 13544 24200
rect 13219 24160 13544 24188
rect 13219 24157 13231 24160
rect 13173 24151 13231 24157
rect 13538 24148 13544 24160
rect 13596 24148 13602 24200
rect 13630 24148 13636 24200
rect 13688 24188 13694 24200
rect 14737 24191 14795 24197
rect 14737 24188 14749 24191
rect 13688 24160 14749 24188
rect 13688 24148 13694 24160
rect 14737 24157 14749 24160
rect 14783 24157 14795 24191
rect 14737 24151 14795 24157
rect 15749 24191 15807 24197
rect 15749 24157 15761 24191
rect 15795 24188 15807 24191
rect 16850 24188 16856 24200
rect 15795 24160 16856 24188
rect 15795 24157 15807 24160
rect 15749 24151 15807 24157
rect 12618 24129 12624 24132
rect 12345 24123 12403 24129
rect 12345 24120 12357 24123
rect 11624 24092 12357 24120
rect 12345 24089 12357 24092
rect 12391 24089 12403 24123
rect 12345 24083 12403 24089
rect 12561 24123 12624 24129
rect 12561 24089 12573 24123
rect 12607 24089 12624 24123
rect 12561 24083 12624 24089
rect 12618 24080 12624 24083
rect 12676 24080 12682 24132
rect 14752 24120 14780 24151
rect 16850 24148 16856 24160
rect 16908 24188 16914 24200
rect 17788 24197 17816 24364
rect 18509 24361 18521 24364
rect 18555 24392 18567 24395
rect 19058 24392 19064 24404
rect 18555 24364 19064 24392
rect 18555 24361 18567 24364
rect 18509 24355 18567 24361
rect 19058 24352 19064 24364
rect 19116 24352 19122 24404
rect 19429 24395 19487 24401
rect 19429 24361 19441 24395
rect 19475 24392 19487 24395
rect 19610 24392 19616 24404
rect 19475 24364 19616 24392
rect 19475 24361 19487 24364
rect 19429 24355 19487 24361
rect 19610 24352 19616 24364
rect 19668 24352 19674 24404
rect 26970 24352 26976 24404
rect 27028 24392 27034 24404
rect 28169 24395 28227 24401
rect 28169 24392 28181 24395
rect 27028 24364 28181 24392
rect 27028 24352 27034 24364
rect 28169 24361 28181 24364
rect 28215 24392 28227 24395
rect 28258 24392 28264 24404
rect 28215 24364 28264 24392
rect 28215 24361 28227 24364
rect 28169 24355 28227 24361
rect 28258 24352 28264 24364
rect 28316 24352 28322 24404
rect 28442 24352 28448 24404
rect 28500 24392 28506 24404
rect 28626 24392 28632 24404
rect 28500 24364 28632 24392
rect 28500 24352 28506 24364
rect 28626 24352 28632 24364
rect 28684 24352 28690 24404
rect 30190 24392 30196 24404
rect 30151 24364 30196 24392
rect 30190 24352 30196 24364
rect 30248 24352 30254 24404
rect 30466 24392 30472 24404
rect 30300 24364 30472 24392
rect 18138 24284 18144 24336
rect 18196 24324 18202 24336
rect 18693 24327 18751 24333
rect 18693 24324 18705 24327
rect 18196 24296 18705 24324
rect 18196 24284 18202 24296
rect 18693 24293 18705 24296
rect 18739 24293 18751 24327
rect 27249 24327 27307 24333
rect 27249 24324 27261 24327
rect 18693 24287 18751 24293
rect 26252 24296 27261 24324
rect 18782 24216 18788 24268
rect 18840 24256 18846 24268
rect 19981 24259 20039 24265
rect 19981 24256 19993 24259
rect 18840 24228 19993 24256
rect 18840 24216 18846 24228
rect 19981 24225 19993 24228
rect 20027 24225 20039 24259
rect 19981 24219 20039 24225
rect 25498 24216 25504 24268
rect 25556 24256 25562 24268
rect 25556 24228 26188 24256
rect 25556 24216 25562 24228
rect 16945 24191 17003 24197
rect 16945 24188 16957 24191
rect 16908 24160 16957 24188
rect 16908 24148 16914 24160
rect 16945 24157 16957 24160
rect 16991 24157 17003 24191
rect 17773 24191 17831 24197
rect 17773 24188 17785 24191
rect 16945 24151 17003 24157
rect 17052 24160 17785 24188
rect 16574 24120 16580 24132
rect 14752 24092 16580 24120
rect 16574 24080 16580 24092
rect 16632 24120 16638 24132
rect 17052 24120 17080 24160
rect 17773 24157 17785 24160
rect 17819 24157 17831 24191
rect 17773 24151 17831 24157
rect 17865 24191 17923 24197
rect 17865 24157 17877 24191
rect 17911 24188 17923 24191
rect 19337 24191 19395 24197
rect 17911 24160 19104 24188
rect 17911 24157 17923 24160
rect 17865 24151 17923 24157
rect 16632 24092 17080 24120
rect 17589 24123 17647 24129
rect 16632 24080 16638 24092
rect 17589 24089 17601 24123
rect 17635 24120 17647 24123
rect 18325 24123 18383 24129
rect 18325 24120 18337 24123
rect 17635 24092 18337 24120
rect 17635 24089 17647 24092
rect 17589 24083 17647 24089
rect 18325 24089 18337 24092
rect 18371 24120 18383 24123
rect 18966 24120 18972 24132
rect 18371 24092 18972 24120
rect 18371 24089 18383 24092
rect 18325 24083 18383 24089
rect 18966 24080 18972 24092
rect 19024 24080 19030 24132
rect 10505 24055 10563 24061
rect 10505 24021 10517 24055
rect 10551 24052 10563 24055
rect 11054 24052 11060 24064
rect 10551 24024 11060 24052
rect 10551 24021 10563 24024
rect 10505 24015 10563 24021
rect 11054 24012 11060 24024
rect 11112 24012 11118 24064
rect 11422 24052 11428 24064
rect 11383 24024 11428 24052
rect 11422 24012 11428 24024
rect 11480 24012 11486 24064
rect 11790 24052 11796 24064
rect 11751 24024 11796 24052
rect 11790 24012 11796 24024
rect 11848 24012 11854 24064
rect 13354 24052 13360 24064
rect 13315 24024 13360 24052
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 15194 24012 15200 24064
rect 15252 24052 15258 24064
rect 15749 24055 15807 24061
rect 15749 24052 15761 24055
rect 15252 24024 15761 24052
rect 15252 24012 15258 24024
rect 15749 24021 15761 24024
rect 15795 24021 15807 24055
rect 17678 24052 17684 24064
rect 17736 24061 17742 24064
rect 17645 24024 17684 24052
rect 15749 24015 15807 24021
rect 17678 24012 17684 24024
rect 17736 24015 17745 24061
rect 18535 24055 18593 24061
rect 18535 24021 18547 24055
rect 18581 24052 18593 24055
rect 19076 24052 19104 24160
rect 19337 24157 19349 24191
rect 19383 24188 19395 24191
rect 19886 24188 19892 24200
rect 19383 24160 19892 24188
rect 19383 24157 19395 24160
rect 19337 24151 19395 24157
rect 19886 24148 19892 24160
rect 19944 24148 19950 24200
rect 23106 24148 23112 24200
rect 23164 24188 23170 24200
rect 23385 24191 23443 24197
rect 23385 24188 23397 24191
rect 23164 24160 23397 24188
rect 23164 24148 23170 24160
rect 23385 24157 23397 24160
rect 23431 24157 23443 24191
rect 25958 24188 25964 24200
rect 25919 24160 25964 24188
rect 23385 24151 23443 24157
rect 25958 24148 25964 24160
rect 26016 24148 26022 24200
rect 26160 24197 26188 24228
rect 26252 24197 26280 24296
rect 27249 24293 27261 24296
rect 27295 24293 27307 24327
rect 27249 24287 27307 24293
rect 29546 24284 29552 24336
rect 29604 24324 29610 24336
rect 30300 24324 30328 24364
rect 30466 24352 30472 24364
rect 30524 24352 30530 24404
rect 30558 24352 30564 24404
rect 30616 24392 30622 24404
rect 33229 24395 33287 24401
rect 33229 24392 33241 24395
rect 30616 24364 33241 24392
rect 30616 24352 30622 24364
rect 33229 24361 33241 24364
rect 33275 24361 33287 24395
rect 33229 24355 33287 24361
rect 36262 24352 36268 24404
rect 36320 24392 36326 24404
rect 44266 24392 44272 24404
rect 36320 24364 44272 24392
rect 36320 24352 36326 24364
rect 44266 24352 44272 24364
rect 44324 24352 44330 24404
rect 29604 24296 30328 24324
rect 29604 24284 29610 24296
rect 30374 24284 30380 24336
rect 30432 24324 30438 24336
rect 30432 24296 30972 24324
rect 30432 24284 30438 24296
rect 26973 24259 27031 24265
rect 26973 24225 26985 24259
rect 27019 24256 27031 24259
rect 28074 24256 28080 24268
rect 27019 24228 28080 24256
rect 27019 24225 27031 24228
rect 26973 24219 27031 24225
rect 28074 24216 28080 24228
rect 28132 24216 28138 24268
rect 29641 24259 29699 24265
rect 29641 24225 29653 24259
rect 29687 24256 29699 24259
rect 30944 24256 30972 24296
rect 40034 24284 40040 24336
rect 40092 24324 40098 24336
rect 40862 24324 40868 24336
rect 40092 24296 40868 24324
rect 40092 24284 40098 24296
rect 40862 24284 40868 24296
rect 40920 24324 40926 24336
rect 41509 24327 41567 24333
rect 41509 24324 41521 24327
rect 40920 24296 41521 24324
rect 40920 24284 40926 24296
rect 41509 24293 41521 24296
rect 41555 24293 41567 24327
rect 41509 24287 41567 24293
rect 45922 24284 45928 24336
rect 45980 24324 45986 24336
rect 45980 24296 46704 24324
rect 45980 24284 45986 24296
rect 31757 24259 31815 24265
rect 31757 24256 31769 24259
rect 29687 24228 30512 24256
rect 30944 24228 31769 24256
rect 29687 24225 29699 24228
rect 29641 24219 29699 24225
rect 26145 24191 26203 24197
rect 26145 24157 26157 24191
rect 26191 24157 26203 24191
rect 26145 24151 26203 24157
rect 26237 24191 26295 24197
rect 26237 24157 26249 24191
rect 26283 24157 26295 24191
rect 26237 24151 26295 24157
rect 26881 24191 26939 24197
rect 26881 24157 26893 24191
rect 26927 24157 26939 24191
rect 28166 24188 28172 24200
rect 28127 24160 28172 24188
rect 26881 24151 26939 24157
rect 20162 24120 20168 24132
rect 20123 24092 20168 24120
rect 20162 24080 20168 24092
rect 20220 24080 20226 24132
rect 21818 24120 21824 24132
rect 21779 24092 21824 24120
rect 21818 24080 21824 24092
rect 21876 24080 21882 24132
rect 25682 24080 25688 24132
rect 25740 24120 25746 24132
rect 26896 24120 26924 24151
rect 28166 24148 28172 24160
rect 28224 24148 28230 24200
rect 28353 24191 28411 24197
rect 28353 24157 28365 24191
rect 28399 24157 28411 24191
rect 28353 24151 28411 24157
rect 28445 24191 28503 24197
rect 28445 24157 28457 24191
rect 28491 24188 28503 24191
rect 28534 24188 28540 24200
rect 28491 24160 28540 24188
rect 28491 24157 28503 24160
rect 28445 24151 28503 24157
rect 26970 24120 26976 24132
rect 25740 24092 26976 24120
rect 25740 24080 25746 24092
rect 26970 24080 26976 24092
rect 27028 24080 27034 24132
rect 28368 24120 28396 24151
rect 28534 24148 28540 24160
rect 28592 24148 28598 24200
rect 29546 24188 29552 24200
rect 29507 24160 29552 24188
rect 29546 24148 29552 24160
rect 29604 24148 29610 24200
rect 29733 24191 29791 24197
rect 29733 24157 29745 24191
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 28368 24092 28488 24120
rect 28460 24064 28488 24092
rect 20530 24052 20536 24064
rect 18581 24024 20536 24052
rect 18581 24021 18593 24024
rect 18535 24015 18593 24021
rect 17736 24012 17742 24015
rect 20530 24012 20536 24024
rect 20588 24012 20594 24064
rect 23474 24052 23480 24064
rect 23435 24024 23480 24052
rect 23474 24012 23480 24024
rect 23532 24012 23538 24064
rect 25498 24012 25504 24064
rect 25556 24052 25562 24064
rect 25777 24055 25835 24061
rect 25777 24052 25789 24055
rect 25556 24024 25789 24052
rect 25556 24012 25562 24024
rect 25777 24021 25789 24024
rect 25823 24021 25835 24055
rect 25777 24015 25835 24021
rect 28442 24012 28448 24064
rect 28500 24012 28506 24064
rect 29748 24052 29776 24151
rect 29914 24148 29920 24200
rect 29972 24188 29978 24200
rect 30190 24188 30196 24200
rect 29972 24160 30196 24188
rect 29972 24148 29978 24160
rect 30190 24148 30196 24160
rect 30248 24148 30254 24200
rect 30484 24197 30512 24228
rect 31757 24225 31769 24228
rect 31803 24225 31815 24259
rect 37090 24256 37096 24268
rect 37051 24228 37096 24256
rect 31757 24219 31815 24225
rect 37090 24216 37096 24228
rect 37148 24256 37154 24268
rect 37148 24228 40908 24256
rect 37148 24216 37154 24228
rect 30469 24191 30527 24197
rect 30469 24157 30481 24191
rect 30515 24157 30527 24191
rect 31478 24188 31484 24200
rect 31439 24160 31484 24188
rect 30469 24151 30527 24157
rect 31478 24148 31484 24160
rect 31536 24148 31542 24200
rect 32858 24148 32864 24200
rect 32916 24148 32922 24200
rect 35529 24191 35587 24197
rect 35529 24157 35541 24191
rect 35575 24188 35587 24191
rect 36354 24188 36360 24200
rect 35575 24160 36360 24188
rect 35575 24157 35587 24160
rect 35529 24151 35587 24157
rect 36354 24148 36360 24160
rect 36412 24148 36418 24200
rect 38746 24148 38752 24200
rect 38804 24188 38810 24200
rect 40221 24191 40279 24197
rect 40221 24188 40233 24191
rect 38804 24160 40233 24188
rect 38804 24148 38810 24160
rect 40221 24157 40233 24160
rect 40267 24157 40279 24191
rect 40221 24151 40279 24157
rect 30377 24123 30435 24129
rect 30377 24089 30389 24123
rect 30423 24120 30435 24123
rect 31386 24120 31392 24132
rect 30423 24092 31392 24120
rect 30423 24089 30435 24092
rect 30377 24083 30435 24089
rect 31386 24080 31392 24092
rect 31444 24080 31450 24132
rect 40236 24120 40264 24151
rect 40310 24148 40316 24200
rect 40368 24188 40374 24200
rect 40880 24188 40908 24228
rect 40954 24216 40960 24268
rect 41012 24256 41018 24268
rect 41049 24259 41107 24265
rect 41049 24256 41061 24259
rect 41012 24228 41061 24256
rect 41012 24216 41018 24228
rect 41049 24225 41061 24228
rect 41095 24225 41107 24259
rect 43806 24256 43812 24268
rect 41049 24219 41107 24225
rect 41156 24228 43812 24256
rect 41156 24188 41184 24228
rect 43806 24216 43812 24228
rect 43864 24216 43870 24268
rect 45554 24256 45560 24268
rect 45526 24216 45560 24256
rect 45612 24216 45618 24268
rect 46382 24256 46388 24268
rect 46343 24228 46388 24256
rect 46382 24216 46388 24228
rect 46440 24216 46446 24268
rect 46676 24265 46704 24296
rect 46661 24259 46719 24265
rect 46661 24225 46673 24259
rect 46707 24225 46719 24259
rect 46661 24219 46719 24225
rect 40368 24160 40413 24188
rect 40880 24160 41184 24188
rect 41219 24191 41277 24197
rect 40368 24148 40374 24160
rect 41219 24157 41231 24191
rect 41265 24188 41277 24191
rect 43162 24188 43168 24200
rect 41265 24160 43168 24188
rect 41265 24157 41277 24160
rect 41219 24151 41277 24157
rect 43162 24148 43168 24160
rect 43220 24148 43226 24200
rect 43349 24191 43407 24197
rect 43349 24157 43361 24191
rect 43395 24188 43407 24191
rect 43438 24188 43444 24200
rect 43395 24160 43444 24188
rect 43395 24157 43407 24160
rect 43349 24151 43407 24157
rect 43438 24148 43444 24160
rect 43496 24148 43502 24200
rect 43530 24148 43536 24200
rect 43588 24188 43594 24200
rect 43993 24191 44051 24197
rect 43588 24160 43633 24188
rect 43588 24148 43594 24160
rect 43993 24157 44005 24191
rect 44039 24188 44051 24191
rect 45281 24191 45339 24197
rect 45281 24188 45293 24191
rect 44039 24160 45293 24188
rect 44039 24157 44051 24160
rect 43993 24151 44051 24157
rect 45281 24157 45293 24160
rect 45327 24188 45339 24191
rect 45526 24188 45554 24216
rect 45738 24188 45744 24200
rect 45327 24160 45744 24188
rect 45327 24157 45339 24160
rect 45281 24151 45339 24157
rect 45738 24148 45744 24160
rect 45796 24148 45802 24200
rect 46198 24188 46204 24200
rect 46159 24160 46204 24188
rect 46198 24148 46204 24160
rect 46256 24148 46262 24200
rect 44269 24123 44327 24129
rect 44269 24120 44281 24123
rect 40236 24092 44281 24120
rect 44269 24089 44281 24092
rect 44315 24120 44327 24123
rect 44542 24120 44548 24132
rect 44315 24092 44548 24120
rect 44315 24089 44327 24092
rect 44269 24083 44327 24089
rect 44542 24080 44548 24092
rect 44600 24080 44606 24132
rect 45557 24123 45615 24129
rect 45557 24089 45569 24123
rect 45603 24120 45615 24123
rect 45830 24120 45836 24132
rect 45603 24092 45836 24120
rect 45603 24089 45615 24092
rect 45557 24083 45615 24089
rect 45830 24080 45836 24092
rect 45888 24080 45894 24132
rect 30558 24052 30564 24064
rect 29748 24024 30564 24052
rect 30558 24012 30564 24024
rect 30616 24012 30622 24064
rect 35621 24055 35679 24061
rect 35621 24021 35633 24055
rect 35667 24052 35679 24055
rect 36170 24052 36176 24064
rect 35667 24024 36176 24052
rect 35667 24021 35679 24024
rect 35621 24015 35679 24021
rect 36170 24012 36176 24024
rect 36228 24012 36234 24064
rect 42518 24012 42524 24064
rect 42576 24052 42582 24064
rect 43441 24055 43499 24061
rect 43441 24052 43453 24055
rect 42576 24024 43453 24052
rect 42576 24012 42582 24024
rect 43441 24021 43453 24024
rect 43487 24052 43499 24055
rect 43622 24052 43628 24064
rect 43487 24024 43628 24052
rect 43487 24021 43499 24024
rect 43441 24015 43499 24021
rect 43622 24012 43628 24024
rect 43680 24012 43686 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 8754 23848 8760 23860
rect 8715 23820 8760 23848
rect 8754 23808 8760 23820
rect 8812 23808 8818 23860
rect 11054 23808 11060 23860
rect 11112 23848 11118 23860
rect 11882 23848 11888 23860
rect 11112 23820 11888 23848
rect 11112 23808 11118 23820
rect 11882 23808 11888 23820
rect 11940 23808 11946 23860
rect 18046 23848 18052 23860
rect 18007 23820 18052 23848
rect 18046 23808 18052 23820
rect 18104 23808 18110 23860
rect 18966 23848 18972 23860
rect 18927 23820 18972 23848
rect 18966 23808 18972 23820
rect 19024 23808 19030 23860
rect 19058 23808 19064 23860
rect 19116 23848 19122 23860
rect 20073 23851 20131 23857
rect 19116 23820 19161 23848
rect 19116 23808 19122 23820
rect 20073 23817 20085 23851
rect 20119 23848 20131 23851
rect 20162 23848 20168 23860
rect 20119 23820 20168 23848
rect 20119 23817 20131 23820
rect 20073 23811 20131 23817
rect 20162 23808 20168 23820
rect 20220 23808 20226 23860
rect 22278 23808 22284 23860
rect 22336 23848 22342 23860
rect 25130 23848 25136 23860
rect 22336 23820 25136 23848
rect 22336 23808 22342 23820
rect 11517 23783 11575 23789
rect 11517 23749 11529 23783
rect 11563 23780 11575 23783
rect 12434 23780 12440 23792
rect 11563 23752 12440 23780
rect 11563 23749 11575 23752
rect 11517 23743 11575 23749
rect 12434 23740 12440 23752
rect 12492 23740 12498 23792
rect 18693 23783 18751 23789
rect 18693 23749 18705 23783
rect 18739 23780 18751 23783
rect 18782 23780 18788 23792
rect 18739 23752 18788 23780
rect 18739 23749 18751 23752
rect 18693 23743 18751 23749
rect 18782 23740 18788 23752
rect 18840 23740 18846 23792
rect 1394 23712 1400 23724
rect 1355 23684 1400 23712
rect 1394 23672 1400 23684
rect 1452 23672 1458 23724
rect 8665 23715 8723 23721
rect 8665 23681 8677 23715
rect 8711 23712 8723 23715
rect 8938 23712 8944 23724
rect 8711 23684 8944 23712
rect 8711 23681 8723 23684
rect 8665 23675 8723 23681
rect 8938 23672 8944 23684
rect 8996 23672 9002 23724
rect 10965 23715 11023 23721
rect 10965 23681 10977 23715
rect 11011 23681 11023 23715
rect 13630 23712 13636 23724
rect 13591 23684 13636 23712
rect 10965 23675 11023 23681
rect 10980 23644 11008 23675
rect 13630 23672 13636 23684
rect 13688 23672 13694 23724
rect 16666 23712 16672 23724
rect 16627 23684 16672 23712
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 17678 23672 17684 23724
rect 17736 23712 17742 23724
rect 17957 23715 18015 23721
rect 17957 23712 17969 23715
rect 17736 23684 17969 23712
rect 17736 23672 17742 23684
rect 17957 23681 17969 23684
rect 18003 23681 18015 23715
rect 18138 23712 18144 23724
rect 18099 23684 18144 23712
rect 17957 23675 18015 23681
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 18874 23712 18880 23724
rect 18835 23684 18880 23712
rect 18874 23672 18880 23684
rect 18932 23672 18938 23724
rect 19978 23712 19984 23724
rect 19939 23684 19984 23712
rect 19978 23672 19984 23684
rect 20036 23672 20042 23724
rect 22756 23721 22784 23820
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 28166 23808 28172 23860
rect 28224 23808 28230 23860
rect 29546 23808 29552 23860
rect 29604 23848 29610 23860
rect 30745 23851 30803 23857
rect 30745 23848 30757 23851
rect 29604 23820 30757 23848
rect 29604 23808 29610 23820
rect 30745 23817 30757 23820
rect 30791 23848 30803 23851
rect 31294 23848 31300 23860
rect 30791 23820 31300 23848
rect 30791 23817 30803 23820
rect 30745 23811 30803 23817
rect 31294 23808 31300 23820
rect 31352 23848 31358 23860
rect 31389 23851 31447 23857
rect 31389 23848 31401 23851
rect 31352 23820 31401 23848
rect 31352 23808 31358 23820
rect 31389 23817 31401 23820
rect 31435 23817 31447 23851
rect 32858 23848 32864 23860
rect 32819 23820 32864 23848
rect 31389 23811 31447 23817
rect 32858 23808 32864 23820
rect 32916 23808 32922 23860
rect 33597 23851 33655 23857
rect 33597 23817 33609 23851
rect 33643 23848 33655 23851
rect 33778 23848 33784 23860
rect 33643 23820 33784 23848
rect 33643 23817 33655 23820
rect 33597 23811 33655 23817
rect 23014 23780 23020 23792
rect 22975 23752 23020 23780
rect 23014 23740 23020 23752
rect 23072 23740 23078 23792
rect 23474 23740 23480 23792
rect 23532 23740 23538 23792
rect 27985 23783 28043 23789
rect 27985 23749 27997 23783
rect 28031 23780 28043 23783
rect 28184 23780 28212 23808
rect 33226 23780 33232 23792
rect 28031 23752 28212 23780
rect 30024 23752 30512 23780
rect 28031 23749 28043 23752
rect 27985 23743 28043 23749
rect 21913 23715 21971 23721
rect 21913 23681 21925 23715
rect 21959 23681 21971 23715
rect 21913 23675 21971 23681
rect 22741 23715 22799 23721
rect 22741 23681 22753 23715
rect 22787 23681 22799 23715
rect 22741 23675 22799 23681
rect 28169 23715 28227 23721
rect 28169 23681 28181 23715
rect 28215 23712 28227 23715
rect 28442 23712 28448 23724
rect 28215 23684 28448 23712
rect 28215 23681 28227 23684
rect 28169 23675 28227 23681
rect 11977 23647 12035 23653
rect 11977 23644 11989 23647
rect 10980 23616 11989 23644
rect 11977 23613 11989 23616
rect 12023 23613 12035 23647
rect 13814 23644 13820 23656
rect 13775 23616 13820 23644
rect 11977 23607 12035 23613
rect 13814 23604 13820 23616
rect 13872 23604 13878 23656
rect 14090 23644 14096 23656
rect 14051 23616 14096 23644
rect 14090 23604 14096 23616
rect 14148 23604 14154 23656
rect 21928 23644 21956 23675
rect 28442 23672 28448 23684
rect 28500 23672 28506 23724
rect 28626 23672 28632 23724
rect 28684 23712 28690 23724
rect 29638 23712 29644 23724
rect 28684 23684 29644 23712
rect 28684 23672 28690 23684
rect 29638 23672 29644 23684
rect 29696 23712 29702 23724
rect 29733 23715 29791 23721
rect 29733 23712 29745 23715
rect 29696 23684 29745 23712
rect 29696 23672 29702 23684
rect 29733 23681 29745 23684
rect 29779 23681 29791 23715
rect 29733 23675 29791 23681
rect 29917 23715 29975 23721
rect 29917 23681 29929 23715
rect 29963 23712 29975 23715
rect 30024 23712 30052 23752
rect 30484 23724 30512 23752
rect 32784 23752 33232 23780
rect 29963 23684 30052 23712
rect 29963 23681 29975 23684
rect 29917 23675 29975 23681
rect 30098 23672 30104 23724
rect 30156 23712 30162 23724
rect 30377 23715 30435 23721
rect 30377 23712 30389 23715
rect 30156 23684 30389 23712
rect 30156 23672 30162 23684
rect 30377 23681 30389 23684
rect 30423 23681 30435 23715
rect 30377 23675 30435 23681
rect 30466 23672 30472 23724
rect 30524 23712 30530 23724
rect 30561 23715 30619 23721
rect 30561 23712 30573 23715
rect 30524 23684 30573 23712
rect 30524 23672 30530 23684
rect 30561 23681 30573 23684
rect 30607 23681 30619 23715
rect 30561 23675 30619 23681
rect 31018 23672 31024 23724
rect 31076 23712 31082 23724
rect 32784 23721 32812 23752
rect 33226 23740 33232 23752
rect 33284 23780 33290 23792
rect 33612 23780 33640 23811
rect 33778 23808 33784 23820
rect 33836 23808 33842 23860
rect 40954 23848 40960 23860
rect 40915 23820 40960 23848
rect 40954 23808 40960 23820
rect 41012 23808 41018 23860
rect 42518 23848 42524 23860
rect 42479 23820 42524 23848
rect 42518 23808 42524 23820
rect 42576 23808 42582 23860
rect 43162 23848 43168 23860
rect 43123 23820 43168 23848
rect 43162 23808 43168 23820
rect 43220 23808 43226 23860
rect 47486 23848 47492 23860
rect 43272 23820 47492 23848
rect 36262 23780 36268 23792
rect 33284 23752 33640 23780
rect 36223 23752 36268 23780
rect 33284 23740 33290 23752
rect 36262 23740 36268 23752
rect 36320 23740 36326 23792
rect 37642 23740 37648 23792
rect 37700 23780 37706 23792
rect 38105 23783 38163 23789
rect 38105 23780 38117 23783
rect 37700 23752 38117 23780
rect 37700 23740 37706 23752
rect 38105 23749 38117 23752
rect 38151 23780 38163 23783
rect 43272 23780 43300 23820
rect 47486 23808 47492 23820
rect 47544 23808 47550 23860
rect 46198 23780 46204 23792
rect 38151 23752 43300 23780
rect 45204 23752 46204 23780
rect 38151 23749 38163 23752
rect 38105 23743 38163 23749
rect 31205 23715 31263 23721
rect 31205 23712 31217 23715
rect 31076 23684 31217 23712
rect 31076 23672 31082 23684
rect 31205 23681 31217 23684
rect 31251 23681 31263 23715
rect 31205 23675 31263 23681
rect 31481 23715 31539 23721
rect 31481 23681 31493 23715
rect 31527 23681 31539 23715
rect 31481 23675 31539 23681
rect 32769 23715 32827 23721
rect 32769 23681 32781 23715
rect 32815 23681 32827 23715
rect 32769 23675 32827 23681
rect 33413 23715 33471 23721
rect 33413 23681 33425 23715
rect 33459 23712 33471 23715
rect 33962 23712 33968 23724
rect 33459 23684 33968 23712
rect 33459 23681 33471 23684
rect 33413 23675 33471 23681
rect 23106 23644 23112 23656
rect 21928 23616 23112 23644
rect 23106 23604 23112 23616
rect 23164 23604 23170 23656
rect 24489 23647 24547 23653
rect 24489 23613 24501 23647
rect 24535 23644 24547 23647
rect 24854 23644 24860 23656
rect 24535 23616 24860 23644
rect 24535 23613 24547 23616
rect 24489 23607 24547 23613
rect 24854 23604 24860 23616
rect 24912 23604 24918 23656
rect 28074 23604 28080 23656
rect 28132 23644 28138 23656
rect 28353 23647 28411 23653
rect 28353 23644 28365 23647
rect 28132 23616 28365 23644
rect 28132 23604 28138 23616
rect 28353 23613 28365 23616
rect 28399 23613 28411 23647
rect 28353 23607 28411 23613
rect 29825 23647 29883 23653
rect 29825 23613 29837 23647
rect 29871 23644 29883 23647
rect 31496 23644 31524 23675
rect 33962 23672 33968 23684
rect 34020 23672 34026 23724
rect 35529 23715 35587 23721
rect 35529 23681 35541 23715
rect 35575 23712 35587 23715
rect 36354 23712 36360 23724
rect 35575 23684 36360 23712
rect 35575 23681 35587 23684
rect 35529 23675 35587 23681
rect 36354 23672 36360 23684
rect 36412 23712 36418 23724
rect 37277 23715 37335 23721
rect 37277 23712 37289 23715
rect 36412 23684 37289 23712
rect 36412 23672 36418 23684
rect 37277 23681 37289 23684
rect 37323 23681 37335 23715
rect 40586 23712 40592 23724
rect 40547 23684 40592 23712
rect 37277 23675 37335 23681
rect 40586 23672 40592 23684
rect 40644 23672 40650 23724
rect 42981 23715 43039 23721
rect 42981 23681 42993 23715
rect 43027 23712 43039 23715
rect 43346 23712 43352 23724
rect 43027 23684 43352 23712
rect 43027 23681 43039 23684
rect 42981 23675 43039 23681
rect 43346 23672 43352 23684
rect 43404 23712 43410 23724
rect 43717 23715 43775 23721
rect 43717 23712 43729 23715
rect 43404 23684 43729 23712
rect 43404 23672 43410 23684
rect 43717 23681 43729 23684
rect 43763 23681 43775 23715
rect 43898 23712 43904 23724
rect 43859 23684 43904 23712
rect 43717 23675 43775 23681
rect 43898 23672 43904 23684
rect 43956 23672 43962 23724
rect 45204 23721 45232 23752
rect 46198 23740 46204 23752
rect 46256 23740 46262 23792
rect 47762 23780 47768 23792
rect 47723 23752 47768 23780
rect 47762 23740 47768 23752
rect 47820 23740 47826 23792
rect 44729 23715 44787 23721
rect 44729 23681 44741 23715
rect 44775 23712 44787 23715
rect 45189 23715 45247 23721
rect 45189 23712 45201 23715
rect 44775 23684 45201 23712
rect 44775 23681 44787 23684
rect 44729 23675 44787 23681
rect 45189 23681 45201 23684
rect 45235 23681 45247 23715
rect 47578 23712 47584 23724
rect 47539 23684 47584 23712
rect 45189 23675 45247 23681
rect 47578 23672 47584 23684
rect 47636 23672 47642 23724
rect 29871 23616 31524 23644
rect 40681 23647 40739 23653
rect 29871 23613 29883 23616
rect 29825 23607 29883 23613
rect 40681 23613 40693 23647
rect 40727 23613 40739 23647
rect 42886 23644 42892 23656
rect 42847 23616 42892 23644
rect 40681 23607 40739 23613
rect 1578 23576 1584 23588
rect 1539 23548 1584 23576
rect 1578 23536 1584 23548
rect 1636 23536 1642 23588
rect 11422 23536 11428 23588
rect 11480 23576 11486 23588
rect 11793 23579 11851 23585
rect 11793 23576 11805 23579
rect 11480 23548 11805 23576
rect 11480 23536 11486 23548
rect 11793 23545 11805 23548
rect 11839 23545 11851 23579
rect 11793 23539 11851 23545
rect 24394 23536 24400 23588
rect 24452 23576 24458 23588
rect 25222 23576 25228 23588
rect 24452 23548 25228 23576
rect 24452 23536 24458 23548
rect 25222 23536 25228 23548
rect 25280 23536 25286 23588
rect 26510 23536 26516 23588
rect 26568 23576 26574 23588
rect 40402 23576 40408 23588
rect 26568 23548 40408 23576
rect 26568 23536 26574 23548
rect 40402 23536 40408 23548
rect 40460 23536 40466 23588
rect 40696 23576 40724 23607
rect 42886 23604 42892 23616
rect 42944 23604 42950 23656
rect 45370 23644 45376 23656
rect 45331 23616 45376 23644
rect 45370 23604 45376 23616
rect 45428 23604 45434 23656
rect 45554 23604 45560 23656
rect 45612 23644 45618 23656
rect 45649 23647 45707 23653
rect 45649 23644 45661 23647
rect 45612 23616 45661 23644
rect 45612 23604 45618 23616
rect 45649 23613 45661 23616
rect 45695 23613 45707 23647
rect 45649 23607 45707 23613
rect 48038 23576 48044 23588
rect 40696 23548 48044 23576
rect 48038 23536 48044 23548
rect 48096 23536 48102 23588
rect 10781 23511 10839 23517
rect 10781 23477 10793 23511
rect 10827 23508 10839 23511
rect 11698 23508 11704 23520
rect 10827 23480 11704 23508
rect 10827 23477 10839 23480
rect 10781 23471 10839 23477
rect 11698 23468 11704 23480
rect 11756 23468 11762 23520
rect 16758 23508 16764 23520
rect 16719 23480 16764 23508
rect 16758 23468 16764 23480
rect 16816 23468 16822 23520
rect 19245 23511 19303 23517
rect 19245 23477 19257 23511
rect 19291 23508 19303 23511
rect 19426 23508 19432 23520
rect 19291 23480 19432 23508
rect 19291 23477 19303 23480
rect 19245 23471 19303 23477
rect 19426 23468 19432 23480
rect 19484 23468 19490 23520
rect 22005 23511 22063 23517
rect 22005 23477 22017 23511
rect 22051 23508 22063 23511
rect 22278 23508 22284 23520
rect 22051 23480 22284 23508
rect 22051 23477 22063 23480
rect 22005 23471 22063 23477
rect 22278 23468 22284 23480
rect 22336 23468 22342 23520
rect 27154 23468 27160 23520
rect 27212 23508 27218 23520
rect 31018 23508 31024 23520
rect 27212 23480 31024 23508
rect 27212 23468 27218 23480
rect 31018 23468 31024 23480
rect 31076 23468 31082 23520
rect 31205 23511 31263 23517
rect 31205 23477 31217 23511
rect 31251 23508 31263 23511
rect 31386 23508 31392 23520
rect 31251 23480 31392 23508
rect 31251 23477 31263 23480
rect 31205 23471 31263 23477
rect 31386 23468 31392 23480
rect 31444 23468 31450 23520
rect 44726 23468 44732 23520
rect 44784 23508 44790 23520
rect 47949 23511 48007 23517
rect 47949 23508 47961 23511
rect 44784 23480 47961 23508
rect 44784 23468 44790 23480
rect 47949 23477 47961 23480
rect 47995 23477 48007 23511
rect 47949 23471 48007 23477
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 3878 23264 3884 23316
rect 3936 23304 3942 23316
rect 12066 23304 12072 23316
rect 3936 23276 12072 23304
rect 3936 23264 3942 23276
rect 12066 23264 12072 23276
rect 12124 23264 12130 23316
rect 13078 23264 13084 23316
rect 13136 23304 13142 23316
rect 13173 23307 13231 23313
rect 13173 23304 13185 23307
rect 13136 23276 13185 23304
rect 13136 23264 13142 23276
rect 13173 23273 13185 23276
rect 13219 23273 13231 23307
rect 13173 23267 13231 23273
rect 13814 23264 13820 23316
rect 13872 23304 13878 23316
rect 14185 23307 14243 23313
rect 14185 23304 14197 23307
rect 13872 23276 14197 23304
rect 13872 23264 13878 23276
rect 14185 23273 14197 23276
rect 14231 23273 14243 23307
rect 14185 23267 14243 23273
rect 16574 23264 16580 23316
rect 16632 23304 16638 23316
rect 16853 23307 16911 23313
rect 16853 23304 16865 23307
rect 16632 23276 16865 23304
rect 16632 23264 16638 23276
rect 16853 23273 16865 23276
rect 16899 23273 16911 23307
rect 26970 23304 26976 23316
rect 26931 23276 26976 23304
rect 16853 23267 16911 23273
rect 26970 23264 26976 23276
rect 27028 23264 27034 23316
rect 30374 23264 30380 23316
rect 30432 23304 30438 23316
rect 31570 23304 31576 23316
rect 30432 23276 31576 23304
rect 30432 23264 30438 23276
rect 31570 23264 31576 23276
rect 31628 23304 31634 23316
rect 33873 23307 33931 23313
rect 33873 23304 33885 23307
rect 31628 23276 33885 23304
rect 31628 23264 31634 23276
rect 33873 23273 33885 23276
rect 33919 23273 33931 23307
rect 33873 23267 33931 23273
rect 37844 23276 41414 23304
rect 28169 23239 28227 23245
rect 28169 23205 28181 23239
rect 28215 23236 28227 23239
rect 28810 23236 28816 23248
rect 28215 23208 28816 23236
rect 28215 23205 28227 23208
rect 28169 23199 28227 23205
rect 28810 23196 28816 23208
rect 28868 23196 28874 23248
rect 11698 23168 11704 23180
rect 11659 23140 11704 23168
rect 11698 23128 11704 23140
rect 11756 23128 11762 23180
rect 12066 23128 12072 23180
rect 12124 23168 12130 23180
rect 23474 23168 23480 23180
rect 12124 23140 23480 23168
rect 12124 23128 12130 23140
rect 23474 23128 23480 23140
rect 23532 23128 23538 23180
rect 25498 23168 25504 23180
rect 25459 23140 25504 23168
rect 25498 23128 25504 23140
rect 25556 23128 25562 23180
rect 30190 23128 30196 23180
rect 30248 23168 30254 23180
rect 30248 23140 30696 23168
rect 30248 23128 30254 23140
rect 11422 23100 11428 23112
rect 11383 23072 11428 23100
rect 11422 23060 11428 23072
rect 11480 23060 11486 23112
rect 13446 23060 13452 23112
rect 13504 23100 13510 23112
rect 14093 23103 14151 23109
rect 14093 23100 14105 23103
rect 13504 23072 14105 23100
rect 13504 23060 13510 23072
rect 14093 23069 14105 23072
rect 14139 23069 14151 23103
rect 15102 23100 15108 23112
rect 15063 23072 15108 23100
rect 14093 23063 14151 23069
rect 15102 23060 15108 23072
rect 15160 23060 15166 23112
rect 16666 23060 16672 23112
rect 16724 23100 16730 23112
rect 17405 23103 17463 23109
rect 17405 23100 17417 23103
rect 16724 23072 17417 23100
rect 16724 23060 16730 23072
rect 17405 23069 17417 23072
rect 17451 23069 17463 23103
rect 19426 23100 19432 23112
rect 19387 23072 19432 23100
rect 17405 23063 17463 23069
rect 19426 23060 19432 23072
rect 19484 23060 19490 23112
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23100 19671 23103
rect 20530 23100 20536 23112
rect 19659 23072 20536 23100
rect 19659 23069 19671 23072
rect 19613 23063 19671 23069
rect 20530 23060 20536 23072
rect 20588 23060 20594 23112
rect 20898 23100 20904 23112
rect 20859 23072 20904 23100
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 22278 23060 22284 23112
rect 22336 23060 22342 23112
rect 25130 23060 25136 23112
rect 25188 23100 25194 23112
rect 25225 23103 25283 23109
rect 25225 23100 25237 23103
rect 25188 23072 25237 23100
rect 25188 23060 25194 23072
rect 25225 23069 25237 23072
rect 25271 23069 25283 23103
rect 25225 23063 25283 23069
rect 27154 23060 27160 23112
rect 27212 23100 27218 23112
rect 28169 23103 28227 23109
rect 28169 23100 28181 23103
rect 27212 23072 28181 23100
rect 27212 23060 27218 23072
rect 28169 23069 28181 23072
rect 28215 23069 28227 23103
rect 28169 23063 28227 23069
rect 28258 23060 28264 23112
rect 28316 23100 28322 23112
rect 28445 23103 28503 23109
rect 28445 23100 28457 23103
rect 28316 23072 28457 23100
rect 28316 23060 28322 23072
rect 28445 23069 28457 23072
rect 28491 23069 28503 23103
rect 30374 23100 30380 23112
rect 30335 23072 30380 23100
rect 28445 23063 28503 23069
rect 30374 23060 30380 23072
rect 30432 23060 30438 23112
rect 30668 23109 30696 23140
rect 31478 23128 31484 23180
rect 31536 23168 31542 23180
rect 32125 23171 32183 23177
rect 32125 23168 32137 23171
rect 31536 23140 32137 23168
rect 31536 23128 31542 23140
rect 32125 23137 32137 23140
rect 32171 23137 32183 23171
rect 36170 23168 36176 23180
rect 36131 23140 36176 23168
rect 32125 23131 32183 23137
rect 36170 23128 36176 23140
rect 36228 23128 36234 23180
rect 37844 23177 37872 23276
rect 41386 23236 41414 23276
rect 42886 23264 42892 23316
rect 42944 23304 42950 23316
rect 43717 23307 43775 23313
rect 43717 23304 43729 23307
rect 42944 23276 43729 23304
rect 42944 23264 42950 23276
rect 43717 23273 43729 23276
rect 43763 23273 43775 23307
rect 43717 23267 43775 23273
rect 44269 23307 44327 23313
rect 44269 23273 44281 23307
rect 44315 23304 44327 23307
rect 45370 23304 45376 23316
rect 44315 23276 45376 23304
rect 44315 23273 44327 23276
rect 44269 23267 44327 23273
rect 45370 23264 45376 23276
rect 45428 23264 45434 23316
rect 45278 23236 45284 23248
rect 41386 23208 45284 23236
rect 45278 23196 45284 23208
rect 45336 23196 45342 23248
rect 37829 23171 37887 23177
rect 37829 23137 37841 23171
rect 37875 23137 37887 23171
rect 40862 23168 40868 23180
rect 40823 23140 40868 23168
rect 37829 23131 37887 23137
rect 40862 23128 40868 23140
rect 40920 23128 40926 23180
rect 42058 23168 42064 23180
rect 42019 23140 42064 23168
rect 42058 23128 42064 23140
rect 42116 23168 42122 23180
rect 45554 23168 45560 23180
rect 42116 23140 45560 23168
rect 42116 23128 42122 23140
rect 45554 23128 45560 23140
rect 45612 23128 45618 23180
rect 45738 23128 45744 23180
rect 45796 23128 45802 23180
rect 46290 23168 46296 23180
rect 46251 23140 46296 23168
rect 46290 23128 46296 23140
rect 46348 23128 46354 23180
rect 48130 23168 48136 23180
rect 48091 23140 48136 23168
rect 48130 23128 48136 23140
rect 48188 23128 48194 23180
rect 30653 23103 30711 23109
rect 30653 23069 30665 23103
rect 30699 23069 30711 23103
rect 30653 23063 30711 23069
rect 30745 23103 30803 23109
rect 30745 23069 30757 23103
rect 30791 23100 30803 23103
rect 30926 23100 30932 23112
rect 30791 23072 30932 23100
rect 30791 23069 30803 23072
rect 30745 23063 30803 23069
rect 30926 23060 30932 23072
rect 30984 23060 30990 23112
rect 31570 23060 31576 23112
rect 31628 23100 31634 23112
rect 31665 23103 31723 23109
rect 31665 23100 31677 23103
rect 31628 23072 31677 23100
rect 31628 23060 31634 23072
rect 31665 23069 31677 23072
rect 31711 23069 31723 23103
rect 35986 23100 35992 23112
rect 35947 23072 35992 23100
rect 31665 23063 31723 23069
rect 35986 23060 35992 23072
rect 36044 23060 36050 23112
rect 40402 23100 40408 23112
rect 40363 23072 40408 23100
rect 40402 23060 40408 23072
rect 40460 23060 40466 23112
rect 43349 23103 43407 23109
rect 43349 23069 43361 23103
rect 43395 23100 43407 23103
rect 43438 23100 43444 23112
rect 43395 23072 43444 23100
rect 43395 23069 43407 23072
rect 43349 23063 43407 23069
rect 43438 23060 43444 23072
rect 43496 23060 43502 23112
rect 44453 23103 44511 23109
rect 44453 23069 44465 23103
rect 44499 23069 44511 23103
rect 44453 23063 44511 23069
rect 45189 23103 45247 23109
rect 45189 23069 45201 23103
rect 45235 23100 45247 23103
rect 45756 23100 45784 23128
rect 45235 23072 45784 23100
rect 45235 23069 45247 23072
rect 45189 23063 45247 23069
rect 12434 22992 12440 23044
rect 12492 22992 12498 23044
rect 15378 23032 15384 23044
rect 15339 23004 15384 23032
rect 15378 22992 15384 23004
rect 15436 22992 15442 23044
rect 16758 23032 16764 23044
rect 16606 23004 16764 23032
rect 16758 22992 16764 23004
rect 16816 22992 16822 23044
rect 21174 23032 21180 23044
rect 21135 23004 21180 23032
rect 21174 22992 21180 23004
rect 21232 22992 21238 23044
rect 27062 23032 27068 23044
rect 26726 23004 27068 23032
rect 27062 22992 27068 23004
rect 27120 22992 27126 23044
rect 30558 23032 30564 23044
rect 30519 23004 30564 23032
rect 30558 22992 30564 23004
rect 30616 22992 30622 23044
rect 32401 23035 32459 23041
rect 32401 23032 32413 23035
rect 31726 23004 32413 23032
rect 17494 22964 17500 22976
rect 17455 22936 17500 22964
rect 17494 22924 17500 22936
rect 17552 22924 17558 22976
rect 19334 22924 19340 22976
rect 19392 22964 19398 22976
rect 19797 22967 19855 22973
rect 19797 22964 19809 22967
rect 19392 22936 19809 22964
rect 19392 22924 19398 22936
rect 19797 22933 19809 22936
rect 19843 22933 19855 22967
rect 19797 22927 19855 22933
rect 22094 22924 22100 22976
rect 22152 22964 22158 22976
rect 22649 22967 22707 22973
rect 22649 22964 22661 22967
rect 22152 22936 22661 22964
rect 22152 22924 22158 22936
rect 22649 22933 22661 22936
rect 22695 22933 22707 22967
rect 22649 22927 22707 22933
rect 28074 22924 28080 22976
rect 28132 22964 28138 22976
rect 28353 22967 28411 22973
rect 28353 22964 28365 22967
rect 28132 22936 28365 22964
rect 28132 22924 28138 22936
rect 28353 22933 28365 22936
rect 28399 22933 28411 22967
rect 28353 22927 28411 22933
rect 30929 22967 30987 22973
rect 30929 22933 30941 22967
rect 30975 22964 30987 22967
rect 31202 22964 31208 22976
rect 30975 22936 31208 22964
rect 30975 22933 30987 22936
rect 30929 22927 30987 22933
rect 31202 22924 31208 22936
rect 31260 22924 31266 22976
rect 31481 22967 31539 22973
rect 31481 22933 31493 22967
rect 31527 22964 31539 22967
rect 31726 22964 31754 23004
rect 32401 23001 32413 23004
rect 32447 23001 32459 23035
rect 32401 22995 32459 23001
rect 33410 22992 33416 23044
rect 33468 22992 33474 23044
rect 41049 23035 41107 23041
rect 41049 23001 41061 23035
rect 41095 23001 41107 23035
rect 41049 22995 41107 23001
rect 43533 23035 43591 23041
rect 43533 23001 43545 23035
rect 43579 23032 43591 23035
rect 43622 23032 43628 23044
rect 43579 23004 43628 23032
rect 43579 23001 43591 23004
rect 43533 22995 43591 23001
rect 31527 22936 31754 22964
rect 40221 22967 40279 22973
rect 31527 22933 31539 22936
rect 31481 22927 31539 22933
rect 40221 22933 40233 22967
rect 40267 22964 40279 22967
rect 41064 22964 41092 22995
rect 43622 22992 43628 23004
rect 43680 22992 43686 23044
rect 40267 22936 41092 22964
rect 44468 22964 44496 23063
rect 45554 22992 45560 23044
rect 45612 23032 45618 23044
rect 46477 23035 46535 23041
rect 45612 23004 45657 23032
rect 45612 22992 45618 23004
rect 46477 23001 46489 23035
rect 46523 23032 46535 23035
rect 46934 23032 46940 23044
rect 46523 23004 46940 23032
rect 46523 23001 46535 23004
rect 46477 22995 46535 23001
rect 46934 22992 46940 23004
rect 46992 22992 46998 23044
rect 48130 22964 48136 22976
rect 44468 22936 48136 22964
rect 40267 22933 40279 22936
rect 40221 22927 40279 22933
rect 48130 22924 48136 22936
rect 48188 22924 48194 22976
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 12434 22720 12440 22772
rect 12492 22760 12498 22772
rect 12492 22732 12537 22760
rect 12492 22720 12498 22732
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 18417 22763 18475 22769
rect 18417 22760 18429 22763
rect 18012 22732 18429 22760
rect 18012 22720 18018 22732
rect 18417 22729 18429 22732
rect 18463 22760 18475 22763
rect 18874 22760 18880 22772
rect 18463 22732 18880 22760
rect 18463 22729 18475 22732
rect 18417 22723 18475 22729
rect 18874 22720 18880 22732
rect 18932 22760 18938 22772
rect 19150 22760 19156 22772
rect 18932 22732 19156 22760
rect 18932 22720 18938 22732
rect 19150 22720 19156 22732
rect 19208 22720 19214 22772
rect 21174 22760 21180 22772
rect 21135 22732 21180 22760
rect 21174 22720 21180 22732
rect 21232 22720 21238 22772
rect 27062 22760 27068 22772
rect 27023 22732 27068 22760
rect 27062 22720 27068 22732
rect 27120 22720 27126 22772
rect 28258 22760 28264 22772
rect 28219 22732 28264 22760
rect 28258 22720 28264 22732
rect 28316 22720 28322 22772
rect 30558 22760 30564 22772
rect 29104 22732 30564 22760
rect 17218 22692 17224 22704
rect 16592 22664 17224 22692
rect 16592 22636 16620 22664
rect 17218 22652 17224 22664
rect 17276 22652 17282 22704
rect 17494 22652 17500 22704
rect 17552 22652 17558 22704
rect 18230 22652 18236 22704
rect 18288 22692 18294 22704
rect 18288 22664 19288 22692
rect 18288 22652 18294 22664
rect 8938 22624 8944 22636
rect 8899 22596 8944 22624
rect 8938 22584 8944 22596
rect 8996 22584 9002 22636
rect 9766 22624 9772 22636
rect 9727 22596 9772 22624
rect 9766 22584 9772 22596
rect 9824 22584 9830 22636
rect 10597 22627 10655 22633
rect 10597 22593 10609 22627
rect 10643 22624 10655 22627
rect 11330 22624 11336 22636
rect 10643 22596 11336 22624
rect 10643 22593 10655 22596
rect 10597 22587 10655 22593
rect 11330 22584 11336 22596
rect 11388 22584 11394 22636
rect 11517 22627 11575 22633
rect 11517 22593 11529 22627
rect 11563 22624 11575 22627
rect 12345 22627 12403 22633
rect 12345 22624 12357 22627
rect 11563 22596 12357 22624
rect 11563 22593 11575 22596
rect 11517 22587 11575 22593
rect 12345 22593 12357 22596
rect 12391 22624 12403 22627
rect 13354 22624 13360 22636
rect 12391 22596 13360 22624
rect 12391 22593 12403 22596
rect 12345 22587 12403 22593
rect 13354 22584 13360 22596
rect 13412 22584 13418 22636
rect 13906 22624 13912 22636
rect 13867 22596 13912 22624
rect 13906 22584 13912 22596
rect 13964 22624 13970 22636
rect 16574 22624 16580 22636
rect 13964 22596 16580 22624
rect 13964 22584 13970 22596
rect 16574 22584 16580 22596
rect 16632 22584 16638 22636
rect 18782 22584 18788 22636
rect 18840 22624 18846 22636
rect 19260 22633 19288 22664
rect 20898 22652 20904 22704
rect 20956 22692 20962 22704
rect 26878 22692 26884 22704
rect 20956 22664 26884 22692
rect 20956 22652 20962 22664
rect 26878 22652 26884 22664
rect 26936 22652 26942 22704
rect 29104 22701 29132 22732
rect 30558 22720 30564 22732
rect 30616 22720 30622 22772
rect 31570 22760 31576 22772
rect 31531 22732 31576 22760
rect 31570 22720 31576 22732
rect 31628 22720 31634 22772
rect 33321 22763 33379 22769
rect 33321 22729 33333 22763
rect 33367 22760 33379 22763
rect 33410 22760 33416 22772
rect 33367 22732 33416 22760
rect 33367 22729 33379 22732
rect 33321 22723 33379 22729
rect 33410 22720 33416 22732
rect 33468 22720 33474 22772
rect 40402 22720 40408 22772
rect 40460 22760 40466 22772
rect 40773 22763 40831 22769
rect 40773 22760 40785 22763
rect 40460 22732 40785 22760
rect 40460 22720 40466 22732
rect 40773 22729 40785 22732
rect 40819 22729 40831 22763
rect 46934 22760 46940 22772
rect 46895 22732 46940 22760
rect 40773 22723 40831 22729
rect 46934 22720 46940 22732
rect 46992 22720 46998 22772
rect 48130 22760 48136 22772
rect 48091 22732 48136 22760
rect 48130 22720 48136 22732
rect 48188 22720 48194 22772
rect 29089 22695 29147 22701
rect 29089 22661 29101 22695
rect 29135 22661 29147 22695
rect 29089 22655 29147 22661
rect 29181 22695 29239 22701
rect 29181 22661 29193 22695
rect 29227 22692 29239 22695
rect 31202 22692 31208 22704
rect 29227 22664 30236 22692
rect 31163 22664 31208 22692
rect 29227 22661 29239 22664
rect 29181 22655 29239 22661
rect 30208 22636 30236 22664
rect 31202 22652 31208 22664
rect 31260 22652 31266 22704
rect 31386 22692 31392 22704
rect 31347 22664 31392 22692
rect 31386 22652 31392 22664
rect 31444 22652 31450 22704
rect 45465 22695 45523 22701
rect 45465 22661 45477 22695
rect 45511 22692 45523 22695
rect 45738 22692 45744 22704
rect 45511 22664 45744 22692
rect 45511 22661 45523 22664
rect 45465 22655 45523 22661
rect 45738 22652 45744 22664
rect 45796 22652 45802 22704
rect 46293 22695 46351 22701
rect 46293 22661 46305 22695
rect 46339 22692 46351 22695
rect 47302 22692 47308 22704
rect 46339 22664 47308 22692
rect 46339 22661 46351 22664
rect 46293 22655 46351 22661
rect 47302 22652 47308 22664
rect 47360 22652 47366 22704
rect 18969 22627 19027 22633
rect 18969 22624 18981 22627
rect 18840 22596 18981 22624
rect 18840 22584 18846 22596
rect 18969 22593 18981 22596
rect 19015 22593 19027 22627
rect 18969 22587 19027 22593
rect 19245 22627 19303 22633
rect 19245 22593 19257 22627
rect 19291 22593 19303 22627
rect 19245 22587 19303 22593
rect 20441 22627 20499 22633
rect 20441 22593 20453 22627
rect 20487 22593 20499 22627
rect 20441 22587 20499 22593
rect 21085 22627 21143 22633
rect 21085 22593 21097 22627
rect 21131 22593 21143 22627
rect 21085 22587 21143 22593
rect 21913 22627 21971 22633
rect 21913 22593 21925 22627
rect 21959 22624 21971 22627
rect 22186 22624 22192 22636
rect 21959 22596 22192 22624
rect 21959 22593 21971 22596
rect 21913 22587 21971 22593
rect 9861 22559 9919 22565
rect 9861 22525 9873 22559
rect 9907 22556 9919 22559
rect 11054 22556 11060 22568
rect 9907 22528 11060 22556
rect 9907 22525 9919 22528
rect 9861 22519 9919 22525
rect 11054 22516 11060 22528
rect 11112 22556 11118 22568
rect 11882 22556 11888 22568
rect 11112 22528 11888 22556
rect 11112 22516 11118 22528
rect 11882 22516 11888 22528
rect 11940 22516 11946 22568
rect 16666 22556 16672 22568
rect 16627 22528 16672 22556
rect 16666 22516 16672 22528
rect 16724 22516 16730 22568
rect 16942 22556 16948 22568
rect 16903 22528 16948 22556
rect 16942 22516 16948 22528
rect 17000 22516 17006 22568
rect 19058 22516 19064 22568
rect 19116 22556 19122 22568
rect 19978 22556 19984 22568
rect 19116 22528 19984 22556
rect 19116 22516 19122 22528
rect 19978 22516 19984 22528
rect 20036 22556 20042 22568
rect 20456 22556 20484 22587
rect 20036 22528 20484 22556
rect 20036 22516 20042 22528
rect 21100 22488 21128 22587
rect 22186 22584 22192 22596
rect 22244 22584 22250 22636
rect 26973 22627 27031 22633
rect 26973 22593 26985 22627
rect 27019 22624 27031 22627
rect 27338 22624 27344 22636
rect 27019 22596 27344 22624
rect 27019 22593 27031 22596
rect 26973 22587 27031 22593
rect 27338 22584 27344 22596
rect 27396 22584 27402 22636
rect 28077 22627 28135 22633
rect 28077 22593 28089 22627
rect 28123 22624 28135 22627
rect 28166 22624 28172 22636
rect 28123 22596 28172 22624
rect 28123 22593 28135 22596
rect 28077 22587 28135 22593
rect 28166 22584 28172 22596
rect 28224 22584 28230 22636
rect 28261 22627 28319 22633
rect 28261 22593 28273 22627
rect 28307 22624 28319 22627
rect 28442 22624 28448 22636
rect 28307 22596 28448 22624
rect 28307 22593 28319 22596
rect 28261 22587 28319 22593
rect 28442 22584 28448 22596
rect 28500 22624 28506 22636
rect 28902 22624 28908 22636
rect 28500 22596 28908 22624
rect 28500 22584 28506 22596
rect 28902 22584 28908 22596
rect 28960 22584 28966 22636
rect 29273 22627 29331 22633
rect 29273 22593 29285 22627
rect 29319 22593 29331 22627
rect 30190 22624 30196 22636
rect 30151 22596 30196 22624
rect 29273 22587 29331 22593
rect 22925 22559 22983 22565
rect 22925 22525 22937 22559
rect 22971 22525 22983 22559
rect 23106 22556 23112 22568
rect 23067 22528 23112 22556
rect 22925 22519 22983 22525
rect 22940 22488 22968 22519
rect 23106 22516 23112 22528
rect 23164 22516 23170 22568
rect 23474 22556 23480 22568
rect 23435 22528 23480 22556
rect 23474 22516 23480 22528
rect 23532 22516 23538 22568
rect 23842 22488 23848 22500
rect 21100 22460 22784 22488
rect 22940 22460 23848 22488
rect 9033 22423 9091 22429
rect 9033 22389 9045 22423
rect 9079 22420 9091 22423
rect 9122 22420 9128 22432
rect 9079 22392 9128 22420
rect 9079 22389 9091 22392
rect 9033 22383 9091 22389
rect 9122 22380 9128 22392
rect 9180 22380 9186 22432
rect 10134 22420 10140 22432
rect 10095 22392 10140 22420
rect 10134 22380 10140 22392
rect 10192 22380 10198 22432
rect 10686 22420 10692 22432
rect 10647 22392 10692 22420
rect 10686 22380 10692 22392
rect 10744 22380 10750 22432
rect 11606 22420 11612 22432
rect 11567 22392 11612 22420
rect 11606 22380 11612 22392
rect 11664 22380 11670 22432
rect 13998 22380 14004 22432
rect 14056 22420 14062 22432
rect 14093 22423 14151 22429
rect 14093 22420 14105 22423
rect 14056 22392 14105 22420
rect 14056 22380 14062 22392
rect 14093 22389 14105 22392
rect 14139 22389 14151 22423
rect 14093 22383 14151 22389
rect 18506 22380 18512 22432
rect 18564 22420 18570 22432
rect 18969 22423 19027 22429
rect 18969 22420 18981 22423
rect 18564 22392 18981 22420
rect 18564 22380 18570 22392
rect 18969 22389 18981 22392
rect 19015 22389 19027 22423
rect 18969 22383 19027 22389
rect 20533 22423 20591 22429
rect 20533 22389 20545 22423
rect 20579 22420 20591 22423
rect 20990 22420 20996 22432
rect 20579 22392 20996 22420
rect 20579 22389 20591 22392
rect 20533 22383 20591 22389
rect 20990 22380 20996 22392
rect 21048 22380 21054 22432
rect 22002 22420 22008 22432
rect 21963 22392 22008 22420
rect 22002 22380 22008 22392
rect 22060 22380 22066 22432
rect 22756 22420 22784 22460
rect 23842 22448 23848 22460
rect 23900 22448 23906 22500
rect 29288 22488 29316 22587
rect 30190 22584 30196 22596
rect 30248 22584 30254 22636
rect 33226 22624 33232 22636
rect 33187 22596 33232 22624
rect 33226 22584 33232 22596
rect 33284 22584 33290 22636
rect 36081 22627 36139 22633
rect 36081 22593 36093 22627
rect 36127 22624 36139 22627
rect 36354 22624 36360 22636
rect 36127 22596 36360 22624
rect 36127 22593 36139 22596
rect 36081 22587 36139 22593
rect 36354 22584 36360 22596
rect 36412 22584 36418 22636
rect 40310 22624 40316 22636
rect 40271 22596 40316 22624
rect 40310 22584 40316 22596
rect 40368 22584 40374 22636
rect 44821 22627 44879 22633
rect 44821 22593 44833 22627
rect 44867 22593 44879 22627
rect 44821 22587 44879 22593
rect 45005 22627 45063 22633
rect 45005 22593 45017 22627
rect 45051 22593 45063 22627
rect 45005 22587 45063 22593
rect 29822 22516 29828 22568
rect 29880 22556 29886 22568
rect 29917 22559 29975 22565
rect 29917 22556 29929 22559
rect 29880 22528 29929 22556
rect 29880 22516 29886 22528
rect 29917 22525 29929 22528
rect 29963 22525 29975 22559
rect 36630 22556 36636 22568
rect 36591 22528 36636 22556
rect 29917 22519 29975 22525
rect 36630 22516 36636 22528
rect 36688 22516 36694 22568
rect 42794 22516 42800 22568
rect 42852 22556 42858 22568
rect 43349 22559 43407 22565
rect 43349 22556 43361 22559
rect 42852 22528 43361 22556
rect 42852 22516 42858 22528
rect 43349 22525 43361 22528
rect 43395 22525 43407 22559
rect 43349 22519 43407 22525
rect 42886 22488 42892 22500
rect 29288 22460 42892 22488
rect 42886 22448 42892 22460
rect 42944 22448 42950 22500
rect 43530 22448 43536 22500
rect 43588 22488 43594 22500
rect 43625 22491 43683 22497
rect 43625 22488 43637 22491
rect 43588 22460 43637 22488
rect 43588 22448 43594 22460
rect 43625 22457 43637 22460
rect 43671 22457 43683 22491
rect 44836 22488 44864 22587
rect 45020 22556 45048 22587
rect 45554 22584 45560 22636
rect 45612 22624 45618 22636
rect 46845 22627 46903 22633
rect 46845 22624 46857 22627
rect 45612 22596 46857 22624
rect 45612 22584 45618 22596
rect 46845 22593 46857 22596
rect 46891 22593 46903 22627
rect 46845 22587 46903 22593
rect 47581 22627 47639 22633
rect 47581 22593 47593 22627
rect 47627 22624 47639 22627
rect 47762 22624 47768 22636
rect 47627 22596 47768 22624
rect 47627 22593 47639 22596
rect 47581 22587 47639 22593
rect 47762 22584 47768 22596
rect 47820 22584 47826 22636
rect 47210 22556 47216 22568
rect 45020 22528 47216 22556
rect 47210 22516 47216 22528
rect 47268 22516 47274 22568
rect 47854 22556 47860 22568
rect 47815 22528 47860 22556
rect 47854 22516 47860 22528
rect 47912 22516 47918 22568
rect 47946 22488 47952 22500
rect 44836 22460 47952 22488
rect 43625 22451 43683 22457
rect 47946 22448 47952 22460
rect 48004 22448 48010 22500
rect 23474 22420 23480 22432
rect 22756 22392 23480 22420
rect 23474 22380 23480 22392
rect 23532 22380 23538 22432
rect 29454 22420 29460 22432
rect 29415 22392 29460 22420
rect 29454 22380 29460 22392
rect 29512 22380 29518 22432
rect 40037 22423 40095 22429
rect 40037 22389 40049 22423
rect 40083 22420 40095 22423
rect 40494 22420 40500 22432
rect 40083 22392 40500 22420
rect 40083 22389 40095 22392
rect 40037 22383 40095 22389
rect 40494 22380 40500 22392
rect 40552 22380 40558 22432
rect 43714 22380 43720 22432
rect 43772 22420 43778 22432
rect 43809 22423 43867 22429
rect 43809 22420 43821 22423
rect 43772 22392 43821 22420
rect 43772 22380 43778 22392
rect 43809 22389 43821 22392
rect 43855 22389 43867 22423
rect 43809 22383 43867 22389
rect 44913 22423 44971 22429
rect 44913 22389 44925 22423
rect 44959 22420 44971 22423
rect 47578 22420 47584 22432
rect 44959 22392 47584 22420
rect 44959 22389 44971 22392
rect 44913 22383 44971 22389
rect 47578 22380 47584 22392
rect 47636 22420 47642 22432
rect 47673 22423 47731 22429
rect 47673 22420 47685 22423
rect 47636 22392 47685 22420
rect 47636 22380 47642 22392
rect 47673 22389 47685 22392
rect 47719 22389 47731 22423
rect 47673 22383 47731 22389
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 10134 22176 10140 22228
rect 10192 22216 10198 22228
rect 10302 22219 10360 22225
rect 10302 22216 10314 22219
rect 10192 22188 10314 22216
rect 10192 22176 10198 22188
rect 10302 22185 10314 22188
rect 10348 22185 10360 22219
rect 10302 22179 10360 22185
rect 16942 22176 16948 22228
rect 17000 22216 17006 22228
rect 17957 22219 18015 22225
rect 17957 22216 17969 22219
rect 17000 22188 17969 22216
rect 17000 22176 17006 22188
rect 17957 22185 17969 22188
rect 18003 22185 18015 22219
rect 17957 22179 18015 22185
rect 23106 22176 23112 22228
rect 23164 22216 23170 22228
rect 25406 22225 25412 22228
rect 23201 22219 23259 22225
rect 23201 22216 23213 22219
rect 23164 22188 23213 22216
rect 23164 22176 23170 22188
rect 23201 22185 23213 22188
rect 23247 22185 23259 22219
rect 23201 22179 23259 22185
rect 25396 22219 25412 22225
rect 25396 22185 25408 22219
rect 25396 22179 25412 22185
rect 25406 22176 25412 22179
rect 25464 22176 25470 22228
rect 26878 22176 26884 22228
rect 26936 22216 26942 22228
rect 31938 22216 31944 22228
rect 26936 22188 31944 22216
rect 26936 22176 26942 22188
rect 31938 22176 31944 22188
rect 31996 22176 32002 22228
rect 13096 22120 14228 22148
rect 10045 22083 10103 22089
rect 10045 22049 10057 22083
rect 10091 22080 10103 22083
rect 10686 22080 10692 22092
rect 10091 22052 10692 22080
rect 10091 22049 10103 22052
rect 10045 22043 10103 22049
rect 10686 22040 10692 22052
rect 10744 22040 10750 22092
rect 11054 22040 11060 22092
rect 11112 22080 11118 22092
rect 11790 22080 11796 22092
rect 11112 22052 11796 22080
rect 11112 22040 11118 22052
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 13096 22080 13124 22120
rect 12360 22052 13124 22080
rect 12360 22024 12388 22052
rect 13170 22040 13176 22092
rect 13228 22080 13234 22092
rect 14093 22083 14151 22089
rect 14093 22080 14105 22083
rect 13228 22052 14105 22080
rect 13228 22040 13234 22052
rect 14093 22049 14105 22052
rect 14139 22049 14151 22083
rect 14200 22080 14228 22120
rect 42886 22108 42892 22160
rect 42944 22148 42950 22160
rect 42944 22120 44036 22148
rect 42944 22108 42950 22120
rect 17681 22083 17739 22089
rect 14200 22052 16436 22080
rect 14093 22043 14151 22049
rect 8938 22012 8944 22024
rect 8899 21984 8944 22012
rect 8938 21972 8944 21984
rect 8996 21972 9002 22024
rect 12342 22012 12348 22024
rect 12303 21984 12348 22012
rect 12342 21972 12348 21984
rect 12400 21972 12406 22024
rect 13354 22012 13360 22024
rect 13315 21984 13360 22012
rect 13354 21972 13360 21984
rect 13412 22012 13418 22024
rect 13998 22012 14004 22024
rect 13412 21984 14004 22012
rect 13412 21972 13418 21984
rect 13998 21972 14004 21984
rect 14056 21972 14062 22024
rect 16408 22021 16436 22052
rect 17681 22049 17693 22083
rect 17727 22080 17739 22083
rect 18138 22080 18144 22092
rect 17727 22052 18144 22080
rect 17727 22049 17739 22052
rect 17681 22043 17739 22049
rect 18138 22040 18144 22052
rect 18196 22040 18202 22092
rect 20990 22080 20996 22092
rect 20951 22052 20996 22080
rect 20990 22040 20996 22052
rect 21048 22040 21054 22092
rect 24964 22080 25268 22094
rect 26786 22080 26792 22092
rect 24964 22066 26792 22080
rect 16393 22015 16451 22021
rect 16393 21981 16405 22015
rect 16439 22012 16451 22015
rect 17589 22015 17647 22021
rect 16439 21984 16574 22012
rect 16439 21981 16451 21984
rect 16393 21975 16451 21981
rect 14 21904 20 21956
rect 72 21944 78 21956
rect 8846 21944 8852 21956
rect 72 21916 8852 21944
rect 72 21904 78 21916
rect 8846 21904 8852 21916
rect 8904 21904 8910 21956
rect 11606 21944 11612 21956
rect 11546 21916 11612 21944
rect 11606 21904 11612 21916
rect 11664 21904 11670 21956
rect 11716 21916 12572 21944
rect 8754 21836 8760 21888
rect 8812 21876 8818 21888
rect 9033 21879 9091 21885
rect 9033 21876 9045 21879
rect 8812 21848 9045 21876
rect 8812 21836 8818 21848
rect 9033 21845 9045 21848
rect 9079 21845 9091 21879
rect 9033 21839 9091 21845
rect 9766 21836 9772 21888
rect 9824 21876 9830 21888
rect 11054 21876 11060 21888
rect 9824 21848 11060 21876
rect 9824 21836 9830 21848
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 11330 21836 11336 21888
rect 11388 21876 11394 21888
rect 11716 21876 11744 21916
rect 12544 21885 12572 21916
rect 13630 21904 13636 21956
rect 13688 21944 13694 21956
rect 14277 21947 14335 21953
rect 14277 21944 14289 21947
rect 13688 21916 14289 21944
rect 13688 21904 13694 21916
rect 14277 21913 14289 21916
rect 14323 21913 14335 21947
rect 14277 21907 14335 21913
rect 15933 21947 15991 21953
rect 15933 21913 15945 21947
rect 15979 21944 15991 21947
rect 16206 21944 16212 21956
rect 15979 21916 16212 21944
rect 15979 21913 15991 21916
rect 15933 21907 15991 21913
rect 16206 21904 16212 21916
rect 16264 21904 16270 21956
rect 16546 21944 16574 21984
rect 17589 21981 17601 22015
rect 17635 22012 17647 22015
rect 17954 22012 17960 22024
rect 17635 21984 17960 22012
rect 17635 21981 17647 21984
rect 17589 21975 17647 21981
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 18417 22015 18475 22021
rect 18417 21981 18429 22015
rect 18463 22012 18475 22015
rect 18506 22012 18512 22024
rect 18463 21984 18512 22012
rect 18463 21981 18475 21984
rect 18417 21975 18475 21981
rect 18506 21972 18512 21984
rect 18564 21972 18570 22024
rect 18601 22015 18659 22021
rect 18601 21981 18613 22015
rect 18647 22012 18659 22015
rect 19334 22012 19340 22024
rect 18647 21984 19340 22012
rect 18647 21981 18659 21984
rect 18601 21975 18659 21981
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 20806 22012 20812 22024
rect 20767 21984 20812 22012
rect 20806 21972 20812 21984
rect 20864 21972 20870 22024
rect 22186 21972 22192 22024
rect 22244 22012 22250 22024
rect 23109 22015 23167 22021
rect 23109 22012 23121 22015
rect 22244 21984 23121 22012
rect 22244 21972 22250 21984
rect 23109 21981 23121 21984
rect 23155 22012 23167 22015
rect 24964 22012 24992 22066
rect 25240 22052 26792 22066
rect 26786 22040 26792 22052
rect 26844 22040 26850 22092
rect 26881 22083 26939 22089
rect 26881 22049 26893 22083
rect 26927 22080 26939 22083
rect 28074 22080 28080 22092
rect 26927 22052 28080 22080
rect 26927 22049 26939 22052
rect 26881 22043 26939 22049
rect 28074 22040 28080 22052
rect 28132 22040 28138 22092
rect 28997 22083 29055 22089
rect 28997 22080 29009 22083
rect 28184 22052 29009 22080
rect 25130 22012 25136 22024
rect 23155 21984 24992 22012
rect 25091 21984 25136 22012
rect 23155 21981 23167 21984
rect 23109 21975 23167 21981
rect 25130 21972 25136 21984
rect 25188 21972 25194 22024
rect 27338 22012 27344 22024
rect 26542 21984 26924 22012
rect 27299 21984 27344 22012
rect 22649 21947 22707 21953
rect 16546 21916 20944 21944
rect 20916 21888 20944 21916
rect 22649 21913 22661 21947
rect 22695 21944 22707 21947
rect 25682 21944 25688 21956
rect 22695 21916 25688 21944
rect 22695 21913 22707 21916
rect 22649 21907 22707 21913
rect 25682 21904 25688 21916
rect 25740 21904 25746 21956
rect 26896 21944 26924 21984
rect 27338 21972 27344 21984
rect 27396 21972 27402 22024
rect 28184 22021 28212 22052
rect 28997 22049 29009 22052
rect 29043 22049 29055 22083
rect 42794 22080 42800 22092
rect 42755 22052 42800 22080
rect 28997 22043 29055 22049
rect 42794 22040 42800 22052
rect 42852 22080 42858 22092
rect 43901 22083 43959 22089
rect 43901 22080 43913 22083
rect 42852 22052 43913 22080
rect 42852 22040 42858 22052
rect 43901 22049 43913 22052
rect 43947 22049 43959 22083
rect 44008 22080 44036 22120
rect 47581 22083 47639 22089
rect 47581 22080 47593 22083
rect 44008 22052 47593 22080
rect 43901 22043 43959 22049
rect 47581 22049 47593 22052
rect 47627 22049 47639 22083
rect 47581 22043 47639 22049
rect 28169 22015 28227 22021
rect 28169 21981 28181 22015
rect 28215 21981 28227 22015
rect 28810 22012 28816 22024
rect 28771 21984 28816 22012
rect 28169 21975 28227 21981
rect 28810 21972 28816 21984
rect 28868 21972 28874 22024
rect 34146 21972 34152 22024
rect 34204 22012 34210 22024
rect 34885 22015 34943 22021
rect 34885 22012 34897 22015
rect 34204 21984 34897 22012
rect 34204 21972 34210 21984
rect 34885 21981 34897 21984
rect 34931 21981 34943 22015
rect 40310 22012 40316 22024
rect 40271 21984 40316 22012
rect 34885 21975 34943 21981
rect 40310 21972 40316 21984
rect 40368 21972 40374 22024
rect 40494 22012 40500 22024
rect 40455 21984 40500 22012
rect 40494 21972 40500 21984
rect 40552 21972 40558 22024
rect 42610 21972 42616 22024
rect 42668 22012 42674 22024
rect 42705 22015 42763 22021
rect 42705 22012 42717 22015
rect 42668 21984 42717 22012
rect 42668 21972 42674 21984
rect 42705 21981 42717 21984
rect 42751 21981 42763 22015
rect 42705 21975 42763 21981
rect 42889 22015 42947 22021
rect 42889 21981 42901 22015
rect 42935 22012 42947 22015
rect 42978 22012 42984 22024
rect 42935 21984 42984 22012
rect 42935 21981 42947 21984
rect 42889 21975 42947 21981
rect 42978 21972 42984 21984
rect 43036 21972 43042 22024
rect 43349 22015 43407 22021
rect 43349 21981 43361 22015
rect 43395 21981 43407 22015
rect 43530 22012 43536 22024
rect 43491 21984 43536 22012
rect 43349 21975 43407 21981
rect 27433 21947 27491 21953
rect 27433 21944 27445 21947
rect 26896 21916 27445 21944
rect 27433 21913 27445 21916
rect 27479 21913 27491 21947
rect 28629 21947 28687 21953
rect 27433 21907 27491 21913
rect 27816 21916 28580 21944
rect 11388 21848 11744 21876
rect 12529 21879 12587 21885
rect 11388 21836 11394 21848
rect 12529 21845 12541 21879
rect 12575 21845 12587 21879
rect 12529 21839 12587 21845
rect 13449 21879 13507 21885
rect 13449 21845 13461 21879
rect 13495 21876 13507 21879
rect 14366 21876 14372 21888
rect 13495 21848 14372 21876
rect 13495 21845 13507 21848
rect 13449 21839 13507 21845
rect 14366 21836 14372 21848
rect 14424 21836 14430 21888
rect 16577 21879 16635 21885
rect 16577 21845 16589 21879
rect 16623 21876 16635 21879
rect 16850 21876 16856 21888
rect 16623 21848 16856 21876
rect 16623 21845 16635 21848
rect 16577 21839 16635 21845
rect 16850 21836 16856 21848
rect 16908 21836 16914 21888
rect 18138 21836 18144 21888
rect 18196 21876 18202 21888
rect 18509 21879 18567 21885
rect 18509 21876 18521 21879
rect 18196 21848 18521 21876
rect 18196 21836 18202 21848
rect 18509 21845 18521 21848
rect 18555 21845 18567 21879
rect 18509 21839 18567 21845
rect 20898 21836 20904 21888
rect 20956 21876 20962 21888
rect 22094 21876 22100 21888
rect 20956 21848 22100 21876
rect 20956 21836 20962 21848
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 26786 21836 26792 21888
rect 26844 21876 26850 21888
rect 27816 21876 27844 21916
rect 27982 21876 27988 21888
rect 26844 21848 27844 21876
rect 27943 21848 27988 21876
rect 26844 21836 26850 21848
rect 27982 21836 27988 21848
rect 28040 21836 28046 21888
rect 28552 21876 28580 21916
rect 28629 21913 28641 21947
rect 28675 21944 28687 21947
rect 29454 21944 29460 21956
rect 28675 21916 29460 21944
rect 28675 21913 28687 21916
rect 28629 21907 28687 21913
rect 29454 21904 29460 21916
rect 29512 21904 29518 21956
rect 40589 21947 40647 21953
rect 40589 21944 40601 21947
rect 40512 21916 40601 21944
rect 40512 21888 40540 21916
rect 40589 21913 40601 21916
rect 40635 21913 40647 21947
rect 43364 21944 43392 21975
rect 43530 21972 43536 21984
rect 43588 21972 43594 22024
rect 45557 22015 45615 22021
rect 45557 21981 45569 22015
rect 45603 21981 45615 22015
rect 46014 22012 46020 22024
rect 45975 21984 46020 22012
rect 45557 21975 45615 21981
rect 43806 21944 43812 21956
rect 43364 21916 43812 21944
rect 40589 21907 40647 21913
rect 43806 21904 43812 21916
rect 43864 21904 43870 21956
rect 45572 21944 45600 21975
rect 46014 21972 46020 21984
rect 46072 21972 46078 22024
rect 46198 21972 46204 22024
rect 46256 22012 46262 22024
rect 46293 22015 46351 22021
rect 46293 22012 46305 22015
rect 46256 21984 46305 22012
rect 46256 21972 46262 21984
rect 46293 21981 46305 21984
rect 46339 21981 46351 22015
rect 47302 22012 47308 22024
rect 47263 21984 47308 22012
rect 46293 21975 46351 21981
rect 47302 21972 47308 21984
rect 47360 21972 47366 22024
rect 48038 21944 48044 21956
rect 45572 21916 48044 21944
rect 48038 21904 48044 21916
rect 48096 21904 48102 21956
rect 29270 21876 29276 21888
rect 28552 21848 29276 21876
rect 29270 21836 29276 21848
rect 29328 21836 29334 21888
rect 34698 21876 34704 21888
rect 34659 21848 34704 21876
rect 34698 21836 34704 21848
rect 34756 21836 34762 21888
rect 40494 21836 40500 21888
rect 40552 21836 40558 21888
rect 43346 21836 43352 21888
rect 43404 21876 43410 21888
rect 43533 21879 43591 21885
rect 43533 21876 43545 21879
rect 43404 21848 43545 21876
rect 43404 21836 43410 21848
rect 43533 21845 43545 21848
rect 43579 21845 43591 21879
rect 43533 21839 43591 21845
rect 45373 21879 45431 21885
rect 45373 21845 45385 21879
rect 45419 21876 45431 21879
rect 46382 21876 46388 21888
rect 45419 21848 46388 21876
rect 45419 21845 45431 21848
rect 45373 21839 45431 21845
rect 46382 21836 46388 21848
rect 46440 21836 46446 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 3050 21632 3056 21684
rect 3108 21672 3114 21684
rect 33321 21675 33379 21681
rect 33321 21672 33333 21675
rect 3108 21644 33333 21672
rect 3108 21632 3114 21644
rect 33321 21641 33333 21644
rect 33367 21641 33379 21675
rect 34146 21672 34152 21684
rect 34107 21644 34152 21672
rect 33321 21635 33379 21641
rect 8754 21604 8760 21616
rect 8715 21576 8760 21604
rect 8754 21564 8760 21576
rect 8812 21564 8818 21616
rect 8938 21564 8944 21616
rect 8996 21604 9002 21616
rect 13354 21604 13360 21616
rect 8996 21576 13360 21604
rect 8996 21564 9002 21576
rect 13354 21564 13360 21576
rect 13412 21604 13418 21616
rect 13630 21604 13636 21616
rect 13412 21576 13492 21604
rect 13591 21576 13636 21604
rect 13412 21564 13418 21576
rect 11330 21496 11336 21548
rect 11388 21536 11394 21548
rect 11517 21539 11575 21545
rect 11517 21536 11529 21539
rect 11388 21508 11529 21536
rect 11388 21496 11394 21508
rect 11517 21505 11529 21508
rect 11563 21505 11575 21539
rect 13464 21536 13492 21576
rect 13630 21564 13636 21576
rect 13688 21564 13694 21616
rect 14366 21604 14372 21616
rect 14327 21576 14372 21604
rect 14366 21564 14372 21576
rect 14424 21564 14430 21616
rect 18138 21604 18144 21616
rect 18099 21576 18144 21604
rect 18138 21564 18144 21576
rect 18196 21564 18202 21616
rect 22002 21604 22008 21616
rect 21963 21576 22008 21604
rect 22002 21564 22008 21576
rect 22060 21564 22066 21616
rect 27709 21607 27767 21613
rect 27709 21573 27721 21607
rect 27755 21604 27767 21607
rect 27982 21604 27988 21616
rect 27755 21576 27988 21604
rect 27755 21573 27767 21576
rect 27709 21567 27767 21573
rect 27982 21564 27988 21576
rect 28040 21564 28046 21616
rect 28166 21564 28172 21616
rect 28224 21564 28230 21616
rect 13541 21539 13599 21545
rect 13541 21536 13553 21539
rect 13464 21508 13553 21536
rect 11517 21499 11575 21505
rect 13541 21505 13553 21508
rect 13587 21505 13599 21539
rect 16022 21536 16028 21548
rect 15983 21508 16028 21536
rect 13541 21499 13599 21505
rect 16022 21496 16028 21508
rect 16080 21496 16086 21548
rect 16850 21536 16856 21548
rect 16811 21508 16856 21536
rect 16850 21496 16856 21508
rect 16908 21496 16914 21548
rect 19242 21496 19248 21548
rect 19300 21496 19306 21548
rect 20809 21539 20867 21545
rect 20809 21505 20821 21539
rect 20855 21536 20867 21539
rect 20898 21536 20904 21548
rect 20855 21508 20904 21536
rect 20855 21505 20867 21508
rect 20809 21499 20867 21505
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 21726 21496 21732 21548
rect 21784 21536 21790 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21784 21508 21833 21536
rect 21784 21496 21790 21508
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 25130 21496 25136 21548
rect 25188 21536 25194 21548
rect 27433 21539 27491 21545
rect 27433 21536 27445 21539
rect 25188 21508 27445 21536
rect 25188 21496 25194 21508
rect 27433 21505 27445 21508
rect 27479 21505 27491 21539
rect 32306 21536 32312 21548
rect 32267 21508 32312 21536
rect 27433 21499 27491 21505
rect 32306 21496 32312 21508
rect 32364 21496 32370 21548
rect 8573 21471 8631 21477
rect 8573 21437 8585 21471
rect 8619 21437 8631 21471
rect 8573 21431 8631 21437
rect 8588 21400 8616 21431
rect 8846 21428 8852 21480
rect 8904 21468 8910 21480
rect 9033 21471 9091 21477
rect 9033 21468 9045 21471
rect 8904 21440 9045 21468
rect 8904 21428 8910 21440
rect 9033 21437 9045 21440
rect 9079 21437 9091 21471
rect 14182 21468 14188 21480
rect 14143 21440 14188 21468
rect 9033 21431 9091 21437
rect 14182 21428 14188 21440
rect 14240 21428 14246 21480
rect 17218 21428 17224 21480
rect 17276 21468 17282 21480
rect 17865 21471 17923 21477
rect 17865 21468 17877 21471
rect 17276 21440 17877 21468
rect 17276 21428 17282 21440
rect 17865 21437 17877 21440
rect 17911 21437 17923 21471
rect 17865 21431 17923 21437
rect 18782 21428 18788 21480
rect 18840 21468 18846 21480
rect 19613 21471 19671 21477
rect 19613 21468 19625 21471
rect 18840 21440 19625 21468
rect 18840 21428 18846 21440
rect 19613 21437 19625 21440
rect 19659 21437 19671 21471
rect 22281 21471 22339 21477
rect 22281 21468 22293 21471
rect 19613 21431 19671 21437
rect 22066 21440 22293 21468
rect 10962 21400 10968 21412
rect 8588 21372 10968 21400
rect 10962 21360 10968 21372
rect 11020 21360 11026 21412
rect 11422 21360 11428 21412
rect 11480 21400 11486 21412
rect 11517 21403 11575 21409
rect 11517 21400 11529 21403
rect 11480 21372 11529 21400
rect 11480 21360 11486 21372
rect 11517 21369 11529 21372
rect 11563 21369 11575 21403
rect 16666 21400 16672 21412
rect 16627 21372 16672 21400
rect 11517 21363 11575 21369
rect 16666 21360 16672 21372
rect 16724 21360 16730 21412
rect 22066 21400 22094 21440
rect 22281 21437 22293 21440
rect 22327 21437 22339 21471
rect 22281 21431 22339 21437
rect 28902 21428 28908 21480
rect 28960 21468 28966 21480
rect 29181 21471 29239 21477
rect 29181 21468 29193 21471
rect 28960 21440 29193 21468
rect 28960 21428 28966 21440
rect 29181 21437 29193 21440
rect 29227 21437 29239 21471
rect 29181 21431 29239 21437
rect 19168 21372 22094 21400
rect 17034 21292 17040 21344
rect 17092 21332 17098 21344
rect 19168 21332 19196 21372
rect 20898 21332 20904 21344
rect 17092 21304 19196 21332
rect 20859 21304 20904 21332
rect 17092 21292 17098 21304
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 31846 21292 31852 21344
rect 31904 21332 31910 21344
rect 32125 21335 32183 21341
rect 32125 21332 32137 21335
rect 31904 21304 32137 21332
rect 31904 21292 31910 21304
rect 32125 21301 32137 21304
rect 32171 21301 32183 21335
rect 33336 21332 33364 21635
rect 34146 21632 34152 21644
rect 34204 21632 34210 21684
rect 43073 21675 43131 21681
rect 43073 21641 43085 21675
rect 43119 21672 43131 21675
rect 43530 21672 43536 21684
rect 43119 21644 43536 21672
rect 43119 21641 43131 21644
rect 43073 21635 43131 21641
rect 43530 21632 43536 21644
rect 43588 21632 43594 21684
rect 47762 21672 47768 21684
rect 47723 21644 47768 21672
rect 47762 21632 47768 21644
rect 47820 21632 47826 21684
rect 47946 21672 47952 21684
rect 47907 21644 47952 21672
rect 47946 21632 47952 21644
rect 48004 21632 48010 21684
rect 34698 21564 34704 21616
rect 34756 21604 34762 21616
rect 34793 21607 34851 21613
rect 34793 21604 34805 21607
rect 34756 21576 34805 21604
rect 34756 21564 34762 21576
rect 34793 21573 34805 21576
rect 34839 21573 34851 21607
rect 34793 21567 34851 21573
rect 42978 21564 42984 21616
rect 43036 21604 43042 21616
rect 47026 21604 47032 21616
rect 43036 21576 47032 21604
rect 43036 21564 43042 21576
rect 33689 21539 33747 21545
rect 33689 21505 33701 21539
rect 33735 21536 33747 21539
rect 33778 21536 33784 21548
rect 33735 21508 33784 21536
rect 33735 21505 33747 21508
rect 33689 21499 33747 21505
rect 33778 21496 33784 21508
rect 33836 21496 33842 21548
rect 42610 21496 42616 21548
rect 42668 21536 42674 21548
rect 43088 21545 43116 21576
rect 47026 21564 47032 21576
rect 47084 21564 47090 21616
rect 47486 21564 47492 21616
rect 47544 21604 47550 21616
rect 47854 21604 47860 21616
rect 47544 21576 47860 21604
rect 47544 21564 47550 21576
rect 47854 21564 47860 21576
rect 47912 21564 47918 21616
rect 42889 21539 42947 21545
rect 42889 21536 42901 21539
rect 42668 21508 42901 21536
rect 42668 21496 42674 21508
rect 42889 21505 42901 21508
rect 42935 21505 42947 21539
rect 42889 21499 42947 21505
rect 43073 21539 43131 21545
rect 43073 21505 43085 21539
rect 43119 21505 43131 21539
rect 43714 21536 43720 21548
rect 43675 21508 43720 21536
rect 43073 21499 43131 21505
rect 43714 21496 43720 21508
rect 43772 21496 43778 21548
rect 44726 21536 44732 21548
rect 44687 21508 44732 21536
rect 44726 21496 44732 21508
rect 44784 21496 44790 21548
rect 47210 21496 47216 21548
rect 47268 21536 47274 21548
rect 47581 21539 47639 21545
rect 47581 21536 47593 21539
rect 47268 21508 47593 21536
rect 47268 21496 47274 21508
rect 47581 21505 47593 21508
rect 47627 21505 47639 21539
rect 47581 21499 47639 21505
rect 34514 21428 34520 21480
rect 34572 21468 34578 21480
rect 34701 21471 34759 21477
rect 34701 21468 34713 21471
rect 34572 21440 34713 21468
rect 34572 21428 34578 21440
rect 34701 21437 34713 21440
rect 34747 21437 34759 21471
rect 43806 21468 43812 21480
rect 43767 21440 43812 21468
rect 34701 21431 34759 21437
rect 43806 21428 43812 21440
rect 43864 21428 43870 21480
rect 44634 21468 44640 21480
rect 44100 21440 44640 21468
rect 35253 21403 35311 21409
rect 35253 21369 35265 21403
rect 35299 21400 35311 21403
rect 35894 21400 35900 21412
rect 35299 21372 35900 21400
rect 35299 21369 35311 21372
rect 35253 21363 35311 21369
rect 35894 21360 35900 21372
rect 35952 21400 35958 21412
rect 42702 21400 42708 21412
rect 35952 21372 42708 21400
rect 35952 21360 35958 21372
rect 42702 21360 42708 21372
rect 42760 21360 42766 21412
rect 44100 21409 44128 21440
rect 44634 21428 44640 21440
rect 44692 21468 44698 21480
rect 45189 21471 45247 21477
rect 45189 21468 45201 21471
rect 44692 21440 45201 21468
rect 44692 21428 44698 21440
rect 45189 21437 45201 21440
rect 45235 21437 45247 21471
rect 45189 21431 45247 21437
rect 45373 21471 45431 21477
rect 45373 21437 45385 21471
rect 45419 21437 45431 21471
rect 46842 21468 46848 21480
rect 46803 21440 46848 21468
rect 45373 21431 45431 21437
rect 44085 21403 44143 21409
rect 44085 21369 44097 21403
rect 44131 21369 44143 21403
rect 44085 21363 44143 21369
rect 44545 21403 44603 21409
rect 44545 21369 44557 21403
rect 44591 21400 44603 21403
rect 45388 21400 45416 21431
rect 46842 21428 46848 21440
rect 46900 21428 46906 21480
rect 44591 21372 45416 21400
rect 44591 21369 44603 21372
rect 44545 21363 44603 21369
rect 33781 21335 33839 21341
rect 33781 21332 33793 21335
rect 33336 21304 33793 21332
rect 32125 21295 32183 21301
rect 33781 21301 33793 21304
rect 33827 21301 33839 21335
rect 33781 21295 33839 21301
rect 40310 21292 40316 21344
rect 40368 21332 40374 21344
rect 48133 21335 48191 21341
rect 48133 21332 48145 21335
rect 40368 21304 48145 21332
rect 40368 21292 40374 21304
rect 48133 21301 48145 21304
rect 48179 21301 48191 21335
rect 48133 21295 48191 21301
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 3418 21088 3424 21140
rect 3476 21128 3482 21140
rect 17034 21128 17040 21140
rect 3476 21100 17040 21128
rect 3476 21088 3482 21100
rect 17034 21088 17040 21100
rect 17092 21088 17098 21140
rect 17218 21128 17224 21140
rect 17179 21100 17224 21128
rect 17218 21088 17224 21100
rect 17276 21088 17282 21140
rect 19242 21088 19248 21140
rect 19300 21128 19306 21140
rect 19337 21131 19395 21137
rect 19337 21128 19349 21131
rect 19300 21100 19349 21128
rect 19300 21088 19306 21100
rect 19337 21097 19349 21100
rect 19383 21097 19395 21131
rect 23842 21128 23848 21140
rect 23803 21100 23848 21128
rect 19337 21091 19395 21097
rect 23842 21088 23848 21100
rect 23900 21088 23906 21140
rect 26881 21131 26939 21137
rect 26881 21097 26893 21131
rect 26927 21128 26939 21131
rect 27338 21128 27344 21140
rect 26927 21100 27344 21128
rect 26927 21097 26939 21100
rect 26881 21091 26939 21097
rect 27338 21088 27344 21100
rect 27396 21088 27402 21140
rect 27801 21131 27859 21137
rect 27801 21097 27813 21131
rect 27847 21128 27859 21131
rect 28166 21128 28172 21140
rect 27847 21100 28172 21128
rect 27847 21097 27859 21100
rect 27801 21091 27859 21097
rect 28166 21088 28172 21100
rect 28224 21088 28230 21140
rect 46750 21128 46756 21140
rect 28276 21100 46756 21128
rect 2590 21020 2596 21072
rect 2648 21060 2654 21072
rect 2648 21032 6914 21060
rect 2648 21020 2654 21032
rect 6886 20992 6914 21032
rect 25682 21020 25688 21072
rect 25740 21060 25746 21072
rect 28276 21060 28304 21100
rect 46750 21088 46756 21100
rect 46808 21088 46814 21140
rect 46198 21060 46204 21072
rect 25740 21032 28304 21060
rect 28920 21032 30236 21060
rect 25740 21020 25746 21032
rect 28920 20992 28948 21032
rect 30208 21004 30236 21032
rect 31864 21032 46204 21060
rect 30190 20992 30196 21004
rect 6886 20964 28948 20992
rect 30151 20964 30196 20992
rect 30190 20952 30196 20964
rect 30248 20952 30254 21004
rect 31202 20992 31208 21004
rect 31163 20964 31208 20992
rect 31202 20952 31208 20964
rect 31260 20952 31266 21004
rect 31757 20995 31815 21001
rect 31757 20961 31769 20995
rect 31803 20992 31815 20995
rect 31864 20992 31892 21032
rect 46198 21020 46204 21032
rect 46256 21020 46262 21072
rect 32122 20992 32128 21004
rect 31803 20964 31892 20992
rect 32083 20964 32128 20992
rect 31803 20961 31815 20964
rect 31757 20955 31815 20961
rect 32122 20952 32128 20964
rect 32180 20952 32186 21004
rect 35253 20995 35311 21001
rect 35253 20992 35265 20995
rect 32692 20964 35265 20992
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 8956 20788 8984 20887
rect 16850 20884 16856 20936
rect 16908 20924 16914 20936
rect 17129 20927 17187 20933
rect 17129 20924 17141 20927
rect 16908 20896 17141 20924
rect 16908 20884 16914 20896
rect 17129 20893 17141 20896
rect 17175 20893 17187 20927
rect 19242 20924 19248 20936
rect 19203 20896 19248 20924
rect 17129 20887 17187 20893
rect 19242 20884 19248 20896
rect 19300 20884 19306 20936
rect 20898 20884 20904 20936
rect 20956 20924 20962 20936
rect 21361 20927 21419 20933
rect 21361 20924 21373 20927
rect 20956 20896 21373 20924
rect 20956 20884 20962 20896
rect 21361 20893 21373 20896
rect 21407 20893 21419 20927
rect 21361 20887 21419 20893
rect 21637 20927 21695 20933
rect 21637 20893 21649 20927
rect 21683 20924 21695 20927
rect 22097 20927 22155 20933
rect 22097 20924 22109 20927
rect 21683 20896 22109 20924
rect 21683 20893 21695 20896
rect 21637 20887 21695 20893
rect 22097 20893 22109 20896
rect 22143 20893 22155 20927
rect 26694 20924 26700 20936
rect 26655 20896 26700 20924
rect 22097 20887 22155 20893
rect 26694 20884 26700 20896
rect 26752 20884 26758 20936
rect 27338 20884 27344 20936
rect 27396 20924 27402 20936
rect 27709 20927 27767 20933
rect 27709 20924 27721 20927
rect 27396 20896 27721 20924
rect 27396 20884 27402 20896
rect 27709 20893 27721 20896
rect 27755 20893 27767 20927
rect 27709 20887 27767 20893
rect 9122 20856 9128 20868
rect 9083 20828 9128 20856
rect 9122 20816 9128 20828
rect 9180 20816 9186 20868
rect 10778 20856 10784 20868
rect 10739 20828 10784 20856
rect 10778 20816 10784 20828
rect 10836 20816 10842 20868
rect 22373 20859 22431 20865
rect 22373 20825 22385 20859
rect 22419 20856 22431 20859
rect 22646 20856 22652 20868
rect 22419 20828 22652 20856
rect 22419 20825 22431 20828
rect 22373 20819 22431 20825
rect 22646 20816 22652 20828
rect 22704 20816 22710 20868
rect 23382 20816 23388 20868
rect 23440 20816 23446 20868
rect 30282 20816 30288 20868
rect 30340 20856 30346 20868
rect 30340 20828 30385 20856
rect 30340 20816 30346 20828
rect 31846 20816 31852 20868
rect 31904 20856 31910 20868
rect 31904 20828 31949 20856
rect 31904 20816 31910 20828
rect 9766 20788 9772 20800
rect 8956 20760 9772 20788
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 30190 20748 30196 20800
rect 30248 20788 30254 20800
rect 32692 20788 32720 20964
rect 35253 20961 35265 20964
rect 35299 20992 35311 20995
rect 35299 20964 41414 20992
rect 35299 20961 35311 20964
rect 35253 20955 35311 20961
rect 35894 20884 35900 20936
rect 35952 20924 35958 20936
rect 35952 20896 35997 20924
rect 35952 20884 35958 20896
rect 33778 20816 33784 20868
rect 33836 20856 33842 20868
rect 35345 20859 35403 20865
rect 35345 20856 35357 20859
rect 33836 20828 35357 20856
rect 33836 20816 33842 20828
rect 35345 20825 35357 20828
rect 35391 20856 35403 20859
rect 36354 20856 36360 20868
rect 35391 20828 36360 20856
rect 35391 20825 35403 20828
rect 35345 20819 35403 20825
rect 36354 20816 36360 20828
rect 36412 20816 36418 20868
rect 41386 20856 41414 20964
rect 42702 20952 42708 21004
rect 42760 20992 42766 21004
rect 43073 20995 43131 21001
rect 43073 20992 43085 20995
rect 42760 20964 43085 20992
rect 42760 20952 42766 20964
rect 43073 20961 43085 20964
rect 43119 20961 43131 20995
rect 43073 20955 43131 20961
rect 45189 20995 45247 21001
rect 45189 20961 45201 20995
rect 45235 20992 45247 20995
rect 46293 20995 46351 21001
rect 46293 20992 46305 20995
rect 45235 20964 46305 20992
rect 45235 20961 45247 20964
rect 45189 20955 45247 20961
rect 46293 20961 46305 20964
rect 46339 20961 46351 20995
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 46293 20955 46351 20961
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 42334 20884 42340 20936
rect 42392 20924 42398 20936
rect 43257 20927 43315 20933
rect 43257 20924 43269 20927
rect 42392 20896 43269 20924
rect 42392 20884 42398 20896
rect 43257 20893 43269 20896
rect 43303 20893 43315 20927
rect 43257 20887 43315 20893
rect 43441 20927 43499 20933
rect 43441 20893 43453 20927
rect 43487 20924 43499 20927
rect 43898 20924 43904 20936
rect 43487 20896 43904 20924
rect 43487 20893 43499 20896
rect 43441 20887 43499 20893
rect 43898 20884 43904 20896
rect 43956 20884 43962 20936
rect 44082 20924 44088 20936
rect 44043 20896 44088 20924
rect 44082 20884 44088 20896
rect 44140 20884 44146 20936
rect 45646 20924 45652 20936
rect 45607 20896 45652 20924
rect 45646 20884 45652 20896
rect 45704 20884 45710 20936
rect 45741 20859 45799 20865
rect 41386 20828 45554 20856
rect 43990 20788 43996 20800
rect 30248 20760 32720 20788
rect 43951 20760 43996 20788
rect 30248 20748 30254 20760
rect 43990 20748 43996 20760
rect 44048 20748 44054 20800
rect 45526 20788 45554 20828
rect 45741 20825 45753 20859
rect 45787 20856 45799 20859
rect 46477 20859 46535 20865
rect 46477 20856 46489 20859
rect 45787 20828 46489 20856
rect 45787 20825 45799 20828
rect 45741 20819 45799 20825
rect 46477 20825 46489 20828
rect 46523 20825 46535 20859
rect 46477 20819 46535 20825
rect 45922 20788 45928 20800
rect 45526 20760 45928 20788
rect 45922 20748 45928 20760
rect 45980 20748 45986 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 3050 20544 3056 20596
rect 3108 20584 3114 20596
rect 3108 20556 6914 20584
rect 3108 20544 3114 20556
rect 6886 20244 6914 20556
rect 10962 20544 10968 20596
rect 11020 20584 11026 20596
rect 13265 20587 13323 20593
rect 13265 20584 13277 20587
rect 11020 20556 13277 20584
rect 11020 20544 11026 20556
rect 13265 20553 13277 20556
rect 13311 20584 13323 20587
rect 13311 20556 13768 20584
rect 13311 20553 13323 20556
rect 13265 20547 13323 20553
rect 12802 20476 12808 20528
rect 12860 20476 12866 20528
rect 13740 20525 13768 20556
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 13909 20587 13967 20593
rect 13909 20584 13921 20587
rect 13872 20556 13921 20584
rect 13872 20544 13878 20556
rect 13909 20553 13921 20556
rect 13955 20584 13967 20587
rect 14182 20584 14188 20596
rect 13955 20556 14188 20584
rect 13955 20553 13967 20556
rect 13909 20547 13967 20553
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 14274 20544 14280 20596
rect 14332 20584 14338 20596
rect 14332 20556 14377 20584
rect 14332 20544 14338 20556
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 20089 20587 20147 20593
rect 20089 20584 20101 20587
rect 19392 20556 20101 20584
rect 19392 20544 19398 20556
rect 20089 20553 20101 20556
rect 20135 20584 20147 20587
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 20135 20556 21097 20584
rect 20135 20553 20147 20556
rect 20089 20547 20147 20553
rect 21085 20553 21097 20556
rect 21131 20584 21143 20587
rect 21266 20584 21272 20596
rect 21131 20556 21272 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 23293 20587 23351 20593
rect 23293 20553 23305 20587
rect 23339 20584 23351 20587
rect 23382 20584 23388 20596
rect 23339 20556 23388 20584
rect 23339 20553 23351 20556
rect 23293 20547 23351 20553
rect 23382 20544 23388 20556
rect 23440 20544 23446 20596
rect 28276 20556 31754 20584
rect 13725 20519 13783 20525
rect 13725 20485 13737 20519
rect 13771 20485 13783 20519
rect 13725 20479 13783 20485
rect 19889 20519 19947 20525
rect 19889 20485 19901 20519
rect 19935 20516 19947 20519
rect 20901 20519 20959 20525
rect 20901 20516 20913 20519
rect 19935 20488 20913 20516
rect 19935 20485 19947 20488
rect 19889 20479 19947 20485
rect 20901 20485 20913 20488
rect 20947 20516 20959 20519
rect 22094 20516 22100 20528
rect 20947 20488 22100 20516
rect 20947 20485 20959 20488
rect 20901 20479 20959 20485
rect 22094 20476 22100 20488
rect 22152 20476 22158 20528
rect 23842 20516 23848 20528
rect 22388 20488 23848 20516
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20448 10931 20451
rect 11330 20448 11336 20460
rect 10919 20420 11336 20448
rect 10919 20417 10931 20420
rect 10873 20411 10931 20417
rect 11330 20408 11336 20420
rect 11388 20408 11394 20460
rect 13998 20448 14004 20460
rect 13959 20420 14004 20448
rect 13998 20408 14004 20420
rect 14056 20408 14062 20460
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20448 14151 20451
rect 14458 20448 14464 20460
rect 14139 20420 14464 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 14458 20408 14464 20420
rect 14516 20408 14522 20460
rect 15105 20451 15163 20457
rect 15105 20417 15117 20451
rect 15151 20417 15163 20451
rect 15105 20411 15163 20417
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20448 15991 20451
rect 16850 20448 16856 20460
rect 15979 20420 16856 20448
rect 15979 20417 15991 20420
rect 15933 20411 15991 20417
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20380 11023 20383
rect 11517 20383 11575 20389
rect 11517 20380 11529 20383
rect 11011 20352 11529 20380
rect 11011 20349 11023 20352
rect 10965 20343 11023 20349
rect 11517 20349 11529 20352
rect 11563 20349 11575 20383
rect 11790 20380 11796 20392
rect 11751 20352 11796 20380
rect 11517 20343 11575 20349
rect 11790 20340 11796 20352
rect 11848 20340 11854 20392
rect 13538 20340 13544 20392
rect 13596 20380 13602 20392
rect 15120 20380 15148 20411
rect 16850 20408 16856 20420
rect 16908 20408 16914 20460
rect 17037 20451 17095 20457
rect 17037 20417 17049 20451
rect 17083 20417 17095 20451
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 17037 20411 17095 20417
rect 17236 20420 18061 20448
rect 17052 20380 17080 20411
rect 13596 20352 17080 20380
rect 13596 20340 13602 20352
rect 14090 20312 14096 20324
rect 12820 20284 14096 20312
rect 12820 20244 12848 20284
rect 14090 20272 14096 20284
rect 14148 20272 14154 20324
rect 17236 20321 17264 20420
rect 18049 20417 18061 20420
rect 18095 20448 18107 20451
rect 19242 20448 19248 20460
rect 18095 20420 19248 20448
rect 18095 20417 18107 20420
rect 18049 20411 18107 20417
rect 19242 20408 19248 20420
rect 19300 20408 19306 20460
rect 20806 20448 20812 20460
rect 20088 20420 20812 20448
rect 17221 20315 17279 20321
rect 17221 20281 17233 20315
rect 17267 20281 17279 20315
rect 17221 20275 17279 20281
rect 6886 20216 12848 20244
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 13136 20216 15301 20244
rect 13136 20204 13142 20216
rect 15289 20213 15301 20216
rect 15335 20244 15347 20247
rect 15654 20244 15660 20256
rect 15335 20216 15660 20244
rect 15335 20213 15347 20216
rect 15289 20207 15347 20213
rect 15654 20204 15660 20216
rect 15712 20204 15718 20256
rect 16025 20247 16083 20253
rect 16025 20213 16037 20247
rect 16071 20244 16083 20247
rect 16850 20244 16856 20256
rect 16071 20216 16856 20244
rect 16071 20213 16083 20216
rect 16025 20207 16083 20213
rect 16850 20204 16856 20216
rect 16908 20204 16914 20256
rect 18138 20244 18144 20256
rect 18099 20216 18144 20244
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18598 20204 18604 20256
rect 18656 20244 18662 20256
rect 20088 20253 20116 20420
rect 20806 20408 20812 20420
rect 20864 20448 20870 20460
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 20864 20420 21005 20448
rect 20864 20408 20870 20420
rect 20993 20417 21005 20420
rect 21039 20448 21051 20451
rect 21174 20448 21180 20460
rect 21039 20420 21180 20448
rect 21039 20417 21051 20420
rect 20993 20411 21051 20417
rect 21174 20408 21180 20420
rect 21232 20408 21238 20460
rect 22388 20457 22416 20488
rect 23842 20476 23848 20488
rect 23900 20476 23906 20528
rect 22373 20451 22431 20457
rect 22373 20417 22385 20451
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 23201 20451 23259 20457
rect 23201 20417 23213 20451
rect 23247 20417 23259 20451
rect 23201 20411 23259 20417
rect 21269 20383 21327 20389
rect 21269 20349 21281 20383
rect 21315 20380 21327 20383
rect 22281 20383 22339 20389
rect 22281 20380 22293 20383
rect 21315 20352 22293 20380
rect 21315 20349 21327 20352
rect 21269 20343 21327 20349
rect 22281 20349 22293 20352
rect 22327 20349 22339 20383
rect 22281 20343 22339 20349
rect 22646 20340 22652 20392
rect 22704 20380 22710 20392
rect 22741 20383 22799 20389
rect 22741 20380 22753 20383
rect 22704 20352 22753 20380
rect 22704 20340 22710 20352
rect 22741 20349 22753 20352
rect 22787 20349 22799 20383
rect 22741 20343 22799 20349
rect 20717 20315 20775 20321
rect 20717 20281 20729 20315
rect 20763 20312 20775 20315
rect 21726 20312 21732 20324
rect 20763 20284 21732 20312
rect 20763 20281 20775 20284
rect 20717 20275 20775 20281
rect 21726 20272 21732 20284
rect 21784 20272 21790 20324
rect 21818 20272 21824 20324
rect 21876 20312 21882 20324
rect 23216 20312 23244 20411
rect 23474 20408 23480 20460
rect 23532 20448 23538 20460
rect 24486 20448 24492 20460
rect 23532 20420 24492 20448
rect 23532 20408 23538 20420
rect 24486 20408 24492 20420
rect 24544 20448 24550 20460
rect 24857 20451 24915 20457
rect 24857 20448 24869 20451
rect 24544 20420 24869 20448
rect 24544 20408 24550 20420
rect 24857 20417 24869 20420
rect 24903 20417 24915 20451
rect 25774 20448 25780 20460
rect 25735 20420 25780 20448
rect 24857 20411 24915 20417
rect 25774 20408 25780 20420
rect 25832 20408 25838 20460
rect 26237 20451 26295 20457
rect 26237 20417 26249 20451
rect 26283 20448 26295 20451
rect 26973 20451 27031 20457
rect 26973 20448 26985 20451
rect 26283 20420 26985 20448
rect 26283 20417 26295 20420
rect 26237 20411 26295 20417
rect 26973 20417 26985 20420
rect 27019 20448 27031 20451
rect 27338 20448 27344 20460
rect 27019 20420 27344 20448
rect 27019 20417 27031 20420
rect 26973 20411 27031 20417
rect 27338 20408 27344 20420
rect 27396 20408 27402 20460
rect 27614 20408 27620 20460
rect 27672 20448 27678 20460
rect 28276 20457 28304 20556
rect 28353 20519 28411 20525
rect 28353 20485 28365 20519
rect 28399 20516 28411 20519
rect 29089 20519 29147 20525
rect 29089 20516 29101 20519
rect 28399 20488 29101 20516
rect 28399 20485 28411 20488
rect 28353 20479 28411 20485
rect 29089 20485 29101 20488
rect 29135 20485 29147 20519
rect 29089 20479 29147 20485
rect 30282 20476 30288 20528
rect 30340 20516 30346 20528
rect 31726 20516 31754 20556
rect 32306 20544 32312 20596
rect 32364 20584 32370 20596
rect 32585 20587 32643 20593
rect 32585 20584 32597 20587
rect 32364 20556 32597 20584
rect 32364 20544 32370 20556
rect 32585 20553 32597 20556
rect 32631 20553 32643 20587
rect 32585 20547 32643 20553
rect 42521 20587 42579 20593
rect 42521 20553 42533 20587
rect 42567 20584 42579 20587
rect 44082 20584 44088 20596
rect 42567 20556 44088 20584
rect 42567 20553 42579 20556
rect 42521 20547 42579 20553
rect 44082 20544 44088 20556
rect 44140 20544 44146 20596
rect 44177 20587 44235 20593
rect 44177 20553 44189 20587
rect 44223 20584 44235 20587
rect 46474 20584 46480 20596
rect 44223 20556 46480 20584
rect 44223 20553 44235 20556
rect 44177 20547 44235 20553
rect 46474 20544 46480 20556
rect 46532 20544 46538 20596
rect 48038 20584 48044 20596
rect 47999 20556 48044 20584
rect 48038 20544 48044 20556
rect 48096 20544 48102 20596
rect 45554 20516 45560 20528
rect 30340 20488 31340 20516
rect 31726 20488 45560 20516
rect 30340 20476 30346 20488
rect 28261 20451 28319 20457
rect 28261 20448 28273 20451
rect 27672 20420 28273 20448
rect 27672 20408 27678 20420
rect 28261 20417 28273 20420
rect 28307 20417 28319 20451
rect 31202 20448 31208 20460
rect 31163 20420 31208 20448
rect 28261 20411 28319 20417
rect 31202 20408 31208 20420
rect 31260 20408 31266 20460
rect 31312 20448 31340 20488
rect 45554 20476 45560 20488
rect 45612 20476 45618 20528
rect 32125 20451 32183 20457
rect 32125 20448 32137 20451
rect 31312 20420 32137 20448
rect 32125 20417 32137 20420
rect 32171 20417 32183 20451
rect 32125 20411 32183 20417
rect 42334 20408 42340 20460
rect 42392 20448 42398 20460
rect 42429 20451 42487 20457
rect 42429 20448 42441 20451
rect 42392 20420 42441 20448
rect 42392 20408 42398 20420
rect 42429 20417 42441 20420
rect 42475 20417 42487 20451
rect 42429 20411 42487 20417
rect 42613 20451 42671 20457
rect 42613 20417 42625 20451
rect 42659 20448 42671 20451
rect 42702 20448 42708 20460
rect 42659 20420 42708 20448
rect 42659 20417 42671 20420
rect 42613 20411 42671 20417
rect 42702 20408 42708 20420
rect 42760 20408 42766 20460
rect 43346 20408 43352 20460
rect 43404 20448 43410 20460
rect 43441 20451 43499 20457
rect 43441 20448 43453 20451
rect 43404 20420 43453 20448
rect 43404 20408 43410 20420
rect 43441 20417 43453 20420
rect 43487 20448 43499 20451
rect 43990 20448 43996 20460
rect 43487 20420 43996 20448
rect 43487 20417 43499 20420
rect 43441 20411 43499 20417
rect 43990 20408 43996 20420
rect 44048 20408 44054 20460
rect 44634 20448 44640 20460
rect 44595 20420 44640 20448
rect 44634 20408 44640 20420
rect 44692 20408 44698 20460
rect 47581 20451 47639 20457
rect 47581 20417 47593 20451
rect 47627 20448 47639 20451
rect 47946 20448 47952 20460
rect 47627 20420 47952 20448
rect 47627 20417 47639 20420
rect 47581 20411 47639 20417
rect 47946 20408 47952 20420
rect 48004 20408 48010 20460
rect 28905 20383 28963 20389
rect 28905 20349 28917 20383
rect 28951 20380 28963 20383
rect 29914 20380 29920 20392
rect 28951 20352 29920 20380
rect 28951 20349 28963 20352
rect 28905 20343 28963 20349
rect 29914 20340 29920 20352
rect 29972 20340 29978 20392
rect 30006 20340 30012 20392
rect 30064 20380 30070 20392
rect 31220 20380 31248 20408
rect 41046 20380 41052 20392
rect 30064 20352 30109 20380
rect 31220 20352 41052 20380
rect 30064 20340 30070 20352
rect 41046 20340 41052 20352
rect 41104 20340 41110 20392
rect 43530 20380 43536 20392
rect 43491 20352 43536 20380
rect 43530 20340 43536 20352
rect 43588 20340 43594 20392
rect 44821 20383 44879 20389
rect 44821 20349 44833 20383
rect 44867 20380 44879 20383
rect 45186 20380 45192 20392
rect 44867 20352 45192 20380
rect 44867 20349 44879 20352
rect 44821 20343 44879 20349
rect 45186 20340 45192 20352
rect 45244 20340 45250 20392
rect 46014 20380 46020 20392
rect 45975 20352 46020 20380
rect 46014 20340 46020 20352
rect 46072 20340 46078 20392
rect 21876 20284 23244 20312
rect 21876 20272 21882 20284
rect 24578 20272 24584 20324
rect 24636 20312 24642 20324
rect 27154 20312 27160 20324
rect 24636 20284 27160 20312
rect 24636 20272 24642 20284
rect 27154 20272 27160 20284
rect 27212 20272 27218 20324
rect 20073 20247 20131 20253
rect 20073 20244 20085 20247
rect 18656 20216 20085 20244
rect 18656 20204 18662 20216
rect 20073 20213 20085 20216
rect 20119 20213 20131 20247
rect 20254 20244 20260 20256
rect 20215 20216 20260 20244
rect 20073 20207 20131 20213
rect 20254 20204 20260 20216
rect 20312 20204 20318 20256
rect 25041 20247 25099 20253
rect 25041 20213 25053 20247
rect 25087 20244 25099 20247
rect 25222 20244 25228 20256
rect 25087 20216 25228 20244
rect 25087 20213 25099 20216
rect 25041 20207 25099 20213
rect 25222 20204 25228 20216
rect 25280 20204 25286 20256
rect 25498 20204 25504 20256
rect 25556 20244 25562 20256
rect 25593 20247 25651 20253
rect 25593 20244 25605 20247
rect 25556 20216 25605 20244
rect 25556 20204 25562 20216
rect 25593 20213 25605 20216
rect 25639 20213 25651 20247
rect 25593 20207 25651 20213
rect 26234 20204 26240 20256
rect 26292 20244 26298 20256
rect 26329 20247 26387 20253
rect 26329 20244 26341 20247
rect 26292 20216 26341 20244
rect 26292 20204 26298 20216
rect 26329 20213 26341 20216
rect 26375 20213 26387 20247
rect 27062 20244 27068 20256
rect 27023 20216 27068 20244
rect 26329 20207 26387 20213
rect 27062 20204 27068 20216
rect 27120 20204 27126 20256
rect 30190 20204 30196 20256
rect 30248 20244 30254 20256
rect 31297 20247 31355 20253
rect 31297 20244 31309 20247
rect 30248 20216 31309 20244
rect 30248 20204 30254 20216
rect 31297 20213 31309 20216
rect 31343 20213 31355 20247
rect 32306 20244 32312 20256
rect 32267 20216 32312 20244
rect 31297 20207 31355 20213
rect 32306 20204 32312 20216
rect 32364 20204 32370 20256
rect 47210 20204 47216 20256
rect 47268 20244 47274 20256
rect 47673 20247 47731 20253
rect 47673 20244 47685 20247
rect 47268 20216 47685 20244
rect 47268 20204 47274 20216
rect 47673 20213 47685 20216
rect 47719 20213 47731 20247
rect 47673 20207 47731 20213
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 3510 20000 3516 20052
rect 3568 20040 3574 20052
rect 30006 20040 30012 20052
rect 3568 20012 30012 20040
rect 3568 20000 3574 20012
rect 30006 20000 30012 20012
rect 30064 20000 30070 20052
rect 45186 20040 45192 20052
rect 45147 20012 45192 20040
rect 45186 20000 45192 20012
rect 45244 20000 45250 20052
rect 11517 19975 11575 19981
rect 11517 19941 11529 19975
rect 11563 19972 11575 19975
rect 11790 19972 11796 19984
rect 11563 19944 11796 19972
rect 11563 19941 11575 19944
rect 11517 19935 11575 19941
rect 11790 19932 11796 19944
rect 11848 19932 11854 19984
rect 12802 19972 12808 19984
rect 12763 19944 12808 19972
rect 12802 19932 12808 19944
rect 12860 19932 12866 19984
rect 21726 19972 21732 19984
rect 21687 19944 21732 19972
rect 21726 19932 21732 19944
rect 21784 19932 21790 19984
rect 43806 19972 43812 19984
rect 43767 19944 43812 19972
rect 43806 19932 43812 19944
rect 43864 19932 43870 19984
rect 46474 19972 46480 19984
rect 46216 19944 46480 19972
rect 10962 19864 10968 19916
rect 11020 19904 11026 19916
rect 11020 19876 12204 19904
rect 11020 19864 11026 19876
rect 11701 19839 11759 19845
rect 11701 19805 11713 19839
rect 11747 19836 11759 19839
rect 11882 19836 11888 19848
rect 11747 19808 11888 19836
rect 11747 19805 11759 19808
rect 11701 19799 11759 19805
rect 11882 19796 11888 19808
rect 11940 19796 11946 19848
rect 12176 19845 12204 19876
rect 12342 19864 12348 19916
rect 12400 19904 12406 19916
rect 16850 19904 16856 19916
rect 12400 19876 13400 19904
rect 16811 19876 16856 19904
rect 12400 19864 12406 19876
rect 11977 19839 12035 19845
rect 11977 19805 11989 19839
rect 12023 19805 12035 19839
rect 11977 19799 12035 19805
rect 12161 19839 12219 19845
rect 12161 19805 12173 19839
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12713 19839 12771 19845
rect 12713 19805 12725 19839
rect 12759 19836 12771 19839
rect 13078 19836 13084 19848
rect 12759 19808 13084 19836
rect 12759 19805 12771 19808
rect 12713 19799 12771 19805
rect 11992 19768 12020 19799
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13372 19845 13400 19876
rect 16850 19864 16856 19876
rect 16908 19864 16914 19916
rect 17129 19907 17187 19913
rect 17129 19873 17141 19907
rect 17175 19904 17187 19907
rect 18322 19904 18328 19916
rect 17175 19876 18328 19904
rect 17175 19873 17187 19876
rect 17129 19867 17187 19873
rect 18322 19864 18328 19876
rect 18380 19864 18386 19916
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 20990 19904 20996 19916
rect 19484 19876 20996 19904
rect 19484 19864 19490 19876
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 25222 19904 25228 19916
rect 25183 19876 25228 19904
rect 25222 19864 25228 19876
rect 25280 19864 25286 19916
rect 25498 19904 25504 19916
rect 25459 19876 25504 19904
rect 25498 19864 25504 19876
rect 25556 19864 25562 19916
rect 30190 19904 30196 19916
rect 30151 19876 30196 19904
rect 30190 19864 30196 19876
rect 30248 19864 30254 19916
rect 31662 19904 31668 19916
rect 31623 19876 31668 19904
rect 31662 19864 31668 19876
rect 31720 19864 31726 19916
rect 43346 19904 43352 19916
rect 43307 19876 43352 19904
rect 43346 19864 43352 19876
rect 43404 19864 43410 19916
rect 43898 19904 43904 19916
rect 43859 19876 43904 19904
rect 43898 19864 43904 19876
rect 43956 19864 43962 19916
rect 46216 19913 46244 19944
rect 46474 19932 46480 19944
rect 46532 19932 46538 19984
rect 46201 19907 46259 19913
rect 46201 19873 46213 19907
rect 46247 19873 46259 19907
rect 46382 19904 46388 19916
rect 46343 19876 46388 19904
rect 46201 19867 46259 19873
rect 46382 19864 46388 19876
rect 46440 19864 46446 19916
rect 46842 19864 46848 19916
rect 46900 19904 46906 19916
rect 46937 19907 46995 19913
rect 46937 19904 46949 19907
rect 46900 19876 46949 19904
rect 46900 19864 46906 19876
rect 46937 19873 46949 19876
rect 46983 19873 46995 19907
rect 46937 19867 46995 19873
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19805 13415 19839
rect 13357 19799 13415 19805
rect 13449 19839 13507 19845
rect 13449 19805 13461 19839
rect 13495 19836 13507 19839
rect 14461 19839 14519 19845
rect 14461 19836 14473 19839
rect 13495 19808 14473 19836
rect 13495 19805 13507 19808
rect 13449 19799 13507 19805
rect 14461 19805 14473 19808
rect 14507 19805 14519 19839
rect 19978 19836 19984 19848
rect 19939 19808 19984 19836
rect 14461 19799 14519 19805
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 24486 19836 24492 19848
rect 24447 19808 24492 19836
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 27154 19796 27160 19848
rect 27212 19836 27218 19848
rect 30009 19839 30067 19845
rect 30009 19836 30021 19839
rect 27212 19808 30021 19836
rect 27212 19796 27218 19808
rect 30009 19805 30021 19808
rect 30055 19805 30067 19839
rect 30009 19799 30067 19805
rect 42426 19796 42432 19848
rect 42484 19836 42490 19848
rect 43073 19839 43131 19845
rect 43073 19836 43085 19839
rect 42484 19808 43085 19836
rect 42484 19796 42490 19808
rect 43073 19805 43085 19808
rect 43119 19805 43131 19839
rect 43073 19799 43131 19805
rect 43625 19839 43683 19845
rect 43625 19805 43637 19839
rect 43671 19836 43683 19839
rect 43671 19808 43944 19836
rect 43671 19805 43683 19808
rect 43625 19799 43683 19805
rect 43916 19780 43944 19808
rect 44818 19796 44824 19848
rect 44876 19836 44882 19848
rect 45097 19839 45155 19845
rect 45097 19836 45109 19839
rect 44876 19808 45109 19836
rect 44876 19796 44882 19808
rect 45097 19805 45109 19808
rect 45143 19836 45155 19839
rect 45830 19836 45836 19848
rect 45143 19808 45836 19836
rect 45143 19805 45155 19808
rect 45097 19799 45155 19805
rect 45830 19796 45836 19808
rect 45888 19796 45894 19848
rect 13722 19768 13728 19780
rect 11992 19740 13728 19768
rect 13722 19728 13728 19740
rect 13780 19728 13786 19780
rect 14090 19728 14096 19780
rect 14148 19768 14154 19780
rect 14737 19771 14795 19777
rect 14737 19768 14749 19771
rect 14148 19740 14749 19768
rect 14148 19728 14154 19740
rect 14737 19737 14749 19740
rect 14783 19737 14795 19771
rect 14737 19731 14795 19737
rect 15746 19728 15752 19780
rect 15804 19728 15810 19780
rect 18138 19728 18144 19780
rect 18196 19728 18202 19780
rect 20257 19771 20315 19777
rect 20257 19737 20269 19771
rect 20303 19768 20315 19771
rect 20530 19768 20536 19780
rect 20303 19740 20536 19768
rect 20303 19737 20315 19740
rect 20257 19731 20315 19737
rect 20530 19728 20536 19740
rect 20588 19728 20594 19780
rect 21910 19768 21916 19780
rect 21482 19740 21916 19768
rect 21910 19728 21916 19740
rect 21968 19728 21974 19780
rect 24765 19771 24823 19777
rect 24765 19737 24777 19771
rect 24811 19768 24823 19771
rect 25406 19768 25412 19780
rect 24811 19740 25412 19768
rect 24811 19737 24823 19740
rect 24765 19731 24823 19737
rect 25406 19728 25412 19740
rect 25464 19728 25470 19780
rect 26234 19728 26240 19780
rect 26292 19728 26298 19780
rect 43898 19728 43904 19780
rect 43956 19728 43962 19780
rect 13998 19660 14004 19712
rect 14056 19700 14062 19712
rect 14826 19700 14832 19712
rect 14056 19672 14832 19700
rect 14056 19660 14062 19672
rect 14826 19660 14832 19672
rect 14884 19700 14890 19712
rect 16209 19703 16267 19709
rect 16209 19700 16221 19703
rect 14884 19672 16221 19700
rect 14884 19660 14890 19672
rect 16209 19669 16221 19672
rect 16255 19700 16267 19703
rect 16298 19700 16304 19712
rect 16255 19672 16304 19700
rect 16255 19669 16267 19672
rect 16209 19663 16267 19669
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 18598 19700 18604 19712
rect 18559 19672 18604 19700
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 19242 19660 19248 19712
rect 19300 19700 19306 19712
rect 21818 19700 21824 19712
rect 19300 19672 21824 19700
rect 19300 19660 19306 19672
rect 21818 19660 21824 19672
rect 21876 19660 21882 19712
rect 23290 19660 23296 19712
rect 23348 19700 23354 19712
rect 26973 19703 27031 19709
rect 26973 19700 26985 19703
rect 23348 19672 26985 19700
rect 23348 19660 23354 19672
rect 26973 19669 26985 19672
rect 27019 19700 27031 19703
rect 35986 19700 35992 19712
rect 27019 19672 35992 19700
rect 27019 19669 27031 19672
rect 26973 19663 27031 19669
rect 35986 19660 35992 19672
rect 36044 19660 36050 19712
rect 45922 19660 45928 19712
rect 45980 19700 45986 19712
rect 47670 19700 47676 19712
rect 45980 19672 47676 19700
rect 45980 19660 45986 19672
rect 47670 19660 47676 19672
rect 47728 19660 47734 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 1670 19456 1676 19508
rect 1728 19496 1734 19508
rect 23937 19499 23995 19505
rect 1728 19468 22094 19496
rect 1728 19456 1734 19468
rect 2225 19431 2283 19437
rect 2225 19397 2237 19431
rect 2271 19428 2283 19431
rect 3050 19428 3056 19440
rect 2271 19400 3056 19428
rect 2271 19397 2283 19400
rect 2225 19391 2283 19397
rect 3050 19388 3056 19400
rect 3108 19388 3114 19440
rect 13814 19428 13820 19440
rect 13775 19400 13820 19428
rect 13814 19388 13820 19400
rect 13872 19388 13878 19440
rect 13998 19428 14004 19440
rect 13959 19400 14004 19428
rect 13998 19388 14004 19400
rect 14056 19388 14062 19440
rect 14093 19431 14151 19437
rect 14093 19397 14105 19431
rect 14139 19428 14151 19431
rect 14458 19428 14464 19440
rect 14139 19400 14464 19428
rect 14139 19397 14151 19400
rect 14093 19391 14151 19397
rect 14458 19388 14464 19400
rect 14516 19388 14522 19440
rect 14826 19428 14832 19440
rect 14787 19400 14832 19428
rect 14826 19388 14832 19400
rect 14884 19388 14890 19440
rect 15010 19388 15016 19440
rect 15068 19437 15074 19440
rect 15068 19431 15087 19437
rect 15075 19397 15087 19431
rect 15746 19428 15752 19440
rect 15707 19400 15752 19428
rect 15068 19391 15087 19397
rect 15068 19388 15074 19391
rect 15746 19388 15752 19400
rect 15804 19388 15810 19440
rect 17037 19431 17095 19437
rect 17037 19397 17049 19431
rect 17083 19428 17095 19431
rect 18506 19428 18512 19440
rect 17083 19400 18512 19428
rect 17083 19397 17095 19400
rect 17037 19391 17095 19397
rect 18506 19388 18512 19400
rect 18564 19428 18570 19440
rect 19058 19428 19064 19440
rect 18564 19400 19064 19428
rect 18564 19388 18570 19400
rect 19058 19388 19064 19400
rect 19116 19388 19122 19440
rect 19521 19431 19579 19437
rect 19521 19397 19533 19431
rect 19567 19428 19579 19431
rect 19978 19428 19984 19440
rect 19567 19400 19984 19428
rect 19567 19397 19579 19400
rect 19521 19391 19579 19397
rect 19978 19388 19984 19400
rect 20036 19388 20042 19440
rect 21726 19428 21732 19440
rect 20180 19400 21732 19428
rect 11330 19320 11336 19372
rect 11388 19360 11394 19372
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 11388 19332 11897 19360
rect 11388 19320 11394 19332
rect 11885 19329 11897 19332
rect 11931 19360 11943 19363
rect 12342 19360 12348 19372
rect 11931 19332 12348 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 12342 19320 12348 19332
rect 12400 19320 12406 19372
rect 12989 19363 13047 19369
rect 12989 19329 13001 19363
rect 13035 19360 13047 19363
rect 13832 19360 13860 19388
rect 13035 19332 13860 19360
rect 14185 19363 14243 19369
rect 13035 19329 13047 19332
rect 12989 19323 13047 19329
rect 14185 19329 14197 19363
rect 14231 19360 14243 19363
rect 15028 19360 15056 19388
rect 15654 19360 15660 19372
rect 14231 19332 15056 19360
rect 15615 19332 15660 19360
rect 14231 19329 14243 19332
rect 14185 19323 14243 19329
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 16574 19320 16580 19372
rect 16632 19360 16638 19372
rect 16761 19363 16819 19369
rect 16761 19360 16773 19363
rect 16632 19332 16773 19360
rect 16632 19320 16638 19332
rect 16761 19329 16773 19332
rect 16807 19329 16819 19363
rect 16761 19323 16819 19329
rect 17957 19363 18015 19369
rect 17957 19329 17969 19363
rect 18003 19360 18015 19363
rect 18598 19360 18604 19372
rect 18003 19332 18604 19360
rect 18003 19329 18015 19332
rect 17957 19323 18015 19329
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 19426 19360 19432 19372
rect 19387 19332 19432 19360
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 20180 19369 20208 19400
rect 21726 19388 21732 19400
rect 21784 19388 21790 19440
rect 21910 19428 21916 19440
rect 21871 19400 21916 19428
rect 21910 19388 21916 19400
rect 21968 19388 21974 19440
rect 22066 19428 22094 19468
rect 23937 19465 23949 19499
rect 23983 19496 23995 19499
rect 25774 19496 25780 19508
rect 23983 19468 25780 19496
rect 23983 19465 23995 19468
rect 23937 19459 23995 19465
rect 25774 19456 25780 19468
rect 25832 19456 25838 19508
rect 27985 19499 28043 19505
rect 27985 19465 27997 19499
rect 28031 19496 28043 19499
rect 28258 19496 28264 19508
rect 28031 19468 28264 19496
rect 28031 19465 28043 19468
rect 27985 19459 28043 19465
rect 28258 19456 28264 19468
rect 28316 19496 28322 19508
rect 28718 19496 28724 19508
rect 28316 19468 28724 19496
rect 28316 19456 28322 19468
rect 28718 19456 28724 19468
rect 28776 19496 28782 19508
rect 28905 19499 28963 19505
rect 28905 19496 28917 19499
rect 28776 19468 28917 19496
rect 28776 19456 28782 19468
rect 28905 19465 28917 19468
rect 28951 19465 28963 19499
rect 29914 19496 29920 19508
rect 29875 19468 29920 19496
rect 28905 19459 28963 19465
rect 29914 19456 29920 19468
rect 29972 19456 29978 19508
rect 43530 19496 43536 19508
rect 43491 19468 43536 19496
rect 43530 19456 43536 19468
rect 43588 19456 43594 19508
rect 47765 19499 47823 19505
rect 47765 19496 47777 19499
rect 46676 19468 47777 19496
rect 45554 19428 45560 19440
rect 22066 19400 45560 19428
rect 45554 19388 45560 19400
rect 45612 19428 45618 19440
rect 45612 19400 46520 19428
rect 45612 19388 45618 19400
rect 20165 19363 20223 19369
rect 20165 19329 20177 19363
rect 20211 19329 20223 19363
rect 20165 19323 20223 19329
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19329 21051 19363
rect 21174 19360 21180 19372
rect 21135 19332 21180 19360
rect 20993 19323 21051 19329
rect 2038 19292 2044 19304
rect 1999 19264 2044 19292
rect 2038 19252 2044 19264
rect 2096 19252 2102 19304
rect 2774 19292 2780 19304
rect 2735 19264 2780 19292
rect 2774 19252 2780 19264
rect 2832 19252 2838 19304
rect 13081 19295 13139 19301
rect 13081 19261 13093 19295
rect 13127 19292 13139 19295
rect 14274 19292 14280 19304
rect 13127 19264 14280 19292
rect 13127 19261 13139 19264
rect 13081 19255 13139 19261
rect 14274 19252 14280 19264
rect 14332 19252 14338 19304
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19261 18107 19295
rect 18322 19292 18328 19304
rect 18283 19264 18328 19292
rect 18049 19255 18107 19261
rect 14292 19224 14320 19252
rect 15197 19227 15255 19233
rect 15197 19224 15209 19227
rect 14292 19196 15209 19224
rect 15197 19193 15209 19196
rect 15243 19193 15255 19227
rect 18064 19224 18092 19255
rect 18322 19252 18328 19264
rect 18380 19252 18386 19304
rect 20254 19292 20260 19304
rect 20215 19264 20260 19292
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 20530 19292 20536 19304
rect 20491 19264 20536 19292
rect 20530 19252 20536 19264
rect 20588 19252 20594 19304
rect 21008 19292 21036 19323
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 21266 19320 21272 19372
rect 21324 19360 21330 19372
rect 21818 19360 21824 19372
rect 21324 19332 21369 19360
rect 21779 19332 21824 19360
rect 21324 19320 21330 19332
rect 21818 19320 21824 19332
rect 21876 19360 21882 19372
rect 22465 19363 22523 19369
rect 22465 19360 22477 19363
rect 21876 19332 22477 19360
rect 21876 19320 21882 19332
rect 22465 19329 22477 19332
rect 22511 19329 22523 19363
rect 23750 19360 23756 19372
rect 23711 19332 23756 19360
rect 22465 19323 22523 19329
rect 23750 19320 23756 19332
rect 23808 19320 23814 19372
rect 24578 19360 24584 19372
rect 24539 19332 24584 19360
rect 24578 19320 24584 19332
rect 24636 19320 24642 19372
rect 25415 19363 25473 19369
rect 25415 19329 25427 19363
rect 25461 19329 25473 19363
rect 25590 19360 25596 19372
rect 25551 19332 25596 19360
rect 25415 19323 25473 19329
rect 22094 19292 22100 19304
rect 21008 19264 22100 19292
rect 22094 19252 22100 19264
rect 22152 19292 22158 19304
rect 22554 19292 22560 19304
rect 22152 19264 22560 19292
rect 22152 19252 22158 19264
rect 22554 19252 22560 19264
rect 22612 19252 22618 19304
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19292 23627 19295
rect 24673 19295 24731 19301
rect 24673 19292 24685 19295
rect 23615 19264 24685 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 24673 19261 24685 19264
rect 24719 19292 24731 19295
rect 25038 19292 25044 19304
rect 24719 19264 25044 19292
rect 24719 19261 24731 19264
rect 24673 19255 24731 19261
rect 25038 19252 25044 19264
rect 25096 19252 25102 19304
rect 19334 19224 19340 19236
rect 18064 19196 19340 19224
rect 15197 19187 15255 19193
rect 19334 19184 19340 19196
rect 19392 19184 19398 19236
rect 24394 19184 24400 19236
rect 24452 19224 24458 19236
rect 25424 19224 25452 19323
rect 25590 19320 25596 19332
rect 25648 19320 25654 19372
rect 28258 19360 28264 19372
rect 28219 19332 28264 19360
rect 28258 19320 28264 19332
rect 28316 19320 28322 19372
rect 28445 19363 28503 19369
rect 28445 19329 28457 19363
rect 28491 19360 28503 19363
rect 28902 19360 28908 19372
rect 28491 19332 28908 19360
rect 28491 19329 28503 19332
rect 28445 19323 28503 19329
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 29273 19363 29331 19369
rect 29273 19360 29285 19363
rect 29012 19332 29285 19360
rect 28629 19295 28687 19301
rect 28629 19261 28641 19295
rect 28675 19292 28687 19295
rect 29012 19292 29040 19332
rect 29273 19329 29285 19332
rect 29319 19329 29331 19363
rect 29273 19323 29331 19329
rect 29457 19363 29515 19369
rect 29457 19329 29469 19363
rect 29503 19360 29515 19363
rect 30101 19363 30159 19369
rect 30101 19360 30113 19363
rect 29503 19332 30113 19360
rect 29503 19329 29515 19332
rect 29457 19323 29515 19329
rect 30101 19329 30113 19332
rect 30147 19329 30159 19363
rect 30101 19323 30159 19329
rect 42426 19320 42432 19372
rect 42484 19360 42490 19372
rect 43349 19363 43407 19369
rect 43349 19360 43361 19363
rect 42484 19332 43361 19360
rect 42484 19320 42490 19332
rect 43349 19329 43361 19332
rect 43395 19329 43407 19363
rect 43349 19323 43407 19329
rect 43533 19363 43591 19369
rect 43533 19329 43545 19363
rect 43579 19360 43591 19363
rect 43898 19360 43904 19372
rect 43579 19332 43904 19360
rect 43579 19329 43591 19332
rect 43533 19323 43591 19329
rect 43898 19320 43904 19332
rect 43956 19320 43962 19372
rect 45922 19360 45928 19372
rect 45883 19332 45928 19360
rect 45922 19320 45928 19332
rect 45980 19320 45986 19372
rect 46492 19369 46520 19400
rect 46676 19369 46704 19468
rect 47765 19465 47777 19468
rect 47811 19496 47823 19499
rect 47946 19496 47952 19508
rect 47811 19468 47952 19496
rect 47811 19465 47823 19468
rect 47765 19459 47823 19465
rect 47946 19456 47952 19468
rect 48004 19456 48010 19508
rect 48038 19456 48044 19508
rect 48096 19496 48102 19508
rect 48133 19499 48191 19505
rect 48133 19496 48145 19499
rect 48096 19468 48145 19496
rect 48096 19456 48102 19468
rect 48133 19465 48145 19468
rect 48179 19465 48191 19499
rect 48133 19459 48191 19465
rect 47857 19431 47915 19437
rect 47857 19428 47869 19431
rect 46768 19400 47869 19428
rect 46477 19363 46535 19369
rect 46477 19329 46489 19363
rect 46523 19360 46535 19363
rect 46661 19363 46719 19369
rect 46523 19332 46612 19360
rect 46523 19329 46535 19332
rect 46477 19323 46535 19329
rect 28675 19264 29040 19292
rect 28675 19261 28687 19264
rect 28629 19255 28687 19261
rect 29086 19252 29092 19304
rect 29144 19292 29150 19304
rect 46584 19292 46612 19332
rect 46661 19329 46673 19363
rect 46707 19329 46719 19363
rect 46661 19323 46719 19329
rect 46768 19292 46796 19400
rect 47857 19397 47869 19400
rect 47903 19397 47915 19431
rect 47857 19391 47915 19397
rect 46845 19363 46903 19369
rect 46845 19329 46857 19363
rect 46891 19360 46903 19363
rect 46891 19332 47624 19360
rect 46891 19329 46903 19332
rect 46845 19323 46903 19329
rect 29144 19264 29189 19292
rect 46584 19264 46796 19292
rect 29144 19252 29150 19264
rect 47596 19233 47624 19332
rect 47670 19320 47676 19372
rect 47728 19360 47734 19372
rect 47949 19363 48007 19369
rect 47949 19360 47961 19363
rect 47728 19332 47961 19360
rect 47728 19320 47734 19332
rect 47949 19329 47961 19332
rect 47995 19329 48007 19363
rect 47949 19323 48007 19329
rect 24452 19196 25452 19224
rect 47581 19227 47639 19233
rect 24452 19184 24458 19196
rect 47581 19193 47593 19227
rect 47627 19224 47639 19227
rect 47854 19224 47860 19236
rect 47627 19196 47860 19224
rect 47627 19193 47639 19196
rect 47581 19187 47639 19193
rect 47854 19184 47860 19196
rect 47912 19184 47918 19236
rect 11790 19116 11796 19168
rect 11848 19156 11854 19168
rect 11885 19159 11943 19165
rect 11885 19156 11897 19159
rect 11848 19128 11897 19156
rect 11848 19116 11854 19128
rect 11885 19125 11897 19128
rect 11931 19125 11943 19159
rect 11885 19119 11943 19125
rect 12066 19116 12072 19168
rect 12124 19156 12130 19168
rect 13357 19159 13415 19165
rect 13357 19156 13369 19159
rect 12124 19128 13369 19156
rect 12124 19116 12130 19128
rect 13357 19125 13369 19128
rect 13403 19125 13415 19159
rect 13357 19119 13415 19125
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 14369 19159 14427 19165
rect 14369 19156 14381 19159
rect 13780 19128 14381 19156
rect 13780 19116 13786 19128
rect 14369 19125 14381 19128
rect 14415 19125 14427 19159
rect 14369 19119 14427 19125
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 15013 19159 15071 19165
rect 15013 19156 15025 19159
rect 14516 19128 15025 19156
rect 14516 19116 14522 19128
rect 15013 19125 15025 19128
rect 15059 19156 15071 19159
rect 15102 19156 15108 19168
rect 15059 19128 15108 19156
rect 15059 19125 15071 19128
rect 15013 19119 15071 19125
rect 15102 19116 15108 19128
rect 15160 19116 15166 19168
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 20993 19159 21051 19165
rect 20993 19156 21005 19159
rect 20772 19128 21005 19156
rect 20772 19116 20778 19128
rect 20993 19125 21005 19128
rect 21039 19125 21051 19159
rect 20993 19119 21051 19125
rect 22370 19116 22376 19168
rect 22428 19156 22434 19168
rect 22557 19159 22615 19165
rect 22557 19156 22569 19159
rect 22428 19128 22569 19156
rect 22428 19116 22434 19128
rect 22557 19125 22569 19128
rect 22603 19125 22615 19159
rect 24854 19156 24860 19168
rect 24815 19128 24860 19156
rect 22557 19119 22615 19125
rect 24854 19116 24860 19128
rect 24912 19116 24918 19168
rect 25038 19116 25044 19168
rect 25096 19156 25102 19168
rect 25501 19159 25559 19165
rect 25501 19156 25513 19159
rect 25096 19128 25513 19156
rect 25096 19116 25102 19128
rect 25501 19125 25513 19128
rect 25547 19125 25559 19159
rect 45462 19156 45468 19168
rect 45423 19128 45468 19156
rect 25501 19119 25559 19125
rect 45462 19116 45468 19128
rect 45520 19116 45526 19168
rect 46198 19156 46204 19168
rect 46159 19128 46204 19156
rect 46198 19116 46204 19128
rect 46256 19116 46262 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 2038 18912 2044 18964
rect 2096 18952 2102 18964
rect 2317 18955 2375 18961
rect 2317 18952 2329 18955
rect 2096 18924 2329 18952
rect 2096 18912 2102 18924
rect 2317 18921 2329 18924
rect 2363 18921 2375 18955
rect 3050 18952 3056 18964
rect 3011 18924 3056 18952
rect 2317 18915 2375 18921
rect 3050 18912 3056 18924
rect 3108 18912 3114 18964
rect 13541 18955 13599 18961
rect 13541 18921 13553 18955
rect 13587 18952 13599 18955
rect 13814 18952 13820 18964
rect 13587 18924 13820 18952
rect 13587 18921 13599 18924
rect 13541 18915 13599 18921
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 14090 18952 14096 18964
rect 14051 18924 14096 18952
rect 14090 18912 14096 18924
rect 14148 18912 14154 18964
rect 36262 18952 36268 18964
rect 14200 18924 36268 18952
rect 13722 18844 13728 18896
rect 13780 18884 13786 18896
rect 14200 18884 14228 18924
rect 36262 18912 36268 18924
rect 36320 18912 36326 18964
rect 13780 18856 14228 18884
rect 14737 18887 14795 18893
rect 13780 18844 13786 18856
rect 14737 18853 14749 18887
rect 14783 18853 14795 18887
rect 20714 18884 20720 18896
rect 14737 18847 14795 18853
rect 20180 18856 20720 18884
rect 11790 18816 11796 18828
rect 11751 18788 11796 18816
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 12066 18816 12072 18828
rect 12027 18788 12072 18816
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 14752 18816 14780 18847
rect 14108 18788 14780 18816
rect 2958 18748 2964 18760
rect 2919 18720 2964 18748
rect 2958 18708 2964 18720
rect 3016 18708 3022 18760
rect 13170 18708 13176 18760
rect 13228 18708 13234 18760
rect 14108 18757 14136 18788
rect 14093 18751 14151 18757
rect 14093 18717 14105 18751
rect 14139 18717 14151 18751
rect 14274 18748 14280 18760
rect 14235 18720 14280 18748
rect 14093 18711 14151 18717
rect 14274 18708 14280 18720
rect 14332 18708 14338 18760
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18748 14795 18751
rect 14826 18748 14832 18760
rect 14783 18720 14832 18748
rect 14783 18717 14795 18720
rect 14737 18711 14795 18717
rect 14826 18708 14832 18720
rect 14884 18708 14890 18760
rect 15010 18748 15016 18760
rect 14971 18720 15016 18748
rect 15010 18708 15016 18720
rect 15068 18708 15074 18760
rect 16574 18708 16580 18760
rect 16632 18748 16638 18760
rect 20180 18757 20208 18856
rect 20714 18844 20720 18856
rect 20772 18844 20778 18896
rect 23750 18844 23756 18896
rect 23808 18884 23814 18896
rect 24765 18887 24823 18893
rect 24765 18884 24777 18887
rect 23808 18856 24777 18884
rect 23808 18844 23814 18856
rect 24765 18853 24777 18856
rect 24811 18853 24823 18887
rect 27154 18884 27160 18896
rect 27115 18856 27160 18884
rect 24765 18847 24823 18853
rect 27154 18844 27160 18856
rect 27212 18844 27218 18896
rect 28905 18887 28963 18893
rect 28905 18884 28917 18887
rect 28000 18856 28917 18884
rect 20254 18776 20260 18828
rect 20312 18816 20318 18828
rect 20312 18788 20392 18816
rect 20312 18776 20318 18788
rect 20364 18757 20392 18788
rect 24854 18776 24860 18828
rect 24912 18816 24918 18828
rect 25685 18819 25743 18825
rect 25685 18816 25697 18819
rect 24912 18788 25697 18816
rect 24912 18776 24918 18788
rect 25685 18785 25697 18788
rect 25731 18785 25743 18819
rect 25685 18779 25743 18785
rect 27798 18776 27804 18828
rect 27856 18816 27862 18828
rect 27893 18819 27951 18825
rect 27893 18816 27905 18819
rect 27856 18788 27905 18816
rect 27856 18776 27862 18788
rect 27893 18785 27905 18788
rect 27939 18785 27951 18819
rect 27893 18779 27951 18785
rect 17129 18751 17187 18757
rect 17129 18748 17141 18751
rect 16632 18720 17141 18748
rect 16632 18708 16638 18720
rect 17129 18717 17141 18720
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 20165 18751 20223 18757
rect 20165 18717 20177 18751
rect 20211 18717 20223 18751
rect 20165 18711 20223 18717
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18717 20407 18751
rect 20806 18748 20812 18760
rect 20767 18720 20812 18748
rect 20349 18711 20407 18717
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 24394 18748 24400 18760
rect 24355 18720 24400 18748
rect 24394 18708 24400 18720
rect 24452 18708 24458 18760
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18748 24639 18751
rect 24762 18748 24768 18760
rect 24627 18720 24768 18748
rect 24627 18717 24639 18720
rect 24581 18711 24639 18717
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 25406 18748 25412 18760
rect 25367 18720 25412 18748
rect 25406 18708 25412 18720
rect 25464 18708 25470 18760
rect 28000 18757 28028 18856
rect 28905 18853 28917 18856
rect 28951 18884 28963 18887
rect 29086 18884 29092 18896
rect 28951 18856 29092 18884
rect 28951 18853 28963 18856
rect 28905 18847 28963 18853
rect 29086 18844 29092 18856
rect 29144 18844 29150 18896
rect 45649 18887 45707 18893
rect 45649 18884 45661 18887
rect 45020 18856 45661 18884
rect 29914 18776 29920 18828
rect 29972 18816 29978 18828
rect 30285 18819 30343 18825
rect 30285 18816 30297 18819
rect 29972 18788 30297 18816
rect 29972 18776 29978 18788
rect 30285 18785 30297 18788
rect 30331 18785 30343 18819
rect 30285 18779 30343 18785
rect 27985 18751 28043 18757
rect 27985 18717 27997 18751
rect 28031 18717 28043 18751
rect 27985 18711 28043 18717
rect 28718 18708 28724 18760
rect 28776 18748 28782 18760
rect 28813 18751 28871 18757
rect 28813 18748 28825 18751
rect 28776 18720 28825 18748
rect 28776 18708 28782 18720
rect 28813 18717 28825 18720
rect 28859 18717 28871 18751
rect 28994 18748 29000 18760
rect 28955 18720 29000 18748
rect 28813 18711 28871 18717
rect 28994 18708 29000 18720
rect 29052 18708 29058 18760
rect 43254 18708 43260 18760
rect 43312 18748 43318 18760
rect 43717 18751 43775 18757
rect 43717 18748 43729 18751
rect 43312 18720 43729 18748
rect 43312 18708 43318 18720
rect 43717 18717 43729 18720
rect 43763 18717 43775 18751
rect 43898 18748 43904 18760
rect 43859 18720 43904 18748
rect 43717 18711 43775 18717
rect 20257 18683 20315 18689
rect 20257 18649 20269 18683
rect 20303 18680 20315 18683
rect 21085 18683 21143 18689
rect 21085 18680 21097 18683
rect 20303 18652 21097 18680
rect 20303 18649 20315 18652
rect 20257 18643 20315 18649
rect 21085 18649 21097 18652
rect 21131 18649 21143 18683
rect 22370 18680 22376 18692
rect 22310 18652 22376 18680
rect 21085 18643 21143 18649
rect 22370 18640 22376 18652
rect 22428 18640 22434 18692
rect 27062 18680 27068 18692
rect 26910 18652 27068 18680
rect 27062 18640 27068 18652
rect 27120 18640 27126 18692
rect 30006 18640 30012 18692
rect 30064 18680 30070 18692
rect 30282 18680 30288 18692
rect 30064 18652 30288 18680
rect 30064 18640 30070 18652
rect 30282 18640 30288 18652
rect 30340 18640 30346 18692
rect 30469 18683 30527 18689
rect 30469 18649 30481 18683
rect 30515 18680 30527 18683
rect 31110 18680 31116 18692
rect 30515 18652 31116 18680
rect 30515 18649 30527 18652
rect 30469 18643 30527 18649
rect 31110 18640 31116 18652
rect 31168 18640 31174 18692
rect 31938 18640 31944 18692
rect 31996 18680 32002 18692
rect 32122 18680 32128 18692
rect 31996 18652 32128 18680
rect 31996 18640 32002 18652
rect 32122 18640 32128 18652
rect 32180 18680 32186 18692
rect 42058 18680 42064 18692
rect 32180 18652 42064 18680
rect 32180 18640 32186 18652
rect 42058 18640 42064 18652
rect 42116 18640 42122 18692
rect 43732 18680 43760 18711
rect 43898 18708 43904 18720
rect 43956 18708 43962 18760
rect 44910 18708 44916 18760
rect 44968 18748 44974 18760
rect 45020 18757 45048 18856
rect 45649 18853 45661 18856
rect 45695 18853 45707 18887
rect 45649 18847 45707 18853
rect 45462 18776 45468 18828
rect 45520 18816 45526 18828
rect 46293 18819 46351 18825
rect 46293 18816 46305 18819
rect 45520 18788 46305 18816
rect 45520 18776 45526 18788
rect 46293 18785 46305 18788
rect 46339 18785 46351 18819
rect 48130 18816 48136 18828
rect 48091 18788 48136 18816
rect 46293 18779 46351 18785
rect 48130 18776 48136 18788
rect 48188 18776 48194 18828
rect 45005 18751 45063 18757
rect 45005 18748 45017 18751
rect 44968 18720 45017 18748
rect 44968 18708 44974 18720
rect 45005 18717 45017 18720
rect 45051 18717 45063 18751
rect 45005 18711 45063 18717
rect 45094 18708 45100 18760
rect 45152 18748 45158 18760
rect 45189 18751 45247 18757
rect 45189 18748 45201 18751
rect 45152 18720 45201 18748
rect 45152 18708 45158 18720
rect 45189 18717 45201 18720
rect 45235 18717 45247 18751
rect 45830 18748 45836 18760
rect 45791 18720 45836 18748
rect 45189 18711 45247 18717
rect 45830 18708 45836 18720
rect 45888 18708 45894 18760
rect 46477 18683 46535 18689
rect 43732 18652 45140 18680
rect 14921 18615 14979 18621
rect 14921 18581 14933 18615
rect 14967 18612 14979 18615
rect 15102 18612 15108 18624
rect 14967 18584 15108 18612
rect 14967 18581 14979 18584
rect 14921 18575 14979 18581
rect 15102 18572 15108 18584
rect 15160 18572 15166 18624
rect 17310 18612 17316 18624
rect 17271 18584 17316 18612
rect 17310 18572 17316 18584
rect 17368 18572 17374 18624
rect 22554 18612 22560 18624
rect 22467 18584 22560 18612
rect 22554 18572 22560 18584
rect 22612 18612 22618 18624
rect 23106 18612 23112 18624
rect 22612 18584 23112 18612
rect 22612 18572 22618 18584
rect 23106 18572 23112 18584
rect 23164 18572 23170 18624
rect 28166 18572 28172 18624
rect 28224 18612 28230 18624
rect 28353 18615 28411 18621
rect 28353 18612 28365 18615
rect 28224 18584 28365 18612
rect 28224 18572 28230 18584
rect 28353 18581 28365 18584
rect 28399 18612 28411 18615
rect 30190 18612 30196 18624
rect 28399 18584 30196 18612
rect 28399 18581 28411 18584
rect 28353 18575 28411 18581
rect 30190 18572 30196 18584
rect 30248 18572 30254 18624
rect 43806 18612 43812 18624
rect 43767 18584 43812 18612
rect 43806 18572 43812 18584
rect 43864 18572 43870 18624
rect 45112 18621 45140 18652
rect 46477 18649 46489 18683
rect 46523 18680 46535 18683
rect 47670 18680 47676 18692
rect 46523 18652 47676 18680
rect 46523 18649 46535 18652
rect 46477 18643 46535 18649
rect 47670 18640 47676 18652
rect 47728 18640 47734 18692
rect 45097 18615 45155 18621
rect 45097 18581 45109 18615
rect 45143 18581 45155 18615
rect 45097 18575 45155 18581
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 2958 18368 2964 18420
rect 3016 18408 3022 18420
rect 12986 18408 12992 18420
rect 3016 18380 12992 18408
rect 3016 18368 3022 18380
rect 12986 18368 12992 18380
rect 13044 18368 13050 18420
rect 13170 18408 13176 18420
rect 13131 18380 13176 18408
rect 13170 18368 13176 18380
rect 13228 18368 13234 18420
rect 20806 18368 20812 18420
rect 20864 18408 20870 18420
rect 20901 18411 20959 18417
rect 20901 18408 20913 18411
rect 20864 18380 20913 18408
rect 20864 18368 20870 18380
rect 20901 18377 20913 18380
rect 20947 18377 20959 18411
rect 20901 18371 20959 18377
rect 24486 18368 24492 18420
rect 24544 18408 24550 18420
rect 29730 18408 29736 18420
rect 24544 18380 29736 18408
rect 24544 18368 24550 18380
rect 29730 18368 29736 18380
rect 29788 18368 29794 18420
rect 47670 18408 47676 18420
rect 47631 18380 47676 18408
rect 47670 18368 47676 18380
rect 47728 18368 47734 18420
rect 4614 18300 4620 18352
rect 4672 18340 4678 18352
rect 42705 18343 42763 18349
rect 4672 18312 41644 18340
rect 4672 18300 4678 18312
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 13078 18272 13084 18284
rect 13039 18244 13084 18272
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 16298 18232 16304 18284
rect 16356 18272 16362 18284
rect 16945 18275 17003 18281
rect 16945 18272 16957 18275
rect 16356 18244 16957 18272
rect 16356 18232 16362 18244
rect 16945 18241 16957 18244
rect 16991 18241 17003 18275
rect 16945 18235 17003 18241
rect 20901 18275 20959 18281
rect 20901 18241 20913 18275
rect 20947 18272 20959 18275
rect 20990 18272 20996 18284
rect 20947 18244 20996 18272
rect 20947 18241 20959 18244
rect 20901 18235 20959 18241
rect 20990 18232 20996 18244
rect 21048 18232 21054 18284
rect 22186 18232 22192 18284
rect 22244 18272 22250 18284
rect 23290 18272 23296 18284
rect 22244 18244 23296 18272
rect 22244 18232 22250 18244
rect 23290 18232 23296 18244
rect 23348 18232 23354 18284
rect 24765 18275 24823 18281
rect 24765 18241 24777 18275
rect 24811 18272 24823 18275
rect 24854 18272 24860 18284
rect 24811 18244 24860 18272
rect 24811 18241 24823 18244
rect 24765 18235 24823 18241
rect 24854 18232 24860 18244
rect 24912 18232 24918 18284
rect 27522 18272 27528 18284
rect 27483 18244 27528 18272
rect 27522 18232 27528 18244
rect 27580 18232 27586 18284
rect 28166 18272 28172 18284
rect 28127 18244 28172 18272
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 30653 18275 30711 18281
rect 30653 18241 30665 18275
rect 30699 18241 30711 18275
rect 31110 18272 31116 18284
rect 31071 18244 31116 18272
rect 30653 18235 30711 18241
rect 12986 18164 12992 18216
rect 13044 18204 13050 18216
rect 13722 18204 13728 18216
rect 13044 18176 13728 18204
rect 13044 18164 13050 18176
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 17126 18204 17132 18216
rect 17087 18176 17132 18204
rect 17126 18164 17132 18176
rect 17184 18164 17190 18216
rect 18782 18204 18788 18216
rect 18743 18176 18788 18204
rect 18782 18164 18788 18176
rect 18840 18164 18846 18216
rect 23474 18164 23480 18216
rect 23532 18204 23538 18216
rect 23569 18207 23627 18213
rect 23569 18204 23581 18207
rect 23532 18176 23581 18204
rect 23532 18164 23538 18176
rect 23569 18173 23581 18176
rect 23615 18204 23627 18207
rect 24670 18204 24676 18216
rect 23615 18176 24676 18204
rect 23615 18173 23627 18176
rect 23569 18167 23627 18173
rect 24670 18164 24676 18176
rect 24728 18164 24734 18216
rect 28353 18207 28411 18213
rect 28353 18173 28365 18207
rect 28399 18173 28411 18207
rect 28353 18167 28411 18173
rect 28629 18207 28687 18213
rect 28629 18173 28641 18207
rect 28675 18173 28687 18207
rect 30668 18204 30696 18235
rect 31110 18232 31116 18244
rect 31168 18272 31174 18284
rect 40126 18272 40132 18284
rect 31168 18244 40132 18272
rect 31168 18232 31174 18244
rect 40126 18232 40132 18244
rect 40184 18232 40190 18284
rect 40770 18272 40776 18284
rect 40731 18244 40776 18272
rect 40770 18232 40776 18244
rect 40828 18232 40834 18284
rect 40972 18281 41000 18312
rect 41616 18281 41644 18312
rect 42705 18309 42717 18343
rect 42751 18309 42763 18343
rect 42705 18303 42763 18309
rect 45373 18343 45431 18349
rect 45373 18309 45385 18343
rect 45419 18340 45431 18343
rect 46198 18340 46204 18352
rect 45419 18312 46204 18340
rect 45419 18309 45431 18312
rect 45373 18303 45431 18309
rect 40957 18275 41015 18281
rect 40957 18241 40969 18275
rect 41003 18241 41015 18275
rect 40957 18235 41015 18241
rect 41417 18275 41475 18281
rect 41417 18241 41429 18275
rect 41463 18241 41475 18275
rect 41417 18235 41475 18241
rect 41601 18275 41659 18281
rect 41601 18241 41613 18275
rect 41647 18241 41659 18275
rect 41601 18235 41659 18241
rect 42429 18275 42487 18281
rect 42429 18241 42441 18275
rect 42475 18272 42487 18275
rect 42518 18272 42524 18284
rect 42475 18244 42524 18272
rect 42475 18241 42487 18244
rect 42429 18235 42487 18241
rect 31573 18207 31631 18213
rect 31573 18204 31585 18207
rect 30668 18176 31585 18204
rect 28629 18167 28687 18173
rect 31573 18173 31585 18176
rect 31619 18173 31631 18207
rect 40788 18204 40816 18232
rect 41432 18204 41460 18235
rect 42518 18232 42524 18244
rect 42576 18232 42582 18284
rect 42720 18272 42748 18303
rect 46198 18300 46204 18312
rect 46256 18300 46262 18352
rect 43533 18275 43591 18281
rect 43533 18272 43545 18275
rect 42720 18244 43545 18272
rect 43533 18241 43545 18244
rect 43579 18241 43591 18275
rect 43806 18272 43812 18284
rect 43767 18244 43812 18272
rect 43533 18235 43591 18241
rect 43806 18232 43812 18244
rect 43864 18232 43870 18284
rect 47026 18232 47032 18284
rect 47084 18272 47090 18284
rect 47394 18272 47400 18284
rect 47084 18244 47400 18272
rect 47084 18232 47090 18244
rect 47394 18232 47400 18244
rect 47452 18272 47458 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 47452 18244 47593 18272
rect 47452 18232 47458 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47581 18235 47639 18241
rect 40788 18176 41460 18204
rect 41509 18207 41567 18213
rect 31573 18167 31631 18173
rect 41509 18173 41521 18207
rect 41555 18204 41567 18207
rect 42150 18204 42156 18216
rect 41555 18176 42156 18204
rect 41555 18173 41567 18176
rect 41509 18167 41567 18173
rect 3326 18096 3332 18148
rect 3384 18136 3390 18148
rect 27617 18139 27675 18145
rect 3384 18108 26096 18136
rect 3384 18096 3390 18108
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18068 1639 18071
rect 24486 18068 24492 18080
rect 1627 18040 24492 18068
rect 1627 18037 1639 18040
rect 1581 18031 1639 18037
rect 24486 18028 24492 18040
rect 24544 18028 24550 18080
rect 24581 18071 24639 18077
rect 24581 18037 24593 18071
rect 24627 18068 24639 18071
rect 24762 18068 24768 18080
rect 24627 18040 24768 18068
rect 24627 18037 24639 18040
rect 24581 18031 24639 18037
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 26068 18068 26096 18108
rect 27617 18105 27629 18139
rect 27663 18136 27675 18139
rect 28368 18136 28396 18167
rect 27663 18108 28396 18136
rect 27663 18105 27675 18108
rect 27617 18099 27675 18105
rect 28644 18068 28672 18167
rect 42150 18164 42156 18176
rect 42208 18204 42214 18216
rect 42705 18207 42763 18213
rect 42705 18204 42717 18207
rect 42208 18176 42717 18204
rect 42208 18164 42214 18176
rect 42705 18173 42717 18176
rect 42751 18173 42763 18207
rect 42705 18167 42763 18173
rect 44545 18207 44603 18213
rect 44545 18173 44557 18207
rect 44591 18204 44603 18207
rect 45002 18204 45008 18216
rect 44591 18176 45008 18204
rect 44591 18173 44603 18176
rect 44545 18167 44603 18173
rect 45002 18164 45008 18176
rect 45060 18204 45066 18216
rect 45189 18207 45247 18213
rect 45189 18204 45201 18207
rect 45060 18176 45201 18204
rect 45060 18164 45066 18176
rect 45189 18173 45201 18176
rect 45235 18173 45247 18207
rect 46842 18204 46848 18216
rect 46803 18176 46848 18204
rect 45189 18167 45247 18173
rect 46842 18164 46848 18176
rect 46900 18164 46906 18216
rect 40034 18136 40040 18148
rect 31404 18108 40040 18136
rect 26068 18040 28672 18068
rect 30374 18028 30380 18080
rect 30432 18068 30438 18080
rect 31404 18077 31432 18108
rect 40034 18096 40040 18108
rect 40092 18096 40098 18148
rect 42058 18096 42064 18148
rect 42116 18136 42122 18148
rect 44174 18136 44180 18148
rect 42116 18108 44180 18136
rect 42116 18096 42122 18108
rect 44174 18096 44180 18108
rect 44232 18096 44238 18148
rect 30469 18071 30527 18077
rect 30469 18068 30481 18071
rect 30432 18040 30481 18068
rect 30432 18028 30438 18040
rect 30469 18037 30481 18040
rect 30515 18037 30527 18071
rect 30469 18031 30527 18037
rect 31389 18071 31447 18077
rect 31389 18037 31401 18071
rect 31435 18037 31447 18071
rect 31389 18031 31447 18037
rect 40773 18071 40831 18077
rect 40773 18037 40785 18071
rect 40819 18068 40831 18071
rect 40954 18068 40960 18080
rect 40819 18040 40960 18068
rect 40819 18037 40831 18040
rect 40773 18031 40831 18037
rect 40954 18028 40960 18040
rect 41012 18068 41018 18080
rect 42521 18071 42579 18077
rect 42521 18068 42533 18071
rect 41012 18040 42533 18068
rect 41012 18028 41018 18040
rect 42521 18037 42533 18040
rect 42567 18037 42579 18071
rect 42521 18031 42579 18037
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 17126 17824 17132 17876
rect 17184 17864 17190 17876
rect 17221 17867 17279 17873
rect 17221 17864 17233 17867
rect 17184 17836 17233 17864
rect 17184 17824 17190 17836
rect 17221 17833 17233 17836
rect 17267 17833 17279 17867
rect 17221 17827 17279 17833
rect 21729 17867 21787 17873
rect 21729 17833 21741 17867
rect 21775 17864 21787 17867
rect 23566 17864 23572 17876
rect 21775 17836 23572 17864
rect 21775 17833 21787 17836
rect 21729 17827 21787 17833
rect 23566 17824 23572 17836
rect 23624 17864 23630 17876
rect 23750 17864 23756 17876
rect 23624 17836 23756 17864
rect 23624 17824 23630 17836
rect 23750 17824 23756 17836
rect 23808 17824 23814 17876
rect 42518 17864 42524 17876
rect 28920 17836 42524 17864
rect 14826 17756 14832 17808
rect 14884 17796 14890 17808
rect 22738 17796 22744 17808
rect 14884 17768 22744 17796
rect 14884 17756 14890 17768
rect 22738 17756 22744 17768
rect 22796 17756 22802 17808
rect 24578 17756 24584 17808
rect 24636 17796 24642 17808
rect 28920 17805 28948 17836
rect 42518 17824 42524 17836
rect 42576 17864 42582 17876
rect 42702 17864 42708 17876
rect 42576 17836 42708 17864
rect 42576 17824 42582 17836
rect 42702 17824 42708 17836
rect 42760 17824 42766 17876
rect 43898 17824 43904 17876
rect 43956 17864 43962 17876
rect 45373 17867 45431 17873
rect 45373 17864 45385 17867
rect 43956 17836 45385 17864
rect 43956 17824 43962 17836
rect 45373 17833 45385 17836
rect 45419 17833 45431 17867
rect 45373 17827 45431 17833
rect 28905 17799 28963 17805
rect 24636 17768 24808 17796
rect 24636 17756 24642 17768
rect 14642 17728 14648 17740
rect 14555 17700 14648 17728
rect 14642 17688 14648 17700
rect 14700 17728 14706 17740
rect 23382 17728 23388 17740
rect 14700 17700 23388 17728
rect 14700 17688 14706 17700
rect 23382 17688 23388 17700
rect 23440 17688 23446 17740
rect 24670 17728 24676 17740
rect 24631 17700 24676 17728
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 24780 17737 24808 17768
rect 28905 17765 28917 17799
rect 28951 17765 28963 17799
rect 28905 17759 28963 17765
rect 41325 17799 41383 17805
rect 41325 17765 41337 17799
rect 41371 17796 41383 17799
rect 42150 17796 42156 17808
rect 41371 17768 42156 17796
rect 41371 17765 41383 17768
rect 41325 17759 41383 17765
rect 42150 17756 42156 17768
rect 42208 17756 42214 17808
rect 42426 17796 42432 17808
rect 42387 17768 42432 17796
rect 42426 17756 42432 17768
rect 42484 17756 42490 17808
rect 45554 17796 45560 17808
rect 43364 17768 45560 17796
rect 24765 17731 24823 17737
rect 24765 17697 24777 17731
rect 24811 17697 24823 17731
rect 28718 17728 28724 17740
rect 24765 17691 24823 17697
rect 28184 17700 28724 17728
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 1762 17660 1768 17672
rect 1719 17632 1768 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 1762 17620 1768 17632
rect 1820 17620 1826 17672
rect 2130 17660 2136 17672
rect 2091 17632 2136 17660
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 14826 17660 14832 17672
rect 14787 17632 14832 17660
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 17129 17663 17187 17669
rect 17129 17629 17141 17663
rect 17175 17660 17187 17663
rect 17310 17660 17316 17672
rect 17175 17632 17316 17660
rect 17175 17629 17187 17632
rect 17129 17623 17187 17629
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 18506 17660 18512 17672
rect 18467 17632 18512 17660
rect 18506 17620 18512 17632
rect 18564 17620 18570 17672
rect 19150 17620 19156 17672
rect 19208 17660 19214 17672
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 19208 17632 19257 17660
rect 19208 17620 19214 17632
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 20990 17620 20996 17672
rect 21048 17660 21054 17672
rect 21545 17663 21603 17669
rect 21545 17660 21557 17663
rect 21048 17632 21557 17660
rect 21048 17620 21054 17632
rect 21545 17629 21557 17632
rect 21591 17629 21603 17663
rect 21545 17623 21603 17629
rect 23474 17620 23480 17672
rect 23532 17660 23538 17672
rect 23569 17663 23627 17669
rect 23569 17660 23581 17663
rect 23532 17632 23581 17660
rect 23532 17620 23538 17632
rect 23569 17629 23581 17632
rect 23615 17629 23627 17663
rect 23569 17623 23627 17629
rect 23661 17663 23719 17669
rect 23661 17629 23673 17663
rect 23707 17660 23719 17663
rect 24394 17660 24400 17672
rect 23707 17632 24400 17660
rect 23707 17629 23719 17632
rect 23661 17623 23719 17629
rect 24394 17620 24400 17632
rect 24452 17660 24458 17672
rect 24581 17663 24639 17669
rect 24581 17660 24593 17663
rect 24452 17632 24593 17660
rect 24452 17620 24458 17632
rect 24581 17629 24593 17632
rect 24627 17629 24639 17663
rect 24581 17623 24639 17629
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 9030 17592 9036 17604
rect 3568 17564 9036 17592
rect 3568 17552 3574 17564
rect 9030 17552 9036 17564
rect 9088 17552 9094 17604
rect 18601 17595 18659 17601
rect 18601 17561 18613 17595
rect 18647 17592 18659 17595
rect 19429 17595 19487 17601
rect 19429 17592 19441 17595
rect 18647 17564 19441 17592
rect 18647 17561 18659 17564
rect 18601 17555 18659 17561
rect 19429 17561 19441 17564
rect 19475 17561 19487 17595
rect 21082 17592 21088 17604
rect 21043 17564 21088 17592
rect 19429 17555 19487 17561
rect 21082 17552 21088 17564
rect 21140 17552 21146 17604
rect 23290 17592 23296 17604
rect 23251 17564 23296 17592
rect 23290 17552 23296 17564
rect 23348 17552 23354 17604
rect 24780 17592 24808 17691
rect 24857 17663 24915 17669
rect 24857 17629 24869 17663
rect 24903 17660 24915 17663
rect 25130 17660 25136 17672
rect 24903 17632 25136 17660
rect 24903 17629 24915 17632
rect 24857 17623 24915 17629
rect 25130 17620 25136 17632
rect 25188 17620 25194 17672
rect 25409 17663 25467 17669
rect 25409 17629 25421 17663
rect 25455 17660 25467 17663
rect 26694 17660 26700 17672
rect 25455 17632 26700 17660
rect 25455 17629 25467 17632
rect 25409 17623 25467 17629
rect 26694 17620 26700 17632
rect 26752 17620 26758 17672
rect 27798 17660 27804 17672
rect 27759 17632 27804 17660
rect 27798 17620 27804 17632
rect 27856 17620 27862 17672
rect 28184 17669 28212 17700
rect 28718 17688 28724 17700
rect 28776 17688 28782 17740
rect 30190 17728 30196 17740
rect 30151 17700 30196 17728
rect 30190 17688 30196 17700
rect 30248 17688 30254 17740
rect 30374 17728 30380 17740
rect 30335 17700 30380 17728
rect 30374 17688 30380 17700
rect 30432 17688 30438 17740
rect 32033 17731 32091 17737
rect 32033 17697 32045 17731
rect 32079 17728 32091 17731
rect 32122 17728 32128 17740
rect 32079 17700 32128 17728
rect 32079 17697 32091 17700
rect 32033 17691 32091 17697
rect 32122 17688 32128 17700
rect 32180 17688 32186 17740
rect 40954 17728 40960 17740
rect 40915 17700 40960 17728
rect 40954 17688 40960 17700
rect 41012 17728 41018 17740
rect 41012 17700 42380 17728
rect 41012 17688 41018 17700
rect 28169 17663 28227 17669
rect 28169 17629 28181 17663
rect 28215 17629 28227 17663
rect 28169 17623 28227 17629
rect 28445 17663 28503 17669
rect 28445 17629 28457 17663
rect 28491 17629 28503 17663
rect 28626 17660 28632 17672
rect 28587 17632 28632 17660
rect 28445 17623 28503 17629
rect 23492 17564 24808 17592
rect 28460 17592 28488 17623
rect 28626 17620 28632 17632
rect 28684 17620 28690 17672
rect 41877 17663 41935 17669
rect 41877 17629 41889 17663
rect 41923 17629 41935 17663
rect 42150 17660 42156 17672
rect 42111 17632 42156 17660
rect 41877 17623 41935 17629
rect 28994 17592 29000 17604
rect 28460 17564 29000 17592
rect 1946 17484 1952 17536
rect 2004 17524 2010 17536
rect 2225 17527 2283 17533
rect 2225 17524 2237 17527
rect 2004 17496 2237 17524
rect 2004 17484 2010 17496
rect 2225 17493 2237 17496
rect 2271 17493 2283 17527
rect 15010 17524 15016 17536
rect 14971 17496 15016 17524
rect 2225 17487 2283 17493
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 23492 17533 23520 17564
rect 23676 17536 23704 17564
rect 28994 17552 29000 17564
rect 29052 17552 29058 17604
rect 41892 17592 41920 17623
rect 42150 17620 42156 17632
rect 42208 17620 42214 17672
rect 42352 17669 42380 17700
rect 42337 17663 42395 17669
rect 42337 17629 42349 17663
rect 42383 17629 42395 17663
rect 43254 17660 43260 17672
rect 42337 17623 42395 17629
rect 42628 17632 43260 17660
rect 42628 17592 42656 17632
rect 43254 17620 43260 17632
rect 43312 17620 43318 17672
rect 43364 17669 43392 17768
rect 45554 17756 45560 17768
rect 45612 17756 45618 17808
rect 47946 17728 47952 17740
rect 43640 17700 47952 17728
rect 43349 17663 43407 17669
rect 43349 17629 43361 17663
rect 43395 17629 43407 17663
rect 43349 17623 43407 17629
rect 43438 17620 43444 17672
rect 43496 17660 43502 17672
rect 43640 17669 43668 17700
rect 47946 17688 47952 17700
rect 48004 17688 48010 17740
rect 43625 17663 43683 17669
rect 43496 17632 43541 17660
rect 43496 17620 43502 17632
rect 43625 17629 43637 17663
rect 43671 17629 43683 17663
rect 43625 17623 43683 17629
rect 41892 17564 42656 17592
rect 42702 17552 42708 17604
rect 42760 17592 42766 17604
rect 42760 17564 42805 17592
rect 42760 17552 42766 17564
rect 43162 17552 43168 17604
rect 43220 17592 43226 17604
rect 43640 17592 43668 17623
rect 44910 17620 44916 17672
rect 44968 17660 44974 17672
rect 45005 17663 45063 17669
rect 45005 17660 45017 17663
rect 44968 17632 45017 17660
rect 44968 17620 44974 17632
rect 45005 17629 45017 17632
rect 45051 17629 45063 17663
rect 46290 17660 46296 17672
rect 46251 17632 46296 17660
rect 45005 17623 45063 17629
rect 46290 17620 46296 17632
rect 46348 17620 46354 17672
rect 43220 17564 43668 17592
rect 43220 17552 43226 17564
rect 43714 17552 43720 17604
rect 43772 17592 43778 17604
rect 43993 17595 44051 17601
rect 43993 17592 44005 17595
rect 43772 17564 44005 17592
rect 43772 17552 43778 17564
rect 43993 17561 44005 17564
rect 44039 17561 44051 17595
rect 43993 17555 44051 17561
rect 45094 17552 45100 17604
rect 45152 17592 45158 17604
rect 45189 17595 45247 17601
rect 45189 17592 45201 17595
rect 45152 17564 45201 17592
rect 45152 17552 45158 17564
rect 45189 17561 45201 17564
rect 45235 17561 45247 17595
rect 45189 17555 45247 17561
rect 46477 17595 46535 17601
rect 46477 17561 46489 17595
rect 46523 17592 46535 17595
rect 47670 17592 47676 17604
rect 46523 17564 47676 17592
rect 46523 17561 46535 17564
rect 46477 17555 46535 17561
rect 47670 17552 47676 17564
rect 47728 17552 47734 17604
rect 48130 17592 48136 17604
rect 48091 17564 48136 17592
rect 48130 17552 48136 17564
rect 48188 17552 48194 17604
rect 23477 17527 23535 17533
rect 23477 17493 23489 17527
rect 23523 17493 23535 17527
rect 23477 17487 23535 17493
rect 23658 17484 23664 17536
rect 23716 17484 23722 17536
rect 23842 17524 23848 17536
rect 23803 17496 23848 17524
rect 23842 17484 23848 17496
rect 23900 17484 23906 17536
rect 24397 17527 24455 17533
rect 24397 17493 24409 17527
rect 24443 17524 24455 17527
rect 24670 17524 24676 17536
rect 24443 17496 24676 17524
rect 24443 17493 24455 17496
rect 24397 17487 24455 17493
rect 24670 17484 24676 17496
rect 24728 17484 24734 17536
rect 25590 17524 25596 17536
rect 25551 17496 25596 17524
rect 25590 17484 25596 17496
rect 25648 17484 25654 17536
rect 41417 17527 41475 17533
rect 41417 17493 41429 17527
rect 41463 17524 41475 17527
rect 42518 17524 42524 17536
rect 41463 17496 42524 17524
rect 41463 17493 41475 17496
rect 41417 17487 41475 17493
rect 42518 17484 42524 17496
rect 42576 17484 42582 17536
rect 43438 17484 43444 17536
rect 43496 17524 43502 17536
rect 47854 17524 47860 17536
rect 43496 17496 47860 17524
rect 43496 17484 43502 17496
rect 47854 17484 47860 17496
rect 47912 17484 47918 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 2130 17280 2136 17332
rect 2188 17320 2194 17332
rect 37642 17320 37648 17332
rect 2188 17292 37648 17320
rect 2188 17280 2194 17292
rect 37642 17280 37648 17292
rect 37700 17280 37706 17332
rect 40034 17280 40040 17332
rect 40092 17320 40098 17332
rect 43438 17320 43444 17332
rect 40092 17292 43444 17320
rect 40092 17280 40098 17292
rect 43438 17280 43444 17292
rect 43496 17280 43502 17332
rect 47670 17320 47676 17332
rect 43548 17292 46888 17320
rect 47631 17292 47676 17320
rect 1946 17252 1952 17264
rect 1907 17224 1952 17252
rect 1946 17212 1952 17224
rect 2004 17212 2010 17264
rect 20990 17252 20996 17264
rect 20272 17224 20996 17252
rect 1762 17184 1768 17196
rect 1723 17156 1768 17184
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 14829 17187 14887 17193
rect 14829 17153 14841 17187
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17184 15439 17187
rect 15654 17184 15660 17196
rect 15427 17156 15660 17184
rect 15427 17153 15439 17156
rect 15381 17147 15439 17153
rect 2774 17116 2780 17128
rect 2735 17088 2780 17116
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 14844 17116 14872 17147
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 20272 17193 20300 17224
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 22186 17212 22192 17264
rect 22244 17252 22250 17264
rect 22373 17255 22431 17261
rect 22373 17252 22385 17255
rect 22244 17224 22385 17252
rect 22244 17212 22250 17224
rect 22373 17221 22385 17224
rect 22419 17221 22431 17255
rect 22738 17252 22744 17264
rect 22699 17224 22744 17252
rect 22373 17215 22431 17221
rect 22738 17212 22744 17224
rect 22796 17212 22802 17264
rect 23382 17212 23388 17264
rect 23440 17252 23446 17264
rect 23569 17255 23627 17261
rect 23569 17252 23581 17255
rect 23440 17224 23581 17252
rect 23440 17212 23446 17224
rect 23569 17221 23581 17224
rect 23615 17221 23627 17255
rect 24762 17252 24768 17264
rect 24723 17224 24768 17252
rect 23569 17215 23627 17221
rect 24762 17212 24768 17224
rect 24820 17212 24826 17264
rect 25498 17212 25504 17264
rect 25556 17212 25562 17264
rect 27798 17252 27804 17264
rect 27759 17224 27804 17252
rect 27798 17212 27804 17224
rect 27856 17212 27862 17264
rect 40126 17212 40132 17264
rect 40184 17252 40190 17264
rect 43162 17252 43168 17264
rect 40184 17224 43168 17252
rect 40184 17212 40190 17224
rect 43162 17212 43168 17224
rect 43220 17212 43226 17264
rect 27160 17196 27212 17202
rect 17957 17187 18015 17193
rect 17957 17184 17969 17187
rect 16546 17156 17969 17184
rect 14918 17116 14924 17128
rect 14831 17088 14924 17116
rect 14918 17076 14924 17088
rect 14976 17116 14982 17128
rect 16546 17116 16574 17156
rect 17957 17153 17969 17156
rect 18003 17153 18015 17187
rect 17957 17147 18015 17153
rect 20257 17187 20315 17193
rect 20257 17153 20269 17187
rect 20303 17153 20315 17187
rect 22462 17184 22468 17196
rect 22423 17156 22468 17184
rect 20257 17147 20315 17153
rect 14976 17088 16574 17116
rect 14976 17076 14982 17088
rect 17972 17048 18000 17147
rect 22462 17144 22468 17156
rect 22520 17144 22526 17196
rect 22557 17187 22615 17193
rect 22557 17153 22569 17187
rect 22603 17153 22615 17187
rect 23474 17184 23480 17196
rect 23435 17156 23480 17184
rect 22557 17147 22615 17153
rect 20990 17076 20996 17128
rect 21048 17116 21054 17128
rect 22572 17116 22600 17147
rect 23474 17144 23480 17156
rect 23532 17144 23538 17196
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17153 23719 17187
rect 23661 17147 23719 17153
rect 23676 17116 23704 17147
rect 26878 17144 26884 17196
rect 26936 17184 26942 17196
rect 27065 17187 27123 17193
rect 27065 17184 27077 17187
rect 26936 17156 27077 17184
rect 26936 17144 26942 17156
rect 27065 17153 27077 17156
rect 27111 17153 27123 17187
rect 27065 17147 27123 17153
rect 42613 17187 42671 17193
rect 42613 17153 42625 17187
rect 42659 17184 42671 17187
rect 42702 17184 42708 17196
rect 42659 17156 42708 17184
rect 42659 17153 42671 17156
rect 42613 17147 42671 17153
rect 42702 17144 42708 17156
rect 42760 17144 42766 17196
rect 43548 17184 43576 17292
rect 43714 17252 43720 17264
rect 43675 17224 43720 17252
rect 43714 17212 43720 17224
rect 43772 17212 43778 17264
rect 42812 17156 43576 17184
rect 27160 17138 27212 17144
rect 24486 17116 24492 17128
rect 21048 17088 22600 17116
rect 23216 17088 23704 17116
rect 24447 17088 24492 17116
rect 21048 17076 21054 17088
rect 20438 17048 20444 17060
rect 17972 17020 20444 17048
rect 20438 17008 20444 17020
rect 20496 17008 20502 17060
rect 21818 17008 21824 17060
rect 21876 17048 21882 17060
rect 22189 17051 22247 17057
rect 22189 17048 22201 17051
rect 21876 17020 22201 17048
rect 21876 17008 21882 17020
rect 22189 17017 22201 17020
rect 22235 17017 22247 17051
rect 22189 17011 22247 17017
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 14645 16983 14703 16989
rect 14645 16980 14657 16983
rect 14424 16952 14657 16980
rect 14424 16940 14430 16952
rect 14645 16949 14657 16952
rect 14691 16949 14703 16983
rect 14645 16943 14703 16949
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 15473 16983 15531 16989
rect 15473 16980 15485 16983
rect 15436 16952 15485 16980
rect 15436 16940 15442 16952
rect 15473 16949 15485 16952
rect 15519 16949 15531 16983
rect 15473 16943 15531 16949
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 18049 16983 18107 16989
rect 18049 16980 18061 16983
rect 18012 16952 18061 16980
rect 18012 16940 18018 16952
rect 18049 16949 18061 16952
rect 18095 16949 18107 16983
rect 22204 16980 22232 17011
rect 22462 17008 22468 17060
rect 22520 17048 22526 17060
rect 23216 17048 23244 17088
rect 24486 17076 24492 17088
rect 24544 17076 24550 17128
rect 25130 17116 25136 17128
rect 24596 17088 25136 17116
rect 22520 17020 23244 17048
rect 22520 17008 22526 17020
rect 23290 17008 23296 17060
rect 23348 17048 23354 17060
rect 24596 17048 24624 17088
rect 25130 17076 25136 17088
rect 25188 17116 25194 17128
rect 26237 17119 26295 17125
rect 26237 17116 26249 17119
rect 25188 17088 26249 17116
rect 25188 17076 25194 17088
rect 26237 17085 26249 17088
rect 26283 17085 26295 17119
rect 26237 17079 26295 17085
rect 29273 17119 29331 17125
rect 29273 17085 29285 17119
rect 29319 17085 29331 17119
rect 29454 17116 29460 17128
rect 29415 17088 29460 17116
rect 29273 17079 29331 17085
rect 23348 17020 24624 17048
rect 23348 17008 23354 17020
rect 25774 17008 25780 17060
rect 25832 17048 25838 17060
rect 29288 17048 29316 17079
rect 29454 17076 29460 17088
rect 29512 17076 29518 17128
rect 31110 17116 31116 17128
rect 31071 17088 31116 17116
rect 31110 17076 31116 17088
rect 31168 17076 31174 17128
rect 42518 17116 42524 17128
rect 42479 17088 42524 17116
rect 42518 17076 42524 17088
rect 42576 17076 42582 17128
rect 25832 17020 29316 17048
rect 25832 17008 25838 17020
rect 40678 17008 40684 17060
rect 40736 17048 40742 17060
rect 42812 17048 42840 17156
rect 46290 17144 46296 17196
rect 46348 17184 46354 17196
rect 46860 17193 46888 17292
rect 47670 17280 47676 17292
rect 47728 17280 47734 17332
rect 46385 17187 46443 17193
rect 46385 17184 46397 17187
rect 46348 17156 46397 17184
rect 46348 17144 46354 17156
rect 46385 17153 46397 17156
rect 46431 17153 46443 17187
rect 46385 17147 46443 17153
rect 46845 17187 46903 17193
rect 46845 17153 46857 17187
rect 46891 17153 46903 17187
rect 46845 17147 46903 17153
rect 47581 17187 47639 17193
rect 47581 17153 47593 17187
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 43533 17119 43591 17125
rect 43533 17116 43545 17119
rect 42996 17088 43545 17116
rect 42996 17057 43024 17088
rect 43533 17085 43545 17088
rect 43579 17116 43591 17119
rect 43898 17116 43904 17128
rect 43579 17088 43904 17116
rect 43579 17085 43591 17088
rect 43533 17079 43591 17085
rect 43898 17076 43904 17088
rect 43956 17076 43962 17128
rect 44174 17116 44180 17128
rect 44135 17088 44180 17116
rect 44174 17076 44180 17088
rect 44232 17116 44238 17128
rect 46750 17116 46756 17128
rect 44232 17088 46756 17116
rect 44232 17076 44238 17088
rect 46750 17076 46756 17088
rect 46808 17076 46814 17128
rect 47596 17060 47624 17147
rect 40736 17020 42840 17048
rect 42981 17051 43039 17057
rect 40736 17008 40742 17020
rect 42981 17017 42993 17051
rect 43027 17017 43039 17051
rect 42981 17011 43039 17017
rect 44266 17008 44272 17060
rect 44324 17048 44330 17060
rect 47578 17048 47584 17060
rect 44324 17020 47584 17048
rect 44324 17008 44330 17020
rect 47578 17008 47584 17020
rect 47636 17008 47642 17060
rect 23308 16980 23336 17008
rect 22204 16952 23336 16980
rect 18049 16943 18107 16949
rect 23474 16940 23480 16992
rect 23532 16980 23538 16992
rect 23845 16983 23903 16989
rect 23845 16980 23857 16983
rect 23532 16952 23857 16980
rect 23532 16940 23538 16952
rect 23845 16949 23857 16952
rect 23891 16949 23903 16983
rect 46934 16980 46940 16992
rect 46895 16952 46940 16980
rect 23845 16943 23903 16949
rect 46934 16940 46940 16952
rect 46992 16940 46998 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 22554 16736 22560 16788
rect 22612 16776 22618 16788
rect 23017 16779 23075 16785
rect 23017 16776 23029 16779
rect 22612 16748 23029 16776
rect 22612 16736 22618 16748
rect 23017 16745 23029 16748
rect 23063 16745 23075 16779
rect 23017 16739 23075 16745
rect 23106 16736 23112 16788
rect 23164 16776 23170 16788
rect 25774 16776 25780 16788
rect 23164 16748 25780 16776
rect 23164 16736 23170 16748
rect 25774 16736 25780 16748
rect 25832 16736 25838 16788
rect 27249 16779 27307 16785
rect 27249 16745 27261 16779
rect 27295 16776 27307 16779
rect 28626 16776 28632 16788
rect 27295 16748 28632 16776
rect 27295 16745 27307 16748
rect 27249 16739 27307 16745
rect 28626 16736 28632 16748
rect 28684 16736 28690 16788
rect 29454 16736 29460 16788
rect 29512 16776 29518 16788
rect 29641 16779 29699 16785
rect 29641 16776 29653 16779
rect 29512 16748 29653 16776
rect 29512 16736 29518 16748
rect 29641 16745 29653 16748
rect 29687 16745 29699 16779
rect 29641 16739 29699 16745
rect 21836 16680 22094 16708
rect 14366 16640 14372 16652
rect 14327 16612 14372 16640
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 15654 16600 15660 16652
rect 15712 16640 15718 16652
rect 17586 16640 17592 16652
rect 15712 16612 16896 16640
rect 17547 16612 17592 16640
rect 15712 16600 15718 16612
rect 16868 16581 16896 16612
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 18049 16643 18107 16649
rect 18049 16609 18061 16643
rect 18095 16640 18107 16643
rect 18230 16640 18236 16652
rect 18095 16612 18236 16640
rect 18095 16609 18107 16612
rect 18049 16603 18107 16609
rect 18230 16600 18236 16612
rect 18288 16600 18294 16652
rect 19978 16640 19984 16652
rect 19891 16612 19984 16640
rect 19978 16600 19984 16612
rect 20036 16640 20042 16652
rect 21836 16640 21864 16680
rect 20036 16612 21864 16640
rect 22066 16640 22094 16680
rect 22462 16668 22468 16720
rect 22520 16708 22526 16720
rect 23201 16711 23259 16717
rect 23201 16708 23213 16711
rect 22520 16680 23213 16708
rect 22520 16668 22526 16680
rect 23201 16677 23213 16680
rect 23247 16677 23259 16711
rect 24670 16708 24676 16720
rect 23201 16671 23259 16677
rect 23768 16680 24532 16708
rect 24631 16680 24676 16708
rect 23768 16640 23796 16680
rect 22066 16612 23796 16640
rect 20036 16600 20042 16612
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16574 16911 16575
rect 17681 16575 17739 16581
rect 16899 16546 16933 16574
rect 16899 16541 16911 16546
rect 16853 16535 16911 16541
rect 17681 16541 17693 16575
rect 17727 16572 17739 16575
rect 18138 16572 18144 16584
rect 17727 16544 18144 16572
rect 17727 16541 17739 16544
rect 17681 16535 17739 16541
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 19613 16575 19671 16581
rect 19613 16541 19625 16575
rect 19659 16572 19671 16575
rect 19996 16572 20024 16600
rect 21836 16581 21864 16612
rect 23842 16600 23848 16652
rect 23900 16640 23906 16652
rect 24397 16643 24455 16649
rect 24397 16640 24409 16643
rect 23900 16612 24409 16640
rect 23900 16600 23906 16612
rect 24397 16609 24409 16612
rect 24443 16609 24455 16643
rect 24504 16640 24532 16680
rect 24670 16668 24676 16680
rect 24728 16668 24734 16720
rect 25222 16640 25228 16652
rect 24504 16612 25228 16640
rect 24397 16603 24455 16609
rect 25222 16600 25228 16612
rect 25280 16640 25286 16652
rect 25590 16640 25596 16652
rect 25280 16612 25596 16640
rect 25280 16600 25286 16612
rect 25424 16581 25452 16612
rect 25590 16600 25596 16612
rect 25648 16600 25654 16652
rect 26878 16640 26884 16652
rect 26839 16612 26884 16640
rect 26878 16600 26884 16612
rect 26936 16600 26942 16652
rect 27154 16640 27160 16652
rect 27080 16612 27160 16640
rect 19659 16544 20024 16572
rect 21821 16575 21879 16581
rect 19659 16541 19671 16544
rect 19613 16535 19671 16541
rect 21821 16541 21833 16575
rect 21867 16541 21879 16575
rect 25409 16575 25467 16581
rect 21821 16535 21879 16541
rect 21928 16544 25360 16572
rect 14642 16504 14648 16516
rect 14603 16476 14648 16504
rect 14642 16464 14648 16476
rect 14700 16464 14706 16516
rect 15378 16464 15384 16516
rect 15436 16464 15442 16516
rect 16393 16507 16451 16513
rect 16393 16473 16405 16507
rect 16439 16504 16451 16507
rect 16574 16504 16580 16516
rect 16439 16476 16580 16504
rect 16439 16473 16451 16476
rect 16393 16467 16451 16473
rect 16574 16464 16580 16476
rect 16632 16464 16638 16516
rect 18782 16464 18788 16516
rect 18840 16504 18846 16516
rect 21928 16504 21956 16544
rect 18840 16476 21956 16504
rect 18840 16464 18846 16476
rect 22094 16464 22100 16516
rect 22152 16504 22158 16516
rect 22833 16507 22891 16513
rect 22833 16504 22845 16507
rect 22152 16476 22845 16504
rect 22152 16464 22158 16476
rect 22833 16473 22845 16476
rect 22879 16473 22891 16507
rect 22833 16467 22891 16473
rect 23049 16507 23107 16513
rect 23049 16473 23061 16507
rect 23095 16504 23107 16507
rect 23658 16504 23664 16516
rect 23095 16476 23664 16504
rect 23095 16473 23107 16476
rect 23049 16467 23107 16473
rect 23658 16464 23664 16476
rect 23716 16464 23722 16516
rect 25332 16504 25360 16544
rect 25409 16541 25421 16575
rect 25455 16541 25467 16575
rect 25409 16535 25467 16541
rect 25498 16532 25504 16584
rect 25556 16572 25562 16584
rect 27080 16581 27108 16612
rect 27154 16600 27160 16612
rect 27212 16600 27218 16652
rect 29270 16600 29276 16652
rect 29328 16640 29334 16652
rect 29328 16612 29592 16640
rect 29328 16600 29334 16612
rect 29564 16584 29592 16612
rect 44910 16600 44916 16652
rect 44968 16640 44974 16652
rect 46293 16643 46351 16649
rect 44968 16612 45048 16640
rect 44968 16600 44974 16612
rect 27065 16575 27123 16581
rect 25556 16544 25601 16572
rect 25556 16532 25562 16544
rect 27065 16541 27077 16575
rect 27111 16541 27123 16575
rect 29546 16572 29552 16584
rect 29459 16544 29552 16572
rect 27065 16535 27123 16541
rect 29546 16532 29552 16544
rect 29604 16532 29610 16584
rect 45020 16581 45048 16612
rect 46293 16609 46305 16643
rect 46339 16640 46351 16643
rect 47762 16640 47768 16652
rect 46339 16612 47768 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47762 16600 47768 16612
rect 47820 16600 47826 16652
rect 45005 16575 45063 16581
rect 45005 16541 45017 16575
rect 45051 16574 45063 16575
rect 45051 16546 45085 16574
rect 45051 16541 45063 16546
rect 45005 16535 45063 16541
rect 46290 16504 46296 16516
rect 25332 16476 46296 16504
rect 46290 16464 46296 16476
rect 46348 16464 46354 16516
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 46934 16504 46940 16516
rect 46523 16476 46940 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 46934 16464 46940 16476
rect 46992 16464 46998 16516
rect 48130 16504 48136 16516
rect 48091 16476 48136 16504
rect 48130 16464 48136 16476
rect 48188 16464 48194 16516
rect 16942 16436 16948 16448
rect 16903 16408 16948 16436
rect 16942 16396 16948 16408
rect 17000 16396 17006 16448
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 19705 16439 19763 16445
rect 19705 16436 19717 16439
rect 19392 16408 19717 16436
rect 19392 16396 19398 16408
rect 19705 16405 19717 16408
rect 19751 16405 19763 16439
rect 21910 16436 21916 16448
rect 21871 16408 21916 16436
rect 19705 16399 19763 16405
rect 21910 16396 21916 16408
rect 21968 16396 21974 16448
rect 24854 16436 24860 16448
rect 24815 16408 24860 16436
rect 24854 16396 24860 16408
rect 24912 16396 24918 16448
rect 45097 16439 45155 16445
rect 45097 16405 45109 16439
rect 45143 16436 45155 16439
rect 45186 16436 45192 16448
rect 45143 16408 45192 16436
rect 45143 16405 45155 16408
rect 45097 16399 45155 16405
rect 45186 16396 45192 16408
rect 45244 16396 45250 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 15102 16232 15108 16244
rect 13924 16204 15108 16232
rect 13924 16105 13952 16204
rect 15102 16192 15108 16204
rect 15160 16232 15166 16244
rect 16574 16232 16580 16244
rect 15160 16204 16580 16232
rect 15160 16192 15166 16204
rect 16574 16192 16580 16204
rect 16632 16192 16638 16244
rect 17497 16235 17555 16241
rect 17497 16201 17509 16235
rect 17543 16232 17555 16235
rect 20990 16232 20996 16244
rect 17543 16204 20996 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 24486 16192 24492 16244
rect 24544 16232 24550 16244
rect 24581 16235 24639 16241
rect 24581 16232 24593 16235
rect 24544 16204 24593 16232
rect 24544 16192 24550 16204
rect 24581 16201 24593 16204
rect 24627 16201 24639 16235
rect 24581 16195 24639 16201
rect 15010 16164 15016 16176
rect 14016 16136 15016 16164
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16065 13967 16099
rect 13909 16059 13967 16065
rect 14016 16037 14044 16136
rect 15010 16124 15016 16136
rect 15068 16164 15074 16176
rect 17129 16167 17187 16173
rect 17129 16164 17141 16167
rect 15068 16136 15700 16164
rect 15068 16124 15074 16136
rect 14918 16096 14924 16108
rect 14879 16068 14924 16096
rect 14918 16056 14924 16068
rect 14976 16056 14982 16108
rect 15672 16105 15700 16136
rect 16132 16136 17141 16164
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 14277 16031 14335 16037
rect 14277 15997 14289 16031
rect 14323 16028 14335 16031
rect 14642 16028 14648 16040
rect 14323 16000 14648 16028
rect 14323 15997 14335 16000
rect 14277 15991 14335 15997
rect 14642 15988 14648 16000
rect 14700 15988 14706 16040
rect 15948 16028 15976 16059
rect 16022 16056 16028 16108
rect 16080 16096 16086 16108
rect 16132 16105 16160 16136
rect 17129 16133 17141 16136
rect 17175 16133 17187 16167
rect 17129 16127 17187 16133
rect 17345 16167 17403 16173
rect 17345 16133 17357 16167
rect 17391 16164 17403 16167
rect 17862 16164 17868 16176
rect 17391 16136 17868 16164
rect 17391 16133 17403 16136
rect 17345 16127 17403 16133
rect 17862 16124 17868 16136
rect 17920 16124 17926 16176
rect 18230 16164 18236 16176
rect 18191 16136 18236 16164
rect 18230 16124 18236 16136
rect 18288 16124 18294 16176
rect 23842 16164 23848 16176
rect 22664 16136 23848 16164
rect 16117 16099 16175 16105
rect 16117 16096 16129 16099
rect 16080 16068 16129 16096
rect 16080 16056 16086 16068
rect 16117 16065 16129 16068
rect 16163 16065 16175 16099
rect 17954 16096 17960 16108
rect 17915 16068 17960 16096
rect 16117 16059 16175 16065
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 19334 16056 19340 16108
rect 19392 16056 19398 16108
rect 19794 16056 19800 16108
rect 19852 16096 19858 16108
rect 20438 16096 20444 16108
rect 19852 16068 20444 16096
rect 19852 16056 19858 16068
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 22094 16056 22100 16108
rect 22152 16096 22158 16108
rect 22373 16099 22431 16105
rect 22373 16096 22385 16099
rect 22152 16068 22385 16096
rect 22152 16056 22158 16068
rect 22373 16065 22385 16068
rect 22419 16065 22431 16099
rect 22554 16096 22560 16108
rect 22515 16068 22560 16096
rect 22373 16059 22431 16065
rect 22554 16056 22560 16068
rect 22612 16056 22618 16108
rect 22664 16105 22692 16136
rect 23842 16124 23848 16136
rect 23900 16124 23906 16176
rect 22649 16099 22707 16105
rect 22649 16065 22661 16099
rect 22695 16065 22707 16099
rect 22649 16059 22707 16065
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16065 23167 16099
rect 23109 16059 23167 16065
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16096 23351 16099
rect 23474 16096 23480 16108
rect 23339 16068 23480 16096
rect 23339 16065 23351 16068
rect 23293 16059 23351 16065
rect 17770 16028 17776 16040
rect 15948 16000 17776 16028
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 23124 16028 23152 16059
rect 23474 16056 23480 16068
rect 23532 16056 23538 16108
rect 23750 16096 23756 16108
rect 23711 16068 23756 16096
rect 23750 16056 23756 16068
rect 23808 16096 23814 16108
rect 24397 16099 24455 16105
rect 24397 16096 24409 16099
rect 23808 16068 24409 16096
rect 23808 16056 23814 16068
rect 24397 16065 24409 16068
rect 24443 16065 24455 16099
rect 43898 16096 43904 16108
rect 43859 16068 43904 16096
rect 24397 16059 24455 16065
rect 43898 16056 43904 16068
rect 43956 16056 43962 16108
rect 47762 16096 47768 16108
rect 47723 16068 47768 16096
rect 47762 16056 47768 16068
rect 47820 16056 47826 16108
rect 44082 16028 44088 16040
rect 22388 16000 23152 16028
rect 44043 16000 44088 16028
rect 22388 15969 22416 16000
rect 44082 15988 44088 16000
rect 44140 15988 44146 16040
rect 45462 16028 45468 16040
rect 45423 16000 45468 16028
rect 45462 15988 45468 16000
rect 45520 15988 45526 16040
rect 22373 15963 22431 15969
rect 22373 15929 22385 15963
rect 22419 15929 22431 15963
rect 22373 15923 22431 15929
rect 14918 15892 14924 15904
rect 14879 15864 14924 15892
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 15194 15852 15200 15904
rect 15252 15892 15258 15904
rect 15473 15895 15531 15901
rect 15473 15892 15485 15895
rect 15252 15864 15485 15892
rect 15252 15852 15258 15864
rect 15473 15861 15485 15864
rect 15519 15861 15531 15895
rect 15473 15855 15531 15861
rect 17313 15895 17371 15901
rect 17313 15861 17325 15895
rect 17359 15892 17371 15895
rect 17954 15892 17960 15904
rect 17359 15864 17960 15892
rect 17359 15861 17371 15864
rect 17313 15855 17371 15861
rect 17954 15852 17960 15864
rect 18012 15852 18018 15904
rect 18598 15852 18604 15904
rect 18656 15892 18662 15904
rect 19705 15895 19763 15901
rect 19705 15892 19717 15895
rect 18656 15864 19717 15892
rect 18656 15852 18662 15864
rect 19705 15861 19717 15864
rect 19751 15861 19763 15895
rect 19705 15855 19763 15861
rect 20625 15895 20683 15901
rect 20625 15861 20637 15895
rect 20671 15892 20683 15895
rect 20898 15892 20904 15904
rect 20671 15864 20904 15892
rect 20671 15861 20683 15864
rect 20625 15855 20683 15861
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 23106 15892 23112 15904
rect 23067 15864 23112 15892
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 23845 15895 23903 15901
rect 23845 15861 23857 15895
rect 23891 15892 23903 15895
rect 24394 15892 24400 15904
rect 23891 15864 24400 15892
rect 23891 15861 23903 15864
rect 23845 15855 23903 15861
rect 24394 15852 24400 15864
rect 24452 15852 24458 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 17589 15691 17647 15697
rect 17589 15657 17601 15691
rect 17635 15657 17647 15691
rect 17770 15688 17776 15700
rect 17731 15660 17776 15688
rect 17589 15651 17647 15657
rect 17604 15620 17632 15651
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 23474 15688 23480 15700
rect 18708 15660 23480 15688
rect 18138 15620 18144 15632
rect 17604 15592 18144 15620
rect 18138 15580 18144 15592
rect 18196 15620 18202 15632
rect 18196 15592 18644 15620
rect 18196 15580 18202 15592
rect 14918 15552 14924 15564
rect 14879 15524 14924 15552
rect 14918 15512 14924 15524
rect 14976 15512 14982 15564
rect 15194 15552 15200 15564
rect 15155 15524 15200 15552
rect 15194 15512 15200 15524
rect 15252 15512 15258 15564
rect 18616 15496 18644 15592
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 16942 15484 16948 15496
rect 16330 15456 16948 15484
rect 2041 15447 2099 15453
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 18417 15487 18475 15493
rect 18417 15453 18429 15487
rect 18463 15453 18475 15487
rect 18598 15484 18604 15496
rect 18559 15456 18604 15484
rect 18417 15447 18475 15453
rect 17405 15419 17463 15425
rect 17405 15385 17417 15419
rect 17451 15416 17463 15419
rect 17954 15416 17960 15428
rect 17451 15388 17960 15416
rect 17451 15385 17463 15388
rect 17405 15379 17463 15385
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 18432 15416 18460 15447
rect 18598 15444 18604 15456
rect 18656 15444 18662 15496
rect 18708 15416 18736 15660
rect 23474 15648 23480 15660
rect 23532 15648 23538 15700
rect 44082 15688 44088 15700
rect 44043 15660 44088 15688
rect 44082 15648 44088 15660
rect 44140 15648 44146 15700
rect 47302 15620 47308 15632
rect 44008 15592 47308 15620
rect 20898 15552 20904 15564
rect 20859 15524 20904 15552
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 21177 15555 21235 15561
rect 21177 15521 21189 15555
rect 21223 15552 21235 15555
rect 23106 15552 23112 15564
rect 21223 15524 23112 15552
rect 21223 15521 21235 15524
rect 21177 15515 21235 15521
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 23569 15555 23627 15561
rect 23569 15521 23581 15555
rect 23615 15552 23627 15555
rect 23750 15552 23756 15564
rect 23615 15524 23756 15552
rect 23615 15521 23627 15524
rect 23569 15515 23627 15521
rect 23750 15512 23756 15524
rect 23808 15512 23814 15564
rect 23845 15555 23903 15561
rect 23845 15521 23857 15555
rect 23891 15552 23903 15555
rect 24673 15555 24731 15561
rect 24673 15552 24685 15555
rect 23891 15524 24685 15552
rect 23891 15521 23903 15524
rect 23845 15515 23903 15521
rect 24673 15521 24685 15524
rect 24719 15521 24731 15555
rect 24673 15515 24731 15521
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15484 19487 15487
rect 19794 15484 19800 15496
rect 19475 15456 19800 15484
rect 19475 15453 19487 15456
rect 19429 15447 19487 15453
rect 19794 15444 19800 15456
rect 19852 15444 19858 15496
rect 19978 15484 19984 15496
rect 19939 15456 19984 15484
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 22554 15444 22560 15496
rect 22612 15484 22618 15496
rect 23477 15487 23535 15493
rect 23477 15484 23489 15487
rect 22612 15456 23489 15484
rect 22612 15444 22618 15456
rect 23477 15453 23489 15456
rect 23523 15453 23535 15487
rect 24394 15484 24400 15496
rect 24355 15456 24400 15484
rect 23477 15447 23535 15453
rect 18064 15388 18736 15416
rect 15930 15308 15936 15360
rect 15988 15348 15994 15360
rect 16669 15351 16727 15357
rect 16669 15348 16681 15351
rect 15988 15320 16681 15348
rect 15988 15308 15994 15320
rect 16669 15317 16681 15320
rect 16715 15317 16727 15351
rect 17586 15348 17592 15360
rect 17644 15357 17650 15360
rect 17644 15351 17673 15357
rect 17525 15320 17592 15348
rect 16669 15311 16727 15317
rect 17586 15308 17592 15320
rect 17661 15348 17673 15351
rect 18064 15348 18092 15388
rect 21910 15376 21916 15428
rect 21968 15376 21974 15428
rect 17661 15320 18092 15348
rect 17661 15317 17673 15320
rect 17644 15311 17673 15317
rect 17644 15308 17650 15311
rect 18138 15308 18144 15360
rect 18196 15348 18202 15360
rect 18509 15351 18567 15357
rect 18509 15348 18521 15351
rect 18196 15320 18521 15348
rect 18196 15308 18202 15320
rect 18509 15317 18521 15320
rect 18555 15317 18567 15351
rect 19426 15348 19432 15360
rect 19387 15320 19432 15348
rect 18509 15311 18567 15317
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 20073 15351 20131 15357
rect 20073 15317 20085 15351
rect 20119 15348 20131 15351
rect 20162 15348 20168 15360
rect 20119 15320 20168 15348
rect 20119 15317 20131 15320
rect 20073 15311 20131 15317
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 22094 15308 22100 15360
rect 22152 15348 22158 15360
rect 22649 15351 22707 15357
rect 22649 15348 22661 15351
rect 22152 15320 22661 15348
rect 22152 15308 22158 15320
rect 22649 15317 22661 15320
rect 22695 15317 22707 15351
rect 23492 15348 23520 15447
rect 24394 15444 24400 15456
rect 24452 15444 24458 15496
rect 40862 15444 40868 15496
rect 40920 15484 40926 15496
rect 44008 15493 44036 15592
rect 47302 15580 47308 15592
rect 47360 15580 47366 15632
rect 45002 15552 45008 15564
rect 44963 15524 45008 15552
rect 45002 15512 45008 15524
rect 45060 15512 45066 15564
rect 45186 15552 45192 15564
rect 45147 15524 45192 15552
rect 45186 15512 45192 15524
rect 45244 15512 45250 15564
rect 46658 15552 46664 15564
rect 46619 15524 46664 15552
rect 46658 15512 46664 15524
rect 46716 15512 46722 15564
rect 43993 15487 44051 15493
rect 43993 15484 44005 15487
rect 40920 15456 44005 15484
rect 40920 15444 40926 15456
rect 43993 15453 44005 15456
rect 44039 15453 44051 15487
rect 43993 15447 44051 15453
rect 25314 15376 25320 15428
rect 25372 15376 25378 15428
rect 26145 15351 26203 15357
rect 26145 15348 26157 15351
rect 23492 15320 26157 15348
rect 22649 15311 22707 15317
rect 26145 15317 26157 15320
rect 26191 15317 26203 15351
rect 26145 15311 26203 15317
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 18417 15147 18475 15153
rect 18417 15113 18429 15147
rect 18463 15113 18475 15147
rect 25314 15144 25320 15156
rect 25275 15116 25320 15144
rect 18417 15107 18475 15113
rect 18432 15076 18460 15107
rect 25314 15104 25320 15116
rect 25372 15104 25378 15156
rect 19153 15079 19211 15085
rect 19153 15076 19165 15079
rect 18432 15048 19165 15076
rect 19153 15045 19165 15048
rect 19199 15045 19211 15079
rect 19153 15039 19211 15045
rect 20162 15036 20168 15088
rect 20220 15036 20226 15088
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 15008 16727 15011
rect 16758 15008 16764 15020
rect 16715 14980 16764 15008
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 16758 14968 16764 14980
rect 16816 15008 16822 15020
rect 17310 15008 17316 15020
rect 16816 14980 17316 15008
rect 16816 14968 16822 14980
rect 17310 14968 17316 14980
rect 17368 14968 17374 15020
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18049 15011 18107 15017
rect 18049 15008 18061 15011
rect 18012 14980 18061 15008
rect 18012 14968 18018 14980
rect 18049 14977 18061 14980
rect 18095 14977 18107 15011
rect 25222 15008 25228 15020
rect 25183 14980 25228 15008
rect 18049 14971 18107 14977
rect 25222 14968 25228 14980
rect 25280 14968 25286 15020
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 18138 14940 18144 14952
rect 18099 14912 18144 14940
rect 18138 14900 18144 14912
rect 18196 14900 18202 14952
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14940 18935 14943
rect 19518 14940 19524 14952
rect 18923 14912 19524 14940
rect 18923 14909 18935 14912
rect 18877 14903 18935 14909
rect 19518 14900 19524 14912
rect 19576 14900 19582 14952
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 22278 14940 22284 14952
rect 22152 14912 22197 14940
rect 22239 14912 22284 14940
rect 22152 14900 22158 14912
rect 22278 14900 22284 14912
rect 22336 14900 22342 14952
rect 23934 14940 23940 14952
rect 23895 14912 23940 14940
rect 23934 14900 23940 14912
rect 23992 14900 23998 14952
rect 16114 14764 16120 14816
rect 16172 14804 16178 14816
rect 16761 14807 16819 14813
rect 16761 14804 16773 14807
rect 16172 14776 16773 14804
rect 16172 14764 16178 14776
rect 16761 14773 16773 14776
rect 16807 14773 16819 14807
rect 16761 14767 16819 14773
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 20625 14807 20683 14813
rect 20625 14804 20637 14807
rect 18012 14776 20637 14804
rect 18012 14764 18018 14776
rect 20625 14773 20637 14776
rect 20671 14773 20683 14807
rect 20625 14767 20683 14773
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 27522 14600 27528 14612
rect 6886 14572 27528 14600
rect 2130 14396 2136 14408
rect 2091 14368 2136 14396
rect 2130 14356 2136 14368
rect 2188 14396 2194 14408
rect 6886 14396 6914 14572
rect 27522 14560 27528 14572
rect 27580 14560 27586 14612
rect 20809 14535 20867 14541
rect 2188 14368 6914 14396
rect 11624 14504 16436 14532
rect 2188 14356 2194 14368
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 11624 14260 11652 14504
rect 15930 14464 15936 14476
rect 15891 14436 15936 14464
rect 15930 14424 15936 14436
rect 15988 14424 15994 14476
rect 16114 14464 16120 14476
rect 16075 14436 16120 14464
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 16408 14473 16436 14504
rect 20809 14501 20821 14535
rect 20855 14532 20867 14535
rect 22278 14532 22284 14544
rect 20855 14504 22284 14532
rect 20855 14501 20867 14504
rect 20809 14495 20867 14501
rect 22278 14492 22284 14504
rect 22336 14492 22342 14544
rect 31202 14532 31208 14544
rect 22480 14504 31208 14532
rect 22480 14476 22508 14504
rect 31202 14492 31208 14504
rect 31260 14492 31266 14544
rect 16393 14467 16451 14473
rect 16393 14433 16405 14467
rect 16439 14433 16451 14467
rect 22462 14464 22468 14476
rect 16393 14427 16451 14433
rect 21376 14436 22468 14464
rect 21376 14405 21404 14436
rect 22462 14424 22468 14436
rect 22520 14424 22526 14476
rect 23566 14464 23572 14476
rect 23527 14436 23572 14464
rect 23566 14424 23572 14436
rect 23624 14424 23630 14476
rect 20717 14399 20775 14405
rect 20717 14365 20729 14399
rect 20763 14396 20775 14399
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 20763 14368 21373 14396
rect 20763 14365 20775 14368
rect 20717 14359 20775 14365
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 22020 14328 22048 14359
rect 22020 14300 22140 14328
rect 3384 14232 11652 14260
rect 21453 14263 21511 14269
rect 3384 14220 3390 14232
rect 21453 14229 21465 14263
rect 21499 14260 21511 14263
rect 22002 14260 22008 14272
rect 21499 14232 22008 14260
rect 21499 14229 21511 14232
rect 21453 14223 21511 14229
rect 22002 14220 22008 14232
rect 22060 14220 22066 14272
rect 22112 14260 22140 14300
rect 22186 14288 22192 14340
rect 22244 14328 22250 14340
rect 22244 14300 22289 14328
rect 22244 14288 22250 14300
rect 22554 14260 22560 14272
rect 22112 14232 22560 14260
rect 22554 14220 22560 14232
rect 22612 14220 22618 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 18233 13991 18291 13997
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 18969 13991 19027 13997
rect 18969 13988 18981 13991
rect 18279 13960 18981 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 18969 13957 18981 13960
rect 19015 13957 19027 13991
rect 22002 13988 22008 14000
rect 21963 13960 22008 13988
rect 18969 13951 19027 13957
rect 22002 13948 22008 13960
rect 22060 13948 22066 14000
rect 16758 13920 16764 13932
rect 16719 13892 16764 13920
rect 16758 13880 16764 13892
rect 16816 13920 16822 13932
rect 17405 13923 17463 13929
rect 17405 13920 17417 13923
rect 16816 13892 17417 13920
rect 16816 13880 16822 13892
rect 17405 13889 17417 13892
rect 17451 13920 17463 13923
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 17451 13892 18153 13920
rect 17451 13889 17463 13892
rect 17405 13883 17463 13889
rect 18141 13889 18153 13892
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 18598 13880 18604 13932
rect 18656 13920 18662 13932
rect 18785 13923 18843 13929
rect 18785 13920 18797 13923
rect 18656 13892 18797 13920
rect 18656 13880 18662 13892
rect 18785 13889 18797 13892
rect 18831 13889 18843 13923
rect 21818 13920 21824 13932
rect 21779 13892 21824 13920
rect 18785 13883 18843 13889
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 44542 13880 44548 13932
rect 44600 13920 44606 13932
rect 46753 13923 46811 13929
rect 46753 13920 46765 13923
rect 44600 13892 46765 13920
rect 44600 13880 44606 13892
rect 46753 13889 46765 13892
rect 46799 13889 46811 13923
rect 46753 13883 46811 13889
rect 20622 13852 20628 13864
rect 20583 13824 20628 13852
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 22830 13852 22836 13864
rect 22791 13824 22836 13852
rect 22830 13812 22836 13824
rect 22888 13812 22894 13864
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 14550 13784 14556 13796
rect 3476 13756 14556 13784
rect 3476 13744 3482 13756
rect 14550 13744 14556 13756
rect 14608 13744 14614 13796
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 16853 13719 16911 13725
rect 16853 13716 16865 13719
rect 16816 13688 16865 13716
rect 16816 13676 16822 13688
rect 16853 13685 16865 13688
rect 16899 13685 16911 13719
rect 16853 13679 16911 13685
rect 16942 13676 16948 13728
rect 17000 13716 17006 13728
rect 17497 13719 17555 13725
rect 17497 13716 17509 13719
rect 17000 13688 17509 13716
rect 17000 13676 17006 13688
rect 17497 13685 17509 13688
rect 17543 13685 17555 13719
rect 17497 13679 17555 13685
rect 46474 13676 46480 13728
rect 46532 13716 46538 13728
rect 46845 13719 46903 13725
rect 46845 13716 46857 13719
rect 46532 13688 46857 13716
rect 46532 13676 46538 13688
rect 46845 13685 46857 13688
rect 46891 13685 46903 13719
rect 46845 13679 46903 13685
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 22186 13472 22192 13524
rect 22244 13512 22250 13524
rect 22465 13515 22523 13521
rect 22465 13512 22477 13515
rect 22244 13484 22477 13512
rect 22244 13472 22250 13484
rect 22465 13481 22477 13484
rect 22511 13481 22523 13515
rect 22465 13475 22523 13481
rect 14826 13404 14832 13456
rect 14884 13444 14890 13456
rect 14884 13416 17080 13444
rect 14884 13404 14890 13416
rect 16758 13376 16764 13388
rect 16719 13348 16764 13376
rect 16758 13336 16764 13348
rect 16816 13336 16822 13388
rect 17052 13385 17080 13416
rect 17037 13379 17095 13385
rect 17037 13345 17049 13379
rect 17083 13345 17095 13379
rect 46474 13376 46480 13388
rect 46435 13348 46480 13376
rect 17037 13339 17095 13345
rect 46474 13336 46480 13348
rect 46532 13336 46538 13388
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 22373 13311 22431 13317
rect 22373 13277 22385 13311
rect 22419 13308 22431 13311
rect 22462 13308 22468 13320
rect 22419 13280 22468 13308
rect 22419 13277 22431 13280
rect 22373 13271 22431 13277
rect 16592 13240 16620 13271
rect 22462 13268 22468 13280
rect 22520 13268 22526 13320
rect 46290 13308 46296 13320
rect 46251 13280 46296 13308
rect 46290 13268 46296 13280
rect 46348 13268 46354 13320
rect 17954 13240 17960 13252
rect 16592 13212 17960 13240
rect 17954 13200 17960 13212
rect 18012 13200 18018 13252
rect 48130 13240 48136 13252
rect 48091 13212 48136 13240
rect 48130 13200 48136 13212
rect 48188 13200 48194 13252
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 16942 12900 16948 12912
rect 16903 12872 16948 12900
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 16761 12835 16819 12841
rect 16761 12832 16773 12835
rect 16632 12804 16773 12832
rect 16632 12792 16638 12804
rect 16761 12801 16773 12804
rect 16807 12801 16819 12835
rect 16761 12795 16819 12801
rect 46290 12792 46296 12844
rect 46348 12832 46354 12844
rect 47765 12835 47823 12841
rect 47765 12832 47777 12835
rect 46348 12804 47777 12832
rect 46348 12792 46354 12804
rect 47765 12801 47777 12804
rect 47811 12801 47823 12835
rect 47765 12795 47823 12801
rect 18598 12764 18604 12776
rect 18559 12736 18604 12764
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 26418 12628 26424 12640
rect 1627 12600 26424 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 26418 12588 26424 12600
rect 26476 12588 26482 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 46290 11500 46296 11552
rect 46348 11540 46354 11552
rect 47765 11543 47823 11549
rect 47765 11540 47777 11543
rect 46348 11512 47777 11540
rect 46348 11500 46354 11512
rect 47765 11509 47777 11512
rect 47811 11509 47823 11543
rect 47765 11503 47823 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 46290 11200 46296 11212
rect 46251 11172 46296 11200
rect 46290 11160 46296 11172
rect 46348 11160 46354 11212
rect 46474 11064 46480 11076
rect 46435 11036 46480 11064
rect 46474 11024 46480 11036
rect 46532 11024 46538 11076
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 10778 10996 10784 11008
rect 3200 10968 10784 10996
rect 3200 10956 3206 10968
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 46474 10752 46480 10804
rect 46532 10792 46538 10804
rect 46845 10795 46903 10801
rect 46845 10792 46857 10795
rect 46532 10764 46857 10792
rect 46532 10752 46538 10764
rect 46845 10761 46857 10764
rect 46891 10761 46903 10795
rect 46845 10755 46903 10761
rect 29546 10616 29552 10668
rect 29604 10656 29610 10668
rect 36630 10656 36636 10668
rect 29604 10628 36636 10656
rect 29604 10616 29610 10628
rect 36630 10616 36636 10628
rect 36688 10656 36694 10668
rect 46753 10659 46811 10665
rect 46753 10656 46765 10659
rect 36688 10628 46765 10656
rect 36688 10616 36694 10628
rect 46753 10625 46765 10628
rect 46799 10625 46811 10659
rect 46753 10619 46811 10625
rect 47394 10616 47400 10668
rect 47452 10656 47458 10668
rect 47581 10659 47639 10665
rect 47581 10656 47593 10659
rect 47452 10628 47593 10656
rect 47452 10616 47458 10628
rect 47581 10625 47593 10628
rect 47627 10625 47639 10659
rect 47581 10619 47639 10625
rect 46290 10452 46296 10464
rect 46251 10424 46296 10452
rect 46290 10412 46296 10424
rect 46348 10412 46354 10464
rect 46474 10412 46480 10464
rect 46532 10452 46538 10464
rect 47673 10455 47731 10461
rect 47673 10452 47685 10455
rect 46532 10424 47685 10452
rect 46532 10412 46538 10424
rect 47673 10421 47685 10424
rect 47719 10421 47731 10455
rect 47673 10415 47731 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 46474 10112 46480 10124
rect 46435 10084 46480 10112
rect 46474 10072 46480 10084
rect 46532 10072 46538 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 47854 9568 47860 9580
rect 47815 9540 47860 9568
rect 47854 9528 47860 9540
rect 47912 9528 47918 9580
rect 46106 9392 46112 9444
rect 46164 9432 46170 9444
rect 48041 9435 48099 9441
rect 48041 9432 48053 9435
rect 46164 9404 48053 9432
rect 46164 9392 46170 9404
rect 48041 9401 48053 9404
rect 48087 9401 48099 9435
rect 48041 9395 48099 9401
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 47762 8888 47768 8900
rect 47723 8860 47768 8888
rect 47762 8848 47768 8860
rect 47820 8848 47826 8900
rect 29822 8780 29828 8832
rect 29880 8820 29886 8832
rect 47857 8823 47915 8829
rect 47857 8820 47869 8823
rect 29880 8792 47869 8820
rect 29880 8780 29886 8792
rect 47857 8789 47869 8792
rect 47903 8789 47915 8823
rect 47857 8783 47915 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 44913 8483 44971 8489
rect 44913 8449 44925 8483
rect 44959 8480 44971 8483
rect 45278 8480 45284 8492
rect 44959 8452 45284 8480
rect 44959 8449 44971 8452
rect 44913 8443 44971 8449
rect 45278 8440 45284 8452
rect 45336 8440 45342 8492
rect 46017 8483 46075 8489
rect 46017 8480 46029 8483
rect 45526 8452 46029 8480
rect 1854 8372 1860 8424
rect 1912 8412 1918 8424
rect 44545 8415 44603 8421
rect 44545 8412 44557 8415
rect 1912 8384 44557 8412
rect 1912 8372 1918 8384
rect 44545 8381 44557 8384
rect 44591 8381 44603 8415
rect 44545 8375 44603 8381
rect 45373 8415 45431 8421
rect 45373 8381 45385 8415
rect 45419 8412 45431 8415
rect 45526 8412 45554 8452
rect 46017 8449 46029 8452
rect 46063 8449 46075 8483
rect 46017 8443 46075 8449
rect 45419 8384 45554 8412
rect 45419 8381 45431 8384
rect 45373 8375 45431 8381
rect 18598 8236 18604 8288
rect 18656 8276 18662 8288
rect 36170 8276 36176 8288
rect 18656 8248 36176 8276
rect 18656 8236 18662 8248
rect 36170 8236 36176 8248
rect 36228 8236 36234 8288
rect 44560 8276 44588 8375
rect 45005 8279 45063 8285
rect 45005 8276 45017 8279
rect 44560 8248 45017 8276
rect 45005 8245 45017 8248
rect 45051 8245 45063 8279
rect 45005 8239 45063 8245
rect 45738 8236 45744 8288
rect 45796 8276 45802 8288
rect 45833 8279 45891 8285
rect 45833 8276 45845 8279
rect 45796 8248 45845 8276
rect 45796 8236 45802 8248
rect 45833 8245 45845 8248
rect 45879 8245 45891 8279
rect 45833 8239 45891 8245
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 36170 8032 36176 8084
rect 36228 8072 36234 8084
rect 46842 8072 46848 8084
rect 36228 8044 46848 8072
rect 36228 8032 36234 8044
rect 46842 8032 46848 8044
rect 46900 8032 46906 8084
rect 45094 7964 45100 8016
rect 45152 8004 45158 8016
rect 45152 7976 45600 8004
rect 45152 7964 45158 7976
rect 45572 7945 45600 7976
rect 45557 7939 45615 7945
rect 45557 7905 45569 7939
rect 45603 7905 45615 7939
rect 45557 7899 45615 7905
rect 47486 7896 47492 7948
rect 47544 7936 47550 7948
rect 47581 7939 47639 7945
rect 47581 7936 47593 7939
rect 47544 7908 47593 7936
rect 47544 7896 47550 7908
rect 47581 7905 47593 7908
rect 47627 7905 47639 7939
rect 47581 7899 47639 7905
rect 47302 7868 47308 7880
rect 47263 7840 47308 7868
rect 47302 7828 47308 7840
rect 47360 7828 47366 7880
rect 45278 7800 45284 7812
rect 45239 7772 45284 7800
rect 45278 7760 45284 7772
rect 45336 7760 45342 7812
rect 45370 7760 45376 7812
rect 45428 7800 45434 7812
rect 45428 7772 45473 7800
rect 45428 7760 45434 7772
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 45094 7488 45100 7540
rect 45152 7528 45158 7540
rect 45152 7500 46704 7528
rect 45152 7488 45158 7500
rect 45738 7460 45744 7472
rect 45699 7432 45744 7460
rect 45738 7420 45744 7432
rect 45796 7420 45802 7472
rect 46676 7469 46704 7500
rect 46661 7463 46719 7469
rect 46661 7429 46673 7463
rect 46707 7429 46719 7463
rect 46661 7423 46719 7429
rect 48133 7395 48191 7401
rect 48133 7361 48145 7395
rect 48179 7392 48191 7395
rect 48222 7392 48228 7404
rect 48179 7364 48228 7392
rect 48179 7361 48191 7364
rect 48133 7355 48191 7361
rect 48222 7352 48228 7364
rect 48280 7352 48286 7404
rect 45649 7327 45707 7333
rect 45649 7293 45661 7327
rect 45695 7293 45707 7327
rect 45649 7287 45707 7293
rect 45664 7256 45692 7287
rect 47949 7259 48007 7265
rect 47949 7256 47961 7259
rect 45664 7228 47961 7256
rect 47949 7225 47961 7228
rect 47995 7225 48007 7259
rect 47949 7219 48007 7225
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 23934 6848 23940 6860
rect 3476 6820 23940 6848
rect 3476 6808 3482 6820
rect 23934 6808 23940 6820
rect 23992 6808 23998 6860
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 42334 6400 42340 6452
rect 42392 6440 42398 6452
rect 48041 6443 48099 6449
rect 48041 6440 48053 6443
rect 42392 6412 48053 6440
rect 42392 6400 42398 6412
rect 48041 6409 48053 6412
rect 48087 6409 48099 6443
rect 48041 6403 48099 6409
rect 47946 6304 47952 6316
rect 47907 6276 47952 6304
rect 47946 6264 47952 6276
rect 48004 6264 48010 6316
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 40126 5692 40132 5704
rect 40087 5664 40132 5692
rect 40126 5652 40132 5664
rect 40184 5652 40190 5704
rect 40218 5556 40224 5568
rect 40179 5528 40224 5556
rect 40218 5516 40224 5528
rect 40276 5516 40282 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 39669 5355 39727 5361
rect 26206 5324 37596 5352
rect 3970 5244 3976 5296
rect 4028 5284 4034 5296
rect 26206 5284 26234 5324
rect 37458 5284 37464 5296
rect 4028 5256 26234 5284
rect 37419 5256 37464 5284
rect 4028 5244 4034 5256
rect 37458 5244 37464 5256
rect 37516 5244 37522 5296
rect 37568 5284 37596 5324
rect 39669 5321 39681 5355
rect 39715 5352 39727 5355
rect 40126 5352 40132 5364
rect 39715 5324 40132 5352
rect 39715 5321 39727 5324
rect 39669 5315 39727 5321
rect 40126 5312 40132 5324
rect 40184 5312 40190 5364
rect 40310 5312 40316 5364
rect 40368 5352 40374 5364
rect 40586 5352 40592 5364
rect 40368 5324 40592 5352
rect 40368 5312 40374 5324
rect 40586 5312 40592 5324
rect 40644 5312 40650 5364
rect 43809 5355 43867 5361
rect 43809 5352 43821 5355
rect 42352 5324 43821 5352
rect 37568 5256 41414 5284
rect 18322 5216 18328 5228
rect 18283 5188 18328 5216
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 21821 5219 21879 5225
rect 21821 5185 21833 5219
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 22465 5219 22523 5225
rect 22465 5185 22477 5219
rect 22511 5216 22523 5219
rect 23842 5216 23848 5228
rect 22511 5188 23848 5216
rect 22511 5185 22523 5188
rect 22465 5179 22523 5185
rect 21836 5148 21864 5179
rect 23842 5176 23848 5188
rect 23900 5176 23906 5228
rect 38657 5219 38715 5225
rect 38657 5216 38669 5219
rect 38212 5188 38669 5216
rect 23198 5148 23204 5160
rect 21836 5120 23204 5148
rect 23198 5108 23204 5120
rect 23256 5108 23262 5160
rect 37366 5148 37372 5160
rect 37327 5120 37372 5148
rect 37366 5108 37372 5120
rect 37424 5148 37430 5160
rect 38212 5148 38240 5188
rect 38657 5185 38669 5188
rect 38703 5185 38715 5219
rect 38657 5179 38715 5185
rect 39206 5176 39212 5228
rect 39264 5216 39270 5228
rect 39577 5219 39635 5225
rect 39577 5216 39589 5219
rect 39264 5188 39589 5216
rect 39264 5176 39270 5188
rect 39577 5185 39589 5188
rect 39623 5185 39635 5219
rect 39577 5179 39635 5185
rect 40405 5219 40463 5225
rect 40405 5185 40417 5219
rect 40451 5216 40463 5219
rect 40586 5216 40592 5228
rect 40451 5188 40592 5216
rect 40451 5185 40463 5188
rect 40405 5179 40463 5185
rect 40586 5176 40592 5188
rect 40644 5176 40650 5228
rect 40862 5216 40868 5228
rect 40823 5188 40868 5216
rect 40862 5176 40868 5188
rect 40920 5176 40926 5228
rect 37424 5120 38240 5148
rect 38381 5151 38439 5157
rect 37424 5108 37430 5120
rect 38381 5117 38393 5151
rect 38427 5148 38439 5151
rect 38470 5148 38476 5160
rect 38427 5120 38476 5148
rect 38427 5117 38439 5120
rect 38381 5111 38439 5117
rect 38470 5108 38476 5120
rect 38528 5148 38534 5160
rect 40310 5148 40316 5160
rect 38528 5120 40316 5148
rect 38528 5108 38534 5120
rect 40310 5108 40316 5120
rect 40368 5108 40374 5160
rect 41386 5148 41414 5256
rect 42352 5148 42380 5324
rect 43809 5321 43821 5324
rect 43855 5321 43867 5355
rect 43809 5315 43867 5321
rect 42518 5244 42524 5296
rect 42576 5284 42582 5296
rect 42613 5287 42671 5293
rect 42613 5284 42625 5287
rect 42576 5256 42625 5284
rect 42576 5244 42582 5256
rect 42613 5253 42625 5256
rect 42659 5253 42671 5287
rect 42613 5247 42671 5253
rect 47857 5219 47915 5225
rect 47857 5185 47869 5219
rect 47903 5216 47915 5219
rect 47946 5216 47952 5228
rect 47903 5188 47952 5216
rect 47903 5185 47915 5188
rect 47857 5179 47915 5185
rect 47946 5176 47952 5188
rect 48004 5176 48010 5228
rect 42521 5151 42579 5157
rect 42521 5148 42533 5151
rect 41386 5120 42533 5148
rect 42521 5117 42533 5120
rect 42567 5117 42579 5151
rect 42521 5111 42579 5117
rect 43533 5151 43591 5157
rect 43533 5117 43545 5151
rect 43579 5148 43591 5151
rect 43622 5148 43628 5160
rect 43579 5120 43628 5148
rect 43579 5117 43591 5120
rect 43533 5111 43591 5117
rect 43622 5108 43628 5120
rect 43680 5148 43686 5160
rect 43806 5148 43812 5160
rect 43680 5120 43812 5148
rect 43680 5108 43686 5120
rect 43806 5108 43812 5120
rect 43864 5108 43870 5160
rect 24946 5040 24952 5092
rect 25004 5080 25010 5092
rect 48041 5083 48099 5089
rect 48041 5080 48053 5083
rect 25004 5052 48053 5080
rect 25004 5040 25010 5052
rect 48041 5049 48053 5052
rect 48087 5049 48099 5083
rect 48041 5043 48099 5049
rect 18046 4972 18052 5024
rect 18104 5012 18110 5024
rect 18417 5015 18475 5021
rect 18417 5012 18429 5015
rect 18104 4984 18429 5012
rect 18104 4972 18110 4984
rect 18417 4981 18429 4984
rect 18463 4981 18475 5015
rect 18417 4975 18475 4981
rect 21913 5015 21971 5021
rect 21913 4981 21925 5015
rect 21959 5012 21971 5015
rect 22462 5012 22468 5024
rect 21959 4984 22468 5012
rect 21959 4981 21971 4984
rect 21913 4975 21971 4981
rect 22462 4972 22468 4984
rect 22520 4972 22526 5024
rect 22557 5015 22615 5021
rect 22557 4981 22569 5015
rect 22603 5012 22615 5015
rect 22922 5012 22928 5024
rect 22603 4984 22928 5012
rect 22603 4981 22615 4984
rect 22557 4975 22615 4981
rect 22922 4972 22928 4984
rect 22980 4972 22986 5024
rect 40221 5015 40279 5021
rect 40221 4981 40233 5015
rect 40267 5012 40279 5015
rect 40402 5012 40408 5024
rect 40267 4984 40408 5012
rect 40267 4981 40279 4984
rect 40221 4975 40279 4981
rect 40402 4972 40408 4984
rect 40460 4972 40466 5024
rect 40862 5012 40868 5024
rect 40823 4984 40868 5012
rect 40862 4972 40868 4984
rect 40920 4972 40926 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 39206 4808 39212 4820
rect 39167 4780 39212 4808
rect 39206 4768 39212 4780
rect 39264 4768 39270 4820
rect 39298 4768 39304 4820
rect 39356 4808 39362 4820
rect 40862 4808 40868 4820
rect 39356 4780 40868 4808
rect 39356 4768 39362 4780
rect 40862 4768 40868 4780
rect 40920 4768 40926 4820
rect 42518 4808 42524 4820
rect 42479 4780 42524 4808
rect 42518 4768 42524 4780
rect 42576 4768 42582 4820
rect 22189 4743 22247 4749
rect 22189 4709 22201 4743
rect 22235 4740 22247 4743
rect 23658 4740 23664 4752
rect 22235 4712 23664 4740
rect 22235 4709 22247 4712
rect 22189 4703 22247 4709
rect 23658 4700 23664 4712
rect 23716 4700 23722 4752
rect 22833 4675 22891 4681
rect 22833 4641 22845 4675
rect 22879 4672 22891 4675
rect 24394 4672 24400 4684
rect 22879 4644 24400 4672
rect 22879 4641 22891 4644
rect 22833 4635 22891 4641
rect 24394 4632 24400 4644
rect 24452 4632 24458 4684
rect 38470 4672 38476 4684
rect 38431 4644 38476 4672
rect 38470 4632 38476 4644
rect 38528 4632 38534 4684
rect 40218 4672 40224 4684
rect 40179 4644 40224 4672
rect 40218 4632 40224 4644
rect 40276 4632 40282 4684
rect 40402 4672 40408 4684
rect 40363 4644 40408 4672
rect 40402 4632 40408 4644
rect 40460 4632 40466 4684
rect 45370 4632 45376 4684
rect 45428 4672 45434 4684
rect 47581 4675 47639 4681
rect 47581 4672 47593 4675
rect 45428 4644 47593 4672
rect 45428 4632 45434 4644
rect 47581 4641 47593 4644
rect 47627 4641 47639 4675
rect 47581 4635 47639 4641
rect 9490 4604 9496 4616
rect 9451 4576 9496 4604
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4604 18107 4607
rect 18230 4604 18236 4616
rect 18095 4576 18236 4604
rect 18095 4573 18107 4576
rect 18049 4567 18107 4573
rect 18230 4564 18236 4576
rect 18288 4564 18294 4616
rect 19242 4604 19248 4616
rect 19203 4576 19248 4604
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 20073 4607 20131 4613
rect 20073 4573 20085 4607
rect 20119 4573 20131 4607
rect 20073 4567 20131 4573
rect 20165 4607 20223 4613
rect 20165 4573 20177 4607
rect 20211 4604 20223 4607
rect 20809 4607 20867 4613
rect 20809 4604 20821 4607
rect 20211 4576 20821 4604
rect 20211 4573 20223 4576
rect 20165 4567 20223 4573
rect 20809 4573 20821 4576
rect 20855 4573 20867 4607
rect 20809 4567 20867 4573
rect 21453 4607 21511 4613
rect 21453 4573 21465 4607
rect 21499 4604 21511 4607
rect 21910 4604 21916 4616
rect 21499 4576 21916 4604
rect 21499 4573 21511 4576
rect 21453 4567 21511 4573
rect 20088 4536 20116 4567
rect 21910 4564 21916 4576
rect 21968 4564 21974 4616
rect 22094 4604 22100 4616
rect 22055 4576 22100 4604
rect 22094 4564 22100 4576
rect 22152 4564 22158 4616
rect 22462 4564 22468 4616
rect 22520 4604 22526 4616
rect 22741 4607 22799 4613
rect 22741 4604 22753 4607
rect 22520 4576 22753 4604
rect 22520 4564 22526 4576
rect 22741 4573 22753 4576
rect 22787 4573 22799 4607
rect 22741 4567 22799 4573
rect 23474 4564 23480 4616
rect 23532 4604 23538 4616
rect 23569 4607 23627 4613
rect 23569 4604 23581 4607
rect 23532 4576 23581 4604
rect 23532 4564 23538 4576
rect 23569 4573 23581 4576
rect 23615 4573 23627 4607
rect 23569 4567 23627 4573
rect 25498 4564 25504 4616
rect 25556 4604 25562 4616
rect 25777 4607 25835 4613
rect 25777 4604 25789 4607
rect 25556 4576 25789 4604
rect 25556 4564 25562 4576
rect 25777 4573 25789 4576
rect 25823 4573 25835 4607
rect 25777 4567 25835 4573
rect 39117 4607 39175 4613
rect 39117 4573 39129 4607
rect 39163 4604 39175 4607
rect 40126 4604 40132 4616
rect 39163 4576 40132 4604
rect 39163 4573 39175 4576
rect 39117 4567 39175 4573
rect 40126 4564 40132 4576
rect 40184 4564 40190 4616
rect 42705 4607 42763 4613
rect 42705 4573 42717 4607
rect 42751 4604 42763 4607
rect 42886 4604 42892 4616
rect 42751 4576 42892 4604
rect 42751 4573 42763 4576
rect 42705 4567 42763 4573
rect 42886 4564 42892 4576
rect 42944 4564 42950 4616
rect 45002 4564 45008 4616
rect 45060 4604 45066 4616
rect 46661 4607 46719 4613
rect 46661 4604 46673 4607
rect 45060 4576 46673 4604
rect 45060 4564 45066 4576
rect 46661 4573 46673 4576
rect 46707 4573 46719 4607
rect 46661 4567 46719 4573
rect 46842 4564 46848 4616
rect 46900 4604 46906 4616
rect 47305 4607 47363 4613
rect 47305 4604 47317 4607
rect 46900 4576 47317 4604
rect 46900 4564 46906 4576
rect 47305 4573 47317 4576
rect 47351 4573 47363 4607
rect 47305 4567 47363 4573
rect 20990 4536 20996 4548
rect 20088 4508 20996 4536
rect 20990 4496 20996 4508
rect 21048 4496 21054 4548
rect 21545 4539 21603 4545
rect 21545 4505 21557 4539
rect 21591 4536 21603 4539
rect 23014 4536 23020 4548
rect 21591 4508 23020 4536
rect 21591 4505 21603 4508
rect 21545 4499 21603 4505
rect 23014 4496 23020 4508
rect 23072 4496 23078 4548
rect 37274 4496 37280 4548
rect 37332 4536 37338 4548
rect 37461 4539 37519 4545
rect 37461 4536 37473 4539
rect 37332 4508 37473 4536
rect 37332 4496 37338 4508
rect 37461 4505 37473 4508
rect 37507 4505 37519 4539
rect 37461 4499 37519 4505
rect 37550 4496 37556 4548
rect 37608 4536 37614 4548
rect 42061 4539 42119 4545
rect 37608 4508 37653 4536
rect 37608 4496 37614 4508
rect 42061 4505 42073 4539
rect 42107 4536 42119 4539
rect 42150 4536 42156 4548
rect 42107 4508 42156 4536
rect 42107 4505 42119 4508
rect 42061 4499 42119 4505
rect 42150 4496 42156 4508
rect 42208 4536 42214 4548
rect 42610 4536 42616 4548
rect 42208 4508 42616 4536
rect 42208 4496 42214 4508
rect 42610 4496 42616 4508
rect 42668 4496 42674 4548
rect 18138 4468 18144 4480
rect 18099 4440 18144 4468
rect 18138 4428 18144 4440
rect 18196 4428 18202 4480
rect 19334 4468 19340 4480
rect 19295 4440 19340 4468
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 20901 4471 20959 4477
rect 20901 4437 20913 4471
rect 20947 4468 20959 4471
rect 21450 4468 21456 4480
rect 20947 4440 21456 4468
rect 20947 4437 20959 4440
rect 20901 4431 20959 4437
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 23385 4471 23443 4477
rect 23385 4437 23397 4471
rect 23431 4468 23443 4471
rect 24302 4468 24308 4480
rect 23431 4440 24308 4468
rect 23431 4437 23443 4440
rect 23385 4431 23443 4437
rect 24302 4428 24308 4440
rect 24360 4428 24366 4480
rect 46474 4428 46480 4480
rect 46532 4468 46538 4480
rect 46753 4471 46811 4477
rect 46753 4468 46765 4471
rect 46532 4440 46765 4468
rect 46532 4428 46538 4440
rect 46753 4437 46765 4440
rect 46799 4437 46811 4471
rect 46753 4431 46811 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 20990 4264 20996 4276
rect 17276 4236 18552 4264
rect 20951 4236 20996 4264
rect 17276 4224 17282 4236
rect 18138 4196 18144 4208
rect 17880 4168 18144 4196
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 5258 4128 5264 4140
rect 2915 4100 5264 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 8846 4128 8852 4140
rect 8807 4100 8852 4128
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4097 10103 4131
rect 13722 4128 13728 4140
rect 13683 4100 13728 4128
rect 10045 4091 10103 4097
rect 10060 4060 10088 4091
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4128 17371 4131
rect 17880 4128 17908 4168
rect 18138 4156 18144 4168
rect 18196 4156 18202 4208
rect 17359 4100 17908 4128
rect 17359 4097 17371 4100
rect 17313 4091 17371 4097
rect 17954 4088 17960 4140
rect 18012 4128 18018 4140
rect 18012 4100 18057 4128
rect 18012 4088 18018 4100
rect 17405 4063 17463 4069
rect 10060 4032 17356 4060
rect 3418 3952 3424 4004
rect 3476 3992 3482 4004
rect 17218 3992 17224 4004
rect 3476 3964 17224 3992
rect 3476 3952 3482 3964
rect 17218 3952 17224 3964
rect 17276 3952 17282 4004
rect 17328 3992 17356 4032
rect 17405 4029 17417 4063
rect 17451 4060 17463 4063
rect 18322 4060 18328 4072
rect 17451 4032 18328 4060
rect 17451 4029 17463 4032
rect 17405 4023 17463 4029
rect 18322 4020 18328 4032
rect 18380 4020 18386 4072
rect 18524 4060 18552 4236
rect 20990 4224 20996 4236
rect 21048 4224 21054 4276
rect 21910 4264 21916 4276
rect 21871 4236 21916 4264
rect 21910 4224 21916 4236
rect 21968 4224 21974 4276
rect 37277 4267 37335 4273
rect 37277 4233 37289 4267
rect 37323 4264 37335 4267
rect 37458 4264 37464 4276
rect 37323 4236 37464 4264
rect 37323 4233 37335 4236
rect 37277 4227 37335 4233
rect 37458 4224 37464 4236
rect 37516 4224 37522 4276
rect 40586 4224 40592 4276
rect 40644 4264 40650 4276
rect 40865 4267 40923 4273
rect 40865 4264 40877 4267
rect 40644 4236 40877 4264
rect 40644 4224 40650 4236
rect 40865 4233 40877 4236
rect 40911 4233 40923 4267
rect 40865 4227 40923 4233
rect 25225 4199 25283 4205
rect 25225 4196 25237 4199
rect 24964 4168 25237 4196
rect 18966 4128 18972 4140
rect 18927 4100 18972 4128
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19058 4088 19064 4140
rect 19116 4128 19122 4140
rect 19613 4131 19671 4137
rect 19613 4128 19625 4131
rect 19116 4100 19625 4128
rect 19116 4088 19122 4100
rect 19613 4097 19625 4100
rect 19659 4097 19671 4131
rect 20254 4128 20260 4140
rect 20215 4100 20260 4128
rect 19613 4091 19671 4097
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 20901 4131 20959 4137
rect 20901 4097 20913 4131
rect 20947 4128 20959 4131
rect 21358 4128 21364 4140
rect 20947 4100 21364 4128
rect 20947 4097 20959 4100
rect 20901 4091 20959 4097
rect 21358 4088 21364 4100
rect 21416 4088 21422 4140
rect 21450 4088 21456 4140
rect 21508 4128 21514 4140
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 21508 4100 21833 4128
rect 21508 4088 21514 4100
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 21821 4091 21879 4097
rect 22465 4131 22523 4137
rect 22465 4097 22477 4131
rect 22511 4128 22523 4131
rect 23106 4128 23112 4140
rect 22511 4100 22876 4128
rect 23067 4100 23112 4128
rect 22511 4097 22523 4100
rect 22465 4091 22523 4097
rect 18524 4032 21036 4060
rect 18506 3992 18512 4004
rect 17328 3964 18512 3992
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 18598 3952 18604 4004
rect 18656 3992 18662 4004
rect 19705 3995 19763 4001
rect 18656 3964 19196 3992
rect 18656 3952 18662 3964
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1673 3927 1731 3933
rect 1673 3924 1685 3927
rect 1452 3896 1685 3924
rect 1452 3884 1458 3896
rect 1673 3893 1685 3896
rect 1719 3893 1731 3927
rect 2222 3924 2228 3936
rect 2183 3896 2228 3924
rect 1673 3887 1731 3893
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 2958 3924 2964 3936
rect 2919 3896 2964 3924
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 5960 3896 6561 3924
rect 5960 3884 5966 3896
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 6972 3896 7205 3924
rect 6972 3884 6978 3896
rect 7193 3893 7205 3896
rect 7239 3893 7251 3927
rect 7193 3887 7251 3893
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8941 3927 8999 3933
rect 8941 3924 8953 3927
rect 8168 3896 8953 3924
rect 8168 3884 8174 3896
rect 8941 3893 8953 3896
rect 8987 3893 8999 3927
rect 8941 3887 8999 3893
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 10137 3927 10195 3933
rect 10137 3924 10149 3927
rect 9456 3896 10149 3924
rect 9456 3884 9462 3896
rect 10137 3893 10149 3896
rect 10183 3893 10195 3927
rect 10137 3887 10195 3893
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11572 3896 11713 3924
rect 11572 3884 11578 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 13998 3924 14004 3936
rect 13863 3896 14004 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 17494 3884 17500 3936
rect 17552 3924 17558 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17552 3896 18061 3924
rect 17552 3884 17558 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 19061 3927 19119 3933
rect 19061 3924 19073 3927
rect 18840 3896 19073 3924
rect 18840 3884 18846 3896
rect 19061 3893 19073 3896
rect 19107 3893 19119 3927
rect 19168 3924 19196 3964
rect 19705 3961 19717 3995
rect 19751 3992 19763 3995
rect 20806 3992 20812 4004
rect 19751 3964 20812 3992
rect 19751 3961 19763 3964
rect 19705 3955 19763 3961
rect 20806 3952 20812 3964
rect 20864 3952 20870 4004
rect 21008 3992 21036 4032
rect 22848 3992 22876 4100
rect 23106 4088 23112 4100
rect 23164 4088 23170 4140
rect 23198 4088 23204 4140
rect 23256 4128 23262 4140
rect 23753 4131 23811 4137
rect 23256 4100 23301 4128
rect 23256 4088 23262 4100
rect 23753 4097 23765 4131
rect 23799 4128 23811 4131
rect 24486 4128 24492 4140
rect 23799 4100 24492 4128
rect 23799 4097 23811 4100
rect 23753 4091 23811 4097
rect 24486 4088 24492 4100
rect 24544 4088 24550 4140
rect 24854 4088 24860 4140
rect 24912 4128 24918 4140
rect 24964 4128 24992 4168
rect 25225 4165 25237 4168
rect 25271 4165 25283 4199
rect 40034 4196 40040 4208
rect 39995 4168 40040 4196
rect 25225 4159 25283 4165
rect 40034 4156 40040 4168
rect 40092 4156 40098 4208
rect 40494 4196 40500 4208
rect 40455 4168 40500 4196
rect 40494 4156 40500 4168
rect 40552 4156 40558 4208
rect 42794 4156 42800 4208
rect 42852 4196 42858 4208
rect 42889 4199 42947 4205
rect 42889 4196 42901 4199
rect 42852 4168 42901 4196
rect 42852 4156 42858 4168
rect 42889 4165 42901 4168
rect 42935 4165 42947 4199
rect 43806 4196 43812 4208
rect 43767 4168 43812 4196
rect 42889 4159 42947 4165
rect 43806 4156 43812 4168
rect 43864 4156 43870 4208
rect 47762 4196 47768 4208
rect 47723 4168 47768 4196
rect 47762 4156 47768 4168
rect 47820 4156 47826 4208
rect 37461 4131 37519 4137
rect 24912 4100 24992 4128
rect 25976 4100 30052 4128
rect 24912 4088 24918 4100
rect 23842 4060 23848 4072
rect 23803 4032 23848 4060
rect 23842 4020 23848 4032
rect 23900 4020 23906 4072
rect 24946 4020 24952 4072
rect 25004 4060 25010 4072
rect 25133 4063 25191 4069
rect 25133 4060 25145 4063
rect 25004 4032 25145 4060
rect 25004 4020 25010 4032
rect 25133 4029 25145 4032
rect 25179 4060 25191 4063
rect 25976 4060 26004 4100
rect 30024 4072 30052 4100
rect 37461 4097 37473 4131
rect 37507 4128 37519 4131
rect 37734 4128 37740 4140
rect 37507 4100 37740 4128
rect 37507 4097 37519 4100
rect 37461 4091 37519 4097
rect 37734 4088 37740 4100
rect 37792 4088 37798 4140
rect 39577 4131 39635 4137
rect 39577 4097 39589 4131
rect 39623 4128 39635 4131
rect 40218 4128 40224 4140
rect 39623 4100 40224 4128
rect 39623 4097 39635 4100
rect 39577 4091 39635 4097
rect 40218 4088 40224 4100
rect 40276 4128 40282 4140
rect 40681 4131 40739 4137
rect 40681 4128 40693 4131
rect 40276 4100 40693 4128
rect 40276 4088 40282 4100
rect 40681 4097 40693 4100
rect 40727 4097 40739 4131
rect 46750 4128 46756 4140
rect 46711 4100 46756 4128
rect 40681 4091 40739 4097
rect 46750 4088 46756 4100
rect 46808 4088 46814 4140
rect 25179 4032 26004 4060
rect 26053 4063 26111 4069
rect 25179 4029 25191 4032
rect 25133 4023 25191 4029
rect 26053 4029 26065 4063
rect 26099 4060 26111 4063
rect 26234 4060 26240 4072
rect 26099 4032 26240 4060
rect 26099 4029 26111 4032
rect 26053 4023 26111 4029
rect 26234 4020 26240 4032
rect 26292 4060 26298 4072
rect 26878 4060 26884 4072
rect 26292 4032 26884 4060
rect 26292 4020 26298 4032
rect 26878 4020 26884 4032
rect 26936 4020 26942 4072
rect 30006 4020 30012 4072
rect 30064 4060 30070 4072
rect 37274 4060 37280 4072
rect 30064 4032 37280 4060
rect 30064 4020 30070 4032
rect 37274 4020 37280 4032
rect 37332 4060 37338 4072
rect 39393 4063 39451 4069
rect 39393 4060 39405 4063
rect 37332 4032 39405 4060
rect 37332 4020 37338 4032
rect 39393 4029 39405 4032
rect 39439 4060 39451 4063
rect 39942 4060 39948 4072
rect 39439 4032 39948 4060
rect 39439 4029 39451 4032
rect 39393 4023 39451 4029
rect 39942 4020 39948 4032
rect 40000 4060 40006 4072
rect 42797 4063 42855 4069
rect 42797 4060 42809 4063
rect 40000 4032 42809 4060
rect 40000 4020 40006 4032
rect 42797 4029 42809 4032
rect 42843 4060 42855 4063
rect 45278 4060 45284 4072
rect 42843 4032 45284 4060
rect 42843 4029 42855 4032
rect 42797 4023 42855 4029
rect 45278 4020 45284 4032
rect 45336 4020 45342 4072
rect 48041 4063 48099 4069
rect 48041 4060 48053 4063
rect 45526 4032 48053 4060
rect 29546 3992 29552 4004
rect 21008 3964 22692 3992
rect 22848 3964 29552 3992
rect 20070 3924 20076 3936
rect 19168 3896 20076 3924
rect 19061 3887 19119 3893
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20349 3927 20407 3933
rect 20349 3893 20361 3927
rect 20395 3924 20407 3927
rect 20898 3924 20904 3936
rect 20395 3896 20904 3924
rect 20395 3893 20407 3896
rect 20349 3887 20407 3893
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 22462 3884 22468 3936
rect 22520 3924 22526 3936
rect 22557 3927 22615 3933
rect 22557 3924 22569 3927
rect 22520 3896 22569 3924
rect 22520 3884 22526 3896
rect 22557 3893 22569 3896
rect 22603 3893 22615 3927
rect 22664 3924 22692 3964
rect 29546 3952 29552 3964
rect 29604 3952 29610 4004
rect 45526 3992 45554 4032
rect 48041 4029 48053 4032
rect 48087 4029 48099 4063
rect 48041 4023 48099 4029
rect 46937 3995 46995 4001
rect 46937 3992 46949 3995
rect 31726 3964 45554 3992
rect 46124 3964 46949 3992
rect 23566 3924 23572 3936
rect 22664 3896 23572 3924
rect 22557 3887 22615 3893
rect 23566 3884 23572 3896
rect 23624 3884 23630 3936
rect 30926 3884 30932 3936
rect 30984 3924 30990 3936
rect 31726 3924 31754 3964
rect 30984 3896 31754 3924
rect 30984 3884 30990 3896
rect 32674 3884 32680 3936
rect 32732 3924 32738 3936
rect 46124 3924 46152 3964
rect 46937 3961 46949 3964
rect 46983 3961 46995 3995
rect 46937 3955 46995 3961
rect 46290 3924 46296 3936
rect 32732 3896 46152 3924
rect 46251 3896 46296 3924
rect 32732 3884 32738 3896
rect 46290 3884 46296 3896
rect 46348 3884 46354 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 17129 3723 17187 3729
rect 17129 3689 17141 3723
rect 17175 3720 17187 3723
rect 18230 3720 18236 3732
rect 17175 3692 18236 3720
rect 17175 3689 17187 3692
rect 17129 3683 17187 3689
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 20162 3720 20168 3732
rect 18748 3692 20168 3720
rect 18748 3680 18754 3692
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20254 3680 20260 3732
rect 20312 3720 20318 3732
rect 20901 3723 20959 3729
rect 20901 3720 20913 3723
rect 20312 3692 20913 3720
rect 20312 3680 20318 3692
rect 20901 3689 20913 3692
rect 20947 3689 20959 3723
rect 20901 3683 20959 3689
rect 21358 3680 21364 3732
rect 21416 3720 21422 3732
rect 21545 3723 21603 3729
rect 21545 3720 21557 3723
rect 21416 3692 21557 3720
rect 21416 3680 21422 3692
rect 21545 3689 21557 3692
rect 21591 3689 21603 3723
rect 21545 3683 21603 3689
rect 23106 3680 23112 3732
rect 23164 3720 23170 3732
rect 23753 3723 23811 3729
rect 23753 3720 23765 3723
rect 23164 3692 23765 3720
rect 23164 3680 23170 3692
rect 23753 3689 23765 3692
rect 23799 3689 23811 3723
rect 24486 3720 24492 3732
rect 24447 3692 24492 3720
rect 23753 3683 23811 3689
rect 24486 3680 24492 3692
rect 24544 3680 24550 3732
rect 24578 3680 24584 3732
rect 24636 3720 24642 3732
rect 30926 3720 30932 3732
rect 24636 3692 30932 3720
rect 24636 3680 24642 3692
rect 30926 3680 30932 3692
rect 30984 3680 30990 3732
rect 31110 3680 31116 3732
rect 31168 3720 31174 3732
rect 31168 3692 31754 3720
rect 31168 3680 31174 3692
rect 658 3612 664 3664
rect 716 3652 722 3664
rect 716 3624 2360 3652
rect 716 3612 722 3624
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 2222 3584 2228 3596
rect 1627 3556 2228 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2332 3593 2360 3624
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 18138 3652 18144 3664
rect 5316 3624 11744 3652
rect 5316 3612 5322 3624
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3553 2375 3587
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 2317 3547 2375 3553
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 9217 3587 9275 3593
rect 9217 3553 9229 3587
rect 9263 3584 9275 3587
rect 9490 3584 9496 3596
rect 9263 3556 9496 3584
rect 9263 3553 9275 3556
rect 9217 3547 9275 3553
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9640 3556 9689 3584
rect 9640 3544 9646 3556
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 2792 3488 3985 3516
rect 2038 3408 2044 3460
rect 2096 3448 2102 3460
rect 2792 3448 2820 3488
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 5258 3516 5264 3528
rect 5219 3488 5264 3516
rect 3973 3479 4031 3485
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 7984 3488 8401 3516
rect 7984 3476 7990 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 2096 3420 2820 3448
rect 5353 3451 5411 3457
rect 2096 3408 2102 3420
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 6089 3451 6147 3457
rect 6089 3448 6101 3451
rect 5399 3420 6101 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 6089 3417 6101 3420
rect 6135 3417 6147 3451
rect 9398 3448 9404 3460
rect 9359 3420 9404 3448
rect 6089 3411 6147 3417
rect 9398 3408 9404 3420
rect 9456 3408 9462 3460
rect 11716 3448 11744 3624
rect 13648 3624 18144 3652
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3516 12035 3519
rect 13648 3516 13676 3624
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 18322 3612 18328 3664
rect 18380 3652 18386 3664
rect 26694 3652 26700 3664
rect 18380 3624 26700 3652
rect 18380 3612 18386 3624
rect 26694 3612 26700 3624
rect 26752 3612 26758 3664
rect 31726 3652 31754 3692
rect 32858 3680 32864 3732
rect 32916 3720 32922 3732
rect 39298 3720 39304 3732
rect 32916 3692 39304 3720
rect 32916 3680 32922 3692
rect 39298 3680 39304 3692
rect 39356 3680 39362 3732
rect 40126 3720 40132 3732
rect 40087 3692 40132 3720
rect 40126 3680 40132 3692
rect 40184 3680 40190 3732
rect 33778 3652 33784 3664
rect 26804 3624 27200 3652
rect 31726 3624 33784 3652
rect 26804 3584 26832 3624
rect 14384 3556 26832 3584
rect 26881 3587 26939 3593
rect 12023 3488 13676 3516
rect 12023 3485 12035 3488
rect 11977 3479 12035 3485
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13872 3488 14289 3516
rect 13872 3476 13878 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14384 3448 14412 3556
rect 26881 3553 26893 3587
rect 26927 3553 26939 3587
rect 27172 3584 27200 3624
rect 33778 3612 33784 3624
rect 33836 3612 33842 3664
rect 34054 3612 34060 3664
rect 34112 3652 34118 3664
rect 42518 3652 42524 3664
rect 34112 3624 42524 3652
rect 34112 3612 34118 3624
rect 42518 3612 42524 3624
rect 42576 3612 42582 3664
rect 46566 3652 46572 3664
rect 45526 3624 46572 3652
rect 45526 3584 45554 3624
rect 46566 3612 46572 3624
rect 46624 3612 46630 3664
rect 46290 3584 46296 3596
rect 27172 3556 34008 3584
rect 26881 3547 26939 3553
rect 33980 3550 34008 3556
rect 34072 3556 45554 3584
rect 46251 3556 46296 3584
rect 34072 3550 34100 3556
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3516 17095 3519
rect 17494 3516 17500 3528
rect 17083 3488 17500 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3516 17739 3519
rect 17770 3516 17776 3528
rect 17727 3488 17776 3516
rect 17727 3485 17739 3488
rect 17681 3479 17739 3485
rect 17770 3476 17776 3488
rect 17828 3476 17834 3528
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 19334 3516 19340 3528
rect 18371 3488 19340 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 19444 3488 19533 3516
rect 11716 3420 14412 3448
rect 16114 3408 16120 3460
rect 16172 3448 16178 3460
rect 18230 3448 18236 3460
rect 16172 3420 18236 3448
rect 16172 3408 16178 3420
rect 18230 3408 18236 3420
rect 18288 3408 18294 3460
rect 18417 3451 18475 3457
rect 18417 3417 18429 3451
rect 18463 3448 18475 3451
rect 18966 3448 18972 3460
rect 18463 3420 18972 3448
rect 18463 3417 18475 3420
rect 18417 3411 18475 3417
rect 18966 3408 18972 3420
rect 19024 3408 19030 3460
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 12069 3383 12127 3389
rect 12069 3380 12081 3383
rect 11756 3352 12081 3380
rect 11756 3340 11762 3352
rect 12069 3349 12081 3352
rect 12115 3349 12127 3383
rect 12069 3343 12127 3349
rect 17402 3340 17408 3392
rect 17460 3380 17466 3392
rect 17773 3383 17831 3389
rect 17773 3380 17785 3383
rect 17460 3352 17785 3380
rect 17460 3340 17466 3352
rect 17773 3349 17785 3352
rect 17819 3349 17831 3383
rect 17773 3343 17831 3349
rect 18138 3340 18144 3392
rect 18196 3380 18202 3392
rect 19444 3380 19472 3488
rect 19521 3485 19533 3488
rect 19567 3516 19579 3519
rect 20346 3516 20352 3528
rect 19567 3488 20208 3516
rect 20307 3488 20352 3516
rect 19567 3485 19579 3488
rect 19521 3479 19579 3485
rect 20180 3448 20208 3488
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 20806 3516 20812 3528
rect 20767 3488 20812 3516
rect 20806 3476 20812 3488
rect 20864 3476 20870 3528
rect 20898 3476 20904 3528
rect 20956 3516 20962 3528
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 20956 3488 21465 3516
rect 20956 3476 20962 3488
rect 21453 3485 21465 3488
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 22278 3476 22284 3528
rect 22336 3516 22342 3528
rect 22557 3519 22615 3525
rect 22557 3516 22569 3519
rect 22336 3488 22569 3516
rect 22336 3476 22342 3488
rect 22557 3485 22569 3488
rect 22603 3485 22615 3519
rect 23014 3516 23020 3528
rect 22975 3488 23020 3516
rect 22557 3479 22615 3485
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 23658 3516 23664 3528
rect 23619 3488 23664 3516
rect 23658 3476 23664 3488
rect 23716 3476 23722 3528
rect 24394 3516 24400 3528
rect 24355 3488 24400 3516
rect 24394 3476 24400 3488
rect 24452 3476 24458 3528
rect 25498 3516 25504 3528
rect 25459 3488 25504 3516
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 20714 3448 20720 3460
rect 20180 3420 20720 3448
rect 20714 3408 20720 3420
rect 20772 3408 20778 3460
rect 22094 3408 22100 3460
rect 22152 3448 22158 3460
rect 23109 3451 23167 3457
rect 23109 3448 23121 3451
rect 22152 3420 23121 3448
rect 22152 3408 22158 3420
rect 23109 3417 23121 3420
rect 23155 3417 23167 3451
rect 23109 3411 23167 3417
rect 25685 3451 25743 3457
rect 25685 3417 25697 3451
rect 25731 3417 25743 3451
rect 25685 3411 25743 3417
rect 18196 3352 19472 3380
rect 19613 3383 19671 3389
rect 18196 3340 18202 3352
rect 19613 3349 19625 3383
rect 19659 3380 19671 3383
rect 19978 3380 19984 3392
rect 19659 3352 19984 3380
rect 19659 3349 19671 3352
rect 19613 3343 19671 3349
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 20622 3340 20628 3392
rect 20680 3380 20686 3392
rect 24578 3380 24584 3392
rect 20680 3352 24584 3380
rect 20680 3340 20686 3352
rect 24578 3340 24584 3352
rect 24636 3340 24642 3392
rect 25700 3380 25728 3411
rect 25774 3408 25780 3460
rect 25832 3448 25838 3460
rect 26896 3448 26924 3547
rect 33045 3519 33103 3525
rect 33045 3485 33057 3519
rect 33091 3516 33103 3519
rect 33870 3516 33876 3528
rect 33091 3488 33732 3516
rect 33831 3488 33876 3516
rect 33091 3485 33103 3488
rect 33045 3479 33103 3485
rect 25832 3420 26924 3448
rect 25832 3408 25838 3420
rect 32858 3380 32864 3392
rect 25700 3352 32864 3380
rect 32858 3340 32864 3352
rect 32916 3340 32922 3392
rect 33134 3380 33140 3392
rect 33095 3352 33140 3380
rect 33134 3340 33140 3352
rect 33192 3340 33198 3392
rect 33704 3380 33732 3488
rect 33870 3476 33876 3488
rect 33928 3476 33934 3528
rect 33980 3522 34100 3550
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 46474 3584 46480 3596
rect 46435 3556 46480 3584
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 40034 3516 40040 3528
rect 39995 3488 40040 3516
rect 40034 3476 40040 3488
rect 40092 3476 40098 3528
rect 40770 3516 40776 3528
rect 40731 3488 40776 3516
rect 40770 3476 40776 3488
rect 40828 3476 40834 3528
rect 43073 3519 43131 3525
rect 43073 3516 43085 3519
rect 42168 3488 43085 3516
rect 39666 3408 39672 3460
rect 39724 3448 39730 3460
rect 40957 3451 41015 3457
rect 40957 3448 40969 3451
rect 39724 3420 40969 3448
rect 39724 3408 39730 3420
rect 40957 3417 40969 3420
rect 41003 3417 41015 3451
rect 40957 3411 41015 3417
rect 41138 3380 41144 3392
rect 33704 3352 41144 3380
rect 41138 3340 41144 3352
rect 41196 3380 41202 3392
rect 42168 3380 42196 3488
rect 43073 3485 43085 3488
rect 43119 3485 43131 3519
rect 43898 3516 43904 3528
rect 43859 3488 43904 3516
rect 43073 3479 43131 3485
rect 43898 3476 43904 3488
rect 43956 3476 43962 3528
rect 45186 3516 45192 3528
rect 45147 3488 45192 3516
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 45649 3519 45707 3525
rect 45649 3485 45661 3519
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 42610 3448 42616 3460
rect 42571 3420 42616 3448
rect 42610 3408 42616 3420
rect 42668 3408 42674 3460
rect 45664 3448 45692 3479
rect 47486 3448 47492 3460
rect 45664 3420 47492 3448
rect 47486 3408 47492 3420
rect 47544 3408 47550 3460
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 41196 3352 42196 3380
rect 41196 3340 41202 3352
rect 43070 3340 43076 3392
rect 43128 3380 43134 3392
rect 43165 3383 43223 3389
rect 43165 3380 43177 3383
rect 43128 3352 43177 3380
rect 43128 3340 43134 3352
rect 43165 3349 43177 3352
rect 43211 3349 43223 3383
rect 43165 3343 43223 3349
rect 45370 3340 45376 3392
rect 45428 3380 45434 3392
rect 45741 3383 45799 3389
rect 45741 3380 45753 3383
rect 45428 3352 45753 3380
rect 45428 3340 45434 3352
rect 45741 3349 45753 3352
rect 45787 3349 45799 3383
rect 45741 3343 45799 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 37458 3176 37464 3188
rect 8904 3148 37464 3176
rect 8904 3136 8910 3148
rect 37458 3136 37464 3148
rect 37516 3136 37522 3188
rect 37734 3176 37740 3188
rect 37695 3148 37740 3176
rect 37734 3136 37740 3148
rect 37792 3136 37798 3188
rect 39666 3176 39672 3188
rect 39627 3148 39672 3176
rect 39666 3136 39672 3148
rect 39724 3136 39730 3188
rect 40770 3136 40776 3188
rect 40828 3176 40834 3188
rect 40957 3179 41015 3185
rect 40957 3176 40969 3179
rect 40828 3148 40969 3176
rect 40828 3136 40834 3148
rect 40957 3145 40969 3148
rect 41003 3145 41015 3179
rect 40957 3139 41015 3145
rect 47670 3136 47676 3188
rect 47728 3176 47734 3188
rect 47857 3179 47915 3185
rect 47857 3176 47869 3179
rect 47728 3148 47869 3176
rect 47728 3136 47734 3148
rect 47857 3145 47869 3148
rect 47903 3145 47915 3179
rect 47857 3139 47915 3145
rect 2225 3111 2283 3117
rect 2225 3077 2237 3111
rect 2271 3108 2283 3111
rect 2958 3108 2964 3120
rect 2271 3080 2964 3108
rect 2271 3077 2283 3080
rect 2225 3071 2283 3077
rect 2958 3068 2964 3080
rect 3016 3068 3022 3120
rect 8110 3108 8116 3120
rect 8071 3080 8116 3108
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 11698 3108 11704 3120
rect 11659 3080 11704 3108
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 13998 3108 14004 3120
rect 13959 3080 14004 3108
rect 13998 3068 14004 3080
rect 14056 3068 14062 3120
rect 17770 3108 17776 3120
rect 17731 3080 17776 3108
rect 17770 3068 17776 3080
rect 17828 3068 17834 3120
rect 18877 3111 18935 3117
rect 18877 3077 18889 3111
rect 18923 3108 18935 3111
rect 19058 3108 19064 3120
rect 18923 3080 19064 3108
rect 18923 3077 18935 3080
rect 18877 3071 18935 3077
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 19613 3111 19671 3117
rect 19613 3108 19625 3111
rect 19352 3080 19625 3108
rect 2038 3040 2044 3052
rect 1999 3012 2044 3040
rect 2038 3000 2044 3012
rect 2096 3000 2102 3052
rect 6638 3040 6644 3052
rect 6599 3012 6644 3040
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 7926 3040 7932 3052
rect 7887 3012 7932 3040
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 13814 3040 13820 3052
rect 13775 3012 13820 3040
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 17681 3043 17739 3049
rect 17681 3040 17693 3043
rect 16853 3003 16911 3009
rect 17236 3012 17693 3040
rect 2958 2972 2964 2984
rect 2919 2944 2964 2972
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 7800 2944 8401 2972
rect 7800 2932 7806 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11020 2944 11989 2972
rect 11020 2932 11026 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14240 2944 14289 2972
rect 14240 2932 14246 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 15194 2932 15200 2984
rect 15252 2972 15258 2984
rect 16761 2975 16819 2981
rect 16761 2972 16773 2975
rect 15252 2944 16773 2972
rect 15252 2932 15258 2944
rect 16761 2941 16773 2944
rect 16807 2941 16819 2975
rect 16761 2935 16819 2941
rect 6730 2836 6736 2848
rect 6691 2808 6736 2836
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9582 2836 9588 2848
rect 9088 2808 9588 2836
rect 9088 2796 9094 2808
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 16868 2836 16896 3003
rect 17236 2981 17264 3012
rect 17681 3009 17693 3012
rect 17727 3009 17739 3043
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 17681 3003 17739 3009
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 19352 2904 19380 3080
rect 19613 3077 19625 3080
rect 19659 3077 19671 3111
rect 19613 3071 19671 3077
rect 19702 3068 19708 3120
rect 19760 3108 19766 3120
rect 21082 3108 21088 3120
rect 19760 3080 21088 3108
rect 19760 3068 19766 3080
rect 21082 3068 21088 3080
rect 21140 3068 21146 3120
rect 22462 3108 22468 3120
rect 22423 3080 22468 3108
rect 22462 3068 22468 3080
rect 22520 3068 22526 3120
rect 24302 3068 24308 3120
rect 24360 3108 24366 3120
rect 25133 3111 25191 3117
rect 25133 3108 25145 3111
rect 24360 3080 25145 3108
rect 24360 3068 24366 3080
rect 25133 3077 25145 3080
rect 25179 3077 25191 3111
rect 25133 3071 25191 3077
rect 25225 3111 25283 3117
rect 25225 3077 25237 3111
rect 25271 3108 25283 3111
rect 26050 3108 26056 3120
rect 25271 3080 26056 3108
rect 25271 3077 25283 3080
rect 25225 3071 25283 3077
rect 26050 3068 26056 3080
rect 26108 3068 26114 3120
rect 26145 3111 26203 3117
rect 26145 3077 26157 3111
rect 26191 3108 26203 3111
rect 26234 3108 26240 3120
rect 26191 3080 26240 3108
rect 26191 3077 26203 3080
rect 26145 3071 26203 3077
rect 26234 3068 26240 3080
rect 26292 3068 26298 3120
rect 26694 3068 26700 3120
rect 26752 3108 26758 3120
rect 32214 3108 32220 3120
rect 26752 3080 32220 3108
rect 26752 3068 26758 3080
rect 32214 3068 32220 3080
rect 32272 3068 32278 3120
rect 33134 3108 33140 3120
rect 33095 3080 33140 3108
rect 33134 3068 33140 3080
rect 33192 3068 33198 3120
rect 42610 3108 42616 3120
rect 38626 3080 42616 3108
rect 22278 3040 22284 3052
rect 22239 3012 22284 3040
rect 22278 3000 22284 3012
rect 22336 3000 22342 3052
rect 27154 3040 27160 3052
rect 25976 3012 26234 3040
rect 27115 3012 27160 3040
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2972 19487 2975
rect 20346 2972 20352 2984
rect 19475 2944 20352 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 20346 2932 20352 2944
rect 20404 2932 20410 2984
rect 20441 2975 20499 2981
rect 20441 2941 20453 2975
rect 20487 2941 20499 2975
rect 20441 2935 20499 2941
rect 19886 2904 19892 2916
rect 19352 2876 19892 2904
rect 19886 2864 19892 2876
rect 19944 2864 19950 2916
rect 19978 2864 19984 2916
rect 20036 2904 20042 2916
rect 20456 2904 20484 2935
rect 22554 2932 22560 2984
rect 22612 2972 22618 2984
rect 22741 2975 22799 2981
rect 22741 2972 22753 2975
rect 22612 2944 22753 2972
rect 22612 2932 22618 2944
rect 22741 2941 22753 2944
rect 22787 2941 22799 2975
rect 22741 2935 22799 2941
rect 20036 2876 20484 2904
rect 20036 2864 20042 2876
rect 20530 2864 20536 2916
rect 20588 2904 20594 2916
rect 24854 2904 24860 2916
rect 20588 2876 24860 2904
rect 20588 2864 20594 2876
rect 24854 2864 24860 2876
rect 24912 2864 24918 2916
rect 25130 2864 25136 2916
rect 25188 2904 25194 2916
rect 25774 2904 25780 2916
rect 25188 2876 25780 2904
rect 25188 2864 25194 2876
rect 25774 2864 25780 2876
rect 25832 2864 25838 2916
rect 25976 2836 26004 3012
rect 26206 2904 26234 3012
rect 27154 3000 27160 3012
rect 27212 3000 27218 3052
rect 32953 3043 33011 3049
rect 32953 3009 32965 3043
rect 32999 3009 33011 3043
rect 32953 3003 33011 3009
rect 37277 3043 37335 3049
rect 37277 3009 37289 3043
rect 37323 3040 37335 3043
rect 37550 3040 37556 3052
rect 37323 3012 37556 3040
rect 37323 3009 37335 3012
rect 37277 3003 37335 3009
rect 32968 2972 32996 3003
rect 37550 3000 37556 3012
rect 37608 3000 37614 3052
rect 33502 2972 33508 2984
rect 32968 2944 33364 2972
rect 33463 2944 33508 2972
rect 33336 2904 33364 2944
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 38626 2972 38654 3080
rect 42610 3068 42616 3080
rect 42668 3068 42674 3120
rect 43070 3108 43076 3120
rect 43031 3080 43076 3108
rect 43070 3068 43076 3080
rect 43128 3068 43134 3120
rect 45370 3108 45376 3120
rect 45331 3080 45376 3108
rect 45370 3068 45376 3080
rect 45428 3068 45434 3120
rect 39209 3043 39267 3049
rect 39209 3009 39221 3043
rect 39255 3009 39267 3043
rect 39209 3003 39267 3009
rect 39853 3043 39911 3049
rect 39853 3009 39865 3043
rect 39899 3040 39911 3043
rect 40586 3040 40592 3052
rect 39899 3012 40592 3040
rect 39899 3009 39911 3012
rect 39853 3003 39911 3009
rect 33980 2944 38654 2972
rect 39224 2972 39252 3003
rect 40586 3000 40592 3012
rect 40644 3000 40650 3052
rect 41230 3000 41236 3052
rect 41288 3040 41294 3052
rect 41601 3043 41659 3049
rect 41601 3040 41613 3043
rect 41288 3012 41613 3040
rect 41288 3000 41294 3012
rect 41601 3009 41613 3012
rect 41647 3009 41659 3043
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 41601 3003 41659 3009
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 47765 3043 47823 3049
rect 47765 3009 47777 3043
rect 47811 3040 47823 3043
rect 48314 3040 48320 3052
rect 47811 3012 48320 3040
rect 47811 3009 47823 3012
rect 47765 3003 47823 3009
rect 48314 3000 48320 3012
rect 48372 3000 48378 3052
rect 39942 2972 39948 2984
rect 39224 2944 39948 2972
rect 33870 2904 33876 2916
rect 26206 2876 28994 2904
rect 33336 2876 33876 2904
rect 16868 2808 26004 2836
rect 26050 2796 26056 2848
rect 26108 2836 26114 2848
rect 26973 2839 27031 2845
rect 26973 2836 26985 2839
rect 26108 2808 26985 2836
rect 26108 2796 26114 2808
rect 26973 2805 26985 2808
rect 27019 2805 27031 2839
rect 28966 2836 28994 2876
rect 33870 2864 33876 2876
rect 33928 2864 33934 2916
rect 33980 2836 34008 2944
rect 39942 2932 39948 2944
rect 40000 2932 40006 2984
rect 40034 2932 40040 2984
rect 40092 2972 40098 2984
rect 40313 2975 40371 2981
rect 40313 2972 40325 2975
rect 40092 2944 40325 2972
rect 40092 2932 40098 2944
rect 40313 2941 40325 2944
rect 40359 2941 40371 2975
rect 40313 2935 40371 2941
rect 40402 2932 40408 2984
rect 40460 2972 40466 2984
rect 40497 2975 40555 2981
rect 40497 2972 40509 2975
rect 40460 2944 40509 2972
rect 40460 2932 40466 2944
rect 40497 2941 40509 2944
rect 40543 2972 40555 2975
rect 42889 2975 42947 2981
rect 40543 2944 41460 2972
rect 40543 2941 40555 2944
rect 40497 2935 40555 2941
rect 39025 2907 39083 2913
rect 39025 2873 39037 2907
rect 39071 2904 39083 2907
rect 40218 2904 40224 2916
rect 39071 2876 40224 2904
rect 39071 2873 39083 2876
rect 39025 2867 39083 2873
rect 40218 2864 40224 2876
rect 40276 2864 40282 2916
rect 41432 2913 41460 2944
rect 42889 2941 42901 2975
rect 42935 2972 42947 2975
rect 43898 2972 43904 2984
rect 42935 2944 43904 2972
rect 42935 2941 42947 2944
rect 42889 2935 42947 2941
rect 43898 2932 43904 2944
rect 43956 2932 43962 2984
rect 43993 2975 44051 2981
rect 43993 2941 44005 2975
rect 44039 2941 44051 2975
rect 43993 2935 44051 2941
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 41417 2907 41475 2913
rect 41417 2873 41429 2907
rect 41463 2873 41475 2907
rect 41417 2867 41475 2873
rect 43162 2864 43168 2916
rect 43220 2904 43226 2916
rect 44008 2904 44036 2935
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 43220 2876 44036 2904
rect 43220 2864 43226 2876
rect 37366 2836 37372 2848
rect 28966 2808 34008 2836
rect 37327 2808 37372 2836
rect 26973 2799 27031 2805
rect 37366 2796 37372 2808
rect 37424 2796 37430 2848
rect 37458 2796 37464 2848
rect 37516 2836 37522 2848
rect 45646 2836 45652 2848
rect 37516 2808 45652 2836
rect 37516 2796 37522 2808
rect 45646 2796 45652 2808
rect 45704 2796 45710 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 9125 2635 9183 2641
rect 5276 2604 9076 2632
rect 5276 2505 5304 2604
rect 6914 2564 6920 2576
rect 6564 2536 6920 2564
rect 6564 2505 6592 2536
rect 6914 2524 6920 2536
rect 6972 2524 6978 2576
rect 9048 2564 9076 2604
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9306 2632 9312 2644
rect 9171 2604 9312 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 15194 2632 15200 2644
rect 12406 2604 15200 2632
rect 12406 2564 12434 2604
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 17310 2632 17316 2644
rect 16546 2604 17316 2632
rect 9048 2536 12434 2564
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2465 5319 2499
rect 5261 2459 5319 2465
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2465 6607 2499
rect 6730 2496 6736 2508
rect 6691 2468 6736 2496
rect 6549 2459 6607 2465
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 7098 2496 7104 2508
rect 7059 2468 7104 2496
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 16546 2496 16574 2604
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17497 2635 17555 2641
rect 17497 2601 17509 2635
rect 17543 2632 17555 2635
rect 17954 2632 17960 2644
rect 17543 2604 17960 2632
rect 17543 2601 17555 2604
rect 17497 2595 17555 2601
rect 17954 2592 17960 2604
rect 18012 2592 18018 2644
rect 18141 2635 18199 2641
rect 18141 2601 18153 2635
rect 18187 2632 18199 2635
rect 19242 2632 19248 2644
rect 18187 2604 19248 2632
rect 18187 2601 18199 2604
rect 18141 2595 18199 2601
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 20456 2604 24164 2632
rect 16853 2567 16911 2573
rect 16853 2533 16865 2567
rect 16899 2564 16911 2567
rect 20456 2564 20484 2604
rect 16899 2536 20484 2564
rect 20533 2567 20591 2573
rect 16899 2533 16911 2536
rect 16853 2527 16911 2533
rect 20533 2533 20545 2567
rect 20579 2564 20591 2567
rect 21266 2564 21272 2576
rect 20579 2536 21272 2564
rect 20579 2533 20591 2536
rect 20533 2527 20591 2533
rect 21266 2524 21272 2536
rect 21324 2524 21330 2576
rect 24136 2564 24164 2604
rect 24210 2592 24216 2644
rect 24268 2632 24274 2644
rect 24673 2635 24731 2641
rect 24673 2632 24685 2635
rect 24268 2604 24685 2632
rect 24268 2592 24274 2604
rect 24673 2601 24685 2604
rect 24719 2601 24731 2635
rect 24673 2595 24731 2601
rect 25501 2635 25559 2641
rect 25501 2601 25513 2635
rect 25547 2632 25559 2635
rect 26234 2632 26240 2644
rect 25547 2604 26240 2632
rect 25547 2601 25559 2604
rect 25501 2595 25559 2601
rect 26234 2592 26240 2604
rect 26292 2592 26298 2644
rect 26329 2635 26387 2641
rect 26329 2601 26341 2635
rect 26375 2632 26387 2635
rect 26375 2604 27568 2632
rect 26375 2601 26387 2604
rect 26329 2595 26387 2601
rect 25685 2567 25743 2573
rect 24136 2536 24808 2564
rect 24780 2496 24808 2536
rect 25685 2533 25697 2567
rect 25731 2564 25743 2567
rect 27154 2564 27160 2576
rect 25731 2536 27160 2564
rect 25731 2533 25743 2536
rect 25685 2527 25743 2533
rect 27154 2524 27160 2536
rect 27212 2524 27218 2576
rect 27430 2496 27436 2508
rect 7248 2468 16574 2496
rect 20088 2468 24716 2496
rect 24780 2468 27436 2496
rect 7248 2456 7254 2468
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5166 2428 5172 2440
rect 5031 2400 5172 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8536 2400 8953 2428
rect 8536 2388 8542 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 12406 2400 15792 2428
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 1360 2332 1869 2360
rect 1360 2320 1366 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 2777 2363 2835 2369
rect 2777 2360 2789 2363
rect 2648 2332 2789 2360
rect 2648 2320 2654 2332
rect 2777 2329 2789 2332
rect 2823 2329 2835 2363
rect 2777 2323 2835 2329
rect 3145 2363 3203 2369
rect 3145 2329 3157 2363
rect 3191 2360 3203 2363
rect 12406 2360 12434 2400
rect 3191 2332 12434 2360
rect 3191 2329 3203 2332
rect 3145 2323 3203 2329
rect 15470 2320 15476 2372
rect 15528 2360 15534 2372
rect 15657 2363 15715 2369
rect 15657 2360 15669 2363
rect 15528 2332 15669 2360
rect 15528 2320 15534 2332
rect 15657 2329 15669 2332
rect 15703 2329 15715 2363
rect 15764 2360 15792 2400
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16172 2400 16681 2428
rect 16172 2388 16178 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 17402 2428 17408 2440
rect 17363 2400 17408 2428
rect 16669 2391 16727 2397
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 18046 2428 18052 2440
rect 18007 2400 18052 2428
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 20088 2360 20116 2468
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 22097 2431 22155 2437
rect 22097 2428 22109 2431
rect 21315 2400 22109 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 22097 2397 22109 2400
rect 22143 2397 22155 2431
rect 22922 2428 22928 2440
rect 22883 2400 22928 2428
rect 22097 2391 22155 2397
rect 22922 2388 22928 2400
rect 22980 2388 22986 2440
rect 23293 2431 23351 2437
rect 23293 2397 23305 2431
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 15764 2332 20116 2360
rect 20349 2363 20407 2369
rect 15657 2323 15715 2329
rect 20349 2329 20361 2363
rect 20395 2360 20407 2363
rect 20622 2360 20628 2372
rect 20395 2332 20628 2360
rect 20395 2329 20407 2332
rect 20349 2323 20407 2329
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 21085 2363 21143 2369
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 21910 2360 21916 2372
rect 21131 2332 21916 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 21910 2320 21916 2332
rect 21968 2320 21974 2372
rect 2130 2292 2136 2304
rect 2091 2264 2136 2292
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 7190 2292 7196 2304
rect 4120 2264 7196 2292
rect 4120 2252 4126 2264
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 15746 2292 15752 2304
rect 15707 2264 15752 2292
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 17310 2252 17316 2304
rect 17368 2292 17374 2304
rect 22830 2292 22836 2304
rect 17368 2264 22836 2292
rect 17368 2252 17374 2264
rect 22830 2252 22836 2264
rect 22888 2252 22894 2304
rect 23308 2292 23336 2391
rect 24486 2320 24492 2372
rect 24544 2360 24550 2372
rect 24581 2363 24639 2369
rect 24581 2360 24593 2363
rect 24544 2332 24593 2360
rect 24544 2320 24550 2332
rect 24581 2329 24593 2332
rect 24627 2329 24639 2363
rect 24688 2360 24716 2468
rect 27430 2456 27436 2468
rect 27488 2456 27494 2508
rect 27540 2496 27568 2604
rect 28350 2592 28356 2644
rect 28408 2632 28414 2644
rect 28629 2635 28687 2641
rect 28629 2632 28641 2635
rect 28408 2604 28641 2632
rect 28408 2592 28414 2604
rect 28629 2601 28641 2604
rect 28675 2601 28687 2635
rect 29730 2632 29736 2644
rect 29691 2604 29736 2632
rect 28629 2595 28687 2601
rect 29730 2592 29736 2604
rect 29788 2592 29794 2644
rect 32306 2592 32312 2644
rect 32364 2632 32370 2644
rect 35618 2632 35624 2644
rect 32364 2604 35624 2632
rect 32364 2592 32370 2604
rect 35618 2592 35624 2604
rect 35676 2592 35682 2644
rect 36354 2632 36360 2644
rect 36315 2604 36360 2632
rect 36354 2592 36360 2604
rect 36412 2592 36418 2644
rect 40405 2635 40463 2641
rect 40405 2601 40417 2635
rect 40451 2601 40463 2635
rect 40586 2632 40592 2644
rect 40547 2604 40592 2632
rect 40405 2595 40463 2601
rect 27617 2567 27675 2573
rect 27617 2533 27629 2567
rect 27663 2564 27675 2567
rect 30098 2564 30104 2576
rect 27663 2536 30104 2564
rect 27663 2533 27675 2536
rect 27617 2527 27675 2533
rect 30098 2524 30104 2536
rect 30156 2524 30162 2576
rect 35894 2564 35900 2576
rect 32324 2536 35900 2564
rect 27540 2468 32168 2496
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 24912 2400 25237 2428
rect 24912 2388 24918 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2428 26203 2431
rect 26418 2428 26424 2440
rect 26191 2400 26424 2428
rect 26191 2397 26203 2400
rect 26145 2391 26203 2397
rect 26418 2388 26424 2400
rect 26476 2388 26482 2440
rect 27706 2428 27712 2440
rect 26988 2400 27712 2428
rect 26988 2360 27016 2400
rect 27706 2388 27712 2400
rect 27764 2388 27770 2440
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29696 2400 29929 2428
rect 29696 2388 29702 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 32140 2428 32168 2468
rect 32324 2428 32352 2536
rect 35894 2524 35900 2536
rect 35952 2524 35958 2576
rect 35986 2524 35992 2576
rect 36044 2564 36050 2576
rect 40420 2564 40448 2595
rect 40586 2592 40592 2604
rect 40644 2592 40650 2644
rect 42521 2635 42579 2641
rect 42521 2601 42533 2635
rect 42567 2601 42579 2635
rect 42886 2632 42892 2644
rect 42847 2604 42892 2632
rect 42521 2595 42579 2601
rect 40494 2564 40500 2576
rect 36044 2536 39436 2564
rect 40420 2536 40500 2564
rect 36044 2524 36050 2536
rect 33686 2456 33692 2508
rect 33744 2496 33750 2508
rect 38381 2499 38439 2505
rect 38381 2496 38393 2499
rect 33744 2468 38393 2496
rect 33744 2456 33750 2468
rect 38381 2465 38393 2468
rect 38427 2465 38439 2499
rect 38381 2459 38439 2465
rect 39301 2499 39359 2505
rect 39301 2465 39313 2499
rect 39347 2465 39359 2499
rect 39408 2496 39436 2536
rect 40494 2524 40500 2536
rect 40552 2524 40558 2576
rect 41325 2567 41383 2573
rect 41325 2533 41337 2567
rect 41371 2564 41383 2567
rect 42426 2564 42432 2576
rect 41371 2536 42432 2564
rect 41371 2533 41383 2536
rect 41325 2527 41383 2533
rect 42426 2524 42432 2536
rect 42484 2524 42490 2576
rect 42536 2496 42564 2595
rect 42886 2592 42892 2604
rect 42944 2592 42950 2644
rect 46477 2499 46535 2505
rect 46477 2496 46489 2499
rect 39408 2468 42564 2496
rect 43548 2468 46489 2496
rect 39301 2459 39359 2465
rect 32140 2400 32352 2428
rect 29917 2391 29975 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 39316 2428 39344 2459
rect 35713 2391 35771 2397
rect 37568 2400 39344 2428
rect 40037 2431 40095 2437
rect 24688 2332 27016 2360
rect 24581 2323 24639 2329
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 27120 2332 27445 2360
rect 27120 2320 27126 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28537 2363 28595 2369
rect 28537 2360 28549 2363
rect 28408 2332 28549 2360
rect 28408 2320 28414 2332
rect 28537 2329 28549 2332
rect 28583 2329 28595 2363
rect 28537 2323 28595 2329
rect 29730 2320 29736 2372
rect 29788 2360 29794 2372
rect 35986 2360 35992 2372
rect 29788 2332 35992 2360
rect 29788 2320 29794 2332
rect 35986 2320 35992 2332
rect 36044 2320 36050 2372
rect 36078 2320 36084 2372
rect 36136 2360 36142 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 36136 2332 36277 2360
rect 36136 2320 36142 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 36265 2323 36323 2329
rect 24946 2292 24952 2304
rect 23308 2264 24952 2292
rect 24946 2252 24952 2264
rect 25004 2252 25010 2304
rect 26234 2252 26240 2304
rect 26292 2292 26298 2304
rect 35529 2295 35587 2301
rect 35529 2292 35541 2295
rect 26292 2264 35541 2292
rect 26292 2252 26298 2264
rect 35529 2261 35541 2264
rect 35575 2261 35587 2295
rect 35529 2255 35587 2261
rect 35618 2252 35624 2304
rect 35676 2292 35682 2304
rect 37568 2292 37596 2400
rect 40037 2397 40049 2431
rect 40083 2428 40095 2431
rect 40218 2428 40224 2440
rect 40083 2400 40224 2428
rect 40083 2397 40095 2400
rect 40037 2391 40095 2397
rect 40218 2388 40224 2400
rect 40276 2388 40282 2440
rect 40402 2428 40408 2440
rect 40363 2400 40408 2428
rect 40402 2388 40408 2400
rect 40460 2388 40466 2440
rect 40586 2388 40592 2440
rect 40644 2428 40650 2440
rect 41141 2431 41199 2437
rect 41141 2428 41153 2431
rect 40644 2400 41153 2428
rect 40644 2388 40650 2400
rect 41141 2397 41153 2400
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 42429 2431 42487 2437
rect 42429 2397 42441 2431
rect 42475 2428 42487 2431
rect 42794 2428 42800 2440
rect 42475 2400 42800 2428
rect 42475 2397 42487 2400
rect 42429 2391 42487 2397
rect 42794 2388 42800 2400
rect 42852 2428 42858 2440
rect 43548 2428 43576 2468
rect 46477 2465 46489 2468
rect 46523 2465 46535 2499
rect 47854 2496 47860 2508
rect 47815 2468 47860 2496
rect 46477 2459 46535 2465
rect 47854 2456 47860 2468
rect 47912 2456 47918 2508
rect 42852 2400 43576 2428
rect 43625 2431 43683 2437
rect 42852 2388 42858 2400
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43806 2428 43812 2440
rect 43671 2400 43812 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 43901 2431 43959 2437
rect 43901 2397 43913 2431
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 46201 2431 46259 2437
rect 46201 2397 46213 2431
rect 46247 2428 46259 2431
rect 47026 2428 47032 2440
rect 46247 2400 47032 2428
rect 46247 2397 46259 2400
rect 46201 2391 46259 2397
rect 38010 2320 38016 2372
rect 38068 2360 38074 2372
rect 38197 2363 38255 2369
rect 38197 2360 38209 2363
rect 38068 2332 38209 2360
rect 38068 2320 38074 2332
rect 38197 2329 38209 2332
rect 38243 2329 38255 2363
rect 38197 2323 38255 2329
rect 39117 2363 39175 2369
rect 39117 2329 39129 2363
rect 39163 2360 39175 2363
rect 39298 2360 39304 2372
rect 39163 2332 39304 2360
rect 39163 2329 39175 2332
rect 39117 2323 39175 2329
rect 39298 2320 39304 2332
rect 39356 2320 39362 2372
rect 43916 2360 43944 2391
rect 47026 2388 47032 2400
rect 47084 2388 47090 2440
rect 47673 2431 47731 2437
rect 47673 2397 47685 2431
rect 47719 2428 47731 2431
rect 48038 2428 48044 2440
rect 47719 2400 48044 2428
rect 47719 2397 47731 2400
rect 47673 2391 47731 2397
rect 48038 2388 48044 2400
rect 48096 2388 48102 2440
rect 39408 2332 43944 2360
rect 45373 2363 45431 2369
rect 35676 2264 37596 2292
rect 35676 2252 35682 2264
rect 37642 2252 37648 2304
rect 37700 2292 37706 2304
rect 39408 2292 39436 2332
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46382 2360 46388 2372
rect 45419 2332 46388 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46382 2320 46388 2332
rect 46440 2320 46446 2372
rect 37700 2264 39436 2292
rect 37700 2252 37706 2264
rect 41322 2252 41328 2304
rect 41380 2292 41386 2304
rect 45465 2295 45523 2301
rect 45465 2292 45477 2295
rect 41380 2264 45477 2292
rect 41380 2252 41386 2264
rect 45465 2261 45477 2264
rect 45511 2261 45523 2295
rect 45465 2255 45523 2261
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 27430 2048 27436 2100
rect 27488 2088 27494 2100
rect 32030 2088 32036 2100
rect 27488 2060 32036 2088
rect 27488 2048 27494 2060
rect 32030 2048 32036 2060
rect 32088 2048 32094 2100
rect 35894 2048 35900 2100
rect 35952 2088 35958 2100
rect 40678 2088 40684 2100
rect 35952 2060 40684 2088
rect 35952 2048 35958 2060
rect 40678 2048 40684 2060
rect 40736 2048 40742 2100
rect 22370 1980 22376 2032
rect 22428 2020 22434 2032
rect 41322 2020 41328 2032
rect 22428 1992 41328 2020
rect 22428 1980 22434 1992
rect 41322 1980 41328 1992
rect 41380 1980 41386 2032
rect 2130 1912 2136 1964
rect 2188 1952 2194 1964
rect 26970 1952 26976 1964
rect 2188 1924 26976 1952
rect 2188 1912 2194 1924
rect 26970 1912 26976 1924
rect 27028 1912 27034 1964
rect 15746 1844 15752 1896
rect 15804 1884 15810 1896
rect 37366 1884 37372 1896
rect 15804 1856 37372 1884
rect 15804 1844 15810 1856
rect 37366 1844 37372 1856
rect 37424 1844 37430 1896
<< via1 >>
rect 13360 47540 13412 47592
rect 20536 47540 20588 47592
rect 6644 47472 6696 47524
rect 37372 47472 37424 47524
rect 2044 47404 2096 47456
rect 38200 47404 38252 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 13360 47243 13412 47252
rect 13360 47209 13369 47243
rect 13369 47209 13403 47243
rect 13403 47209 13412 47243
rect 13360 47200 13412 47209
rect 38200 47200 38252 47252
rect 40500 47200 40552 47252
rect 29000 47132 29052 47184
rect 29828 47132 29880 47184
rect 33692 47132 33744 47184
rect 2044 47107 2096 47116
rect 2044 47073 2053 47107
rect 2053 47073 2087 47107
rect 2087 47073 2096 47107
rect 2044 47064 2096 47073
rect 6644 47107 6696 47116
rect 6644 47073 6653 47107
rect 6653 47073 6687 47107
rect 6687 47073 6696 47107
rect 6644 47064 6696 47073
rect 1952 46996 2004 47048
rect 3240 46996 3292 47048
rect 4712 47039 4764 47048
rect 4712 47005 4721 47039
rect 4721 47005 4755 47039
rect 4755 47005 4764 47039
rect 4712 46996 4764 47005
rect 5816 46996 5868 47048
rect 2596 46860 2648 46912
rect 3056 46928 3108 46980
rect 4068 46971 4120 46980
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 7288 47039 7340 47048
rect 7288 47005 7297 47039
rect 7297 47005 7331 47039
rect 7331 47005 7340 47039
rect 7288 46996 7340 47005
rect 9036 46996 9088 47048
rect 11612 47039 11664 47048
rect 11612 47005 11621 47039
rect 11621 47005 11655 47039
rect 11655 47005 11664 47039
rect 11612 46996 11664 47005
rect 12256 46996 12308 47048
rect 12900 46996 12952 47048
rect 16488 46996 16540 47048
rect 16948 47039 17000 47048
rect 16948 47005 16957 47039
rect 16957 47005 16991 47039
rect 16991 47005 17000 47039
rect 16948 46996 17000 47005
rect 11704 46928 11756 46980
rect 12440 46928 12492 46980
rect 14740 46971 14792 46980
rect 7472 46903 7524 46912
rect 7472 46869 7481 46903
rect 7481 46869 7515 46903
rect 7515 46869 7524 46903
rect 7472 46860 7524 46869
rect 13544 46860 13596 46912
rect 14740 46937 14749 46971
rect 14749 46937 14783 46971
rect 14783 46937 14792 46971
rect 14740 46928 14792 46937
rect 18696 47064 18748 47116
rect 19984 47064 20036 47116
rect 20352 47039 20404 47048
rect 18696 46971 18748 46980
rect 18696 46937 18705 46971
rect 18705 46937 18739 46971
rect 18739 46937 18748 46971
rect 18696 46928 18748 46937
rect 20352 47005 20361 47039
rect 20361 47005 20395 47039
rect 20395 47005 20404 47039
rect 20352 46996 20404 47005
rect 24860 47039 24912 47048
rect 24860 47005 24869 47039
rect 24869 47005 24903 47039
rect 24903 47005 24912 47039
rect 24860 46996 24912 47005
rect 25504 47039 25556 47048
rect 25504 47005 25513 47039
rect 25513 47005 25547 47039
rect 25547 47005 25556 47039
rect 25504 46996 25556 47005
rect 28908 47064 28960 47116
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 30932 46996 30984 47048
rect 38200 46996 38252 47048
rect 42708 47039 42760 47048
rect 42708 47005 42717 47039
rect 42717 47005 42751 47039
rect 42751 47005 42760 47039
rect 42708 46996 42760 47005
rect 44456 47064 44508 47116
rect 48320 47064 48372 47116
rect 43812 46996 43864 47048
rect 45192 47039 45244 47048
rect 45192 47005 45201 47039
rect 45201 47005 45235 47039
rect 45235 47005 45244 47039
rect 45192 46996 45244 47005
rect 47676 46996 47728 47048
rect 28724 46971 28776 46980
rect 28724 46937 28733 46971
rect 28733 46937 28767 46971
rect 28767 46937 28776 46971
rect 28724 46928 28776 46937
rect 31392 46928 31444 46980
rect 39304 46860 39356 46912
rect 40408 46928 40460 46980
rect 44364 46928 44416 46980
rect 45468 46928 45520 46980
rect 41880 46860 41932 46912
rect 42892 46860 42944 46912
rect 43352 46903 43404 46912
rect 43352 46869 43361 46903
rect 43361 46869 43395 46903
rect 43395 46869 43404 46903
rect 43352 46860 43404 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 1860 46631 1912 46640
rect 1860 46597 1869 46631
rect 1869 46597 1903 46631
rect 1903 46597 1912 46631
rect 1860 46588 1912 46597
rect 24860 46588 24912 46640
rect 43168 46588 43220 46640
rect 47032 46631 47084 46640
rect 47032 46597 47041 46631
rect 47041 46597 47075 46631
rect 47075 46597 47084 46631
rect 47032 46588 47084 46597
rect 38200 46563 38252 46572
rect 38200 46529 38209 46563
rect 38209 46529 38243 46563
rect 38243 46529 38252 46563
rect 38200 46520 38252 46529
rect 42708 46563 42760 46572
rect 42708 46529 42717 46563
rect 42717 46529 42751 46563
rect 42751 46529 42760 46563
rect 42708 46520 42760 46529
rect 47952 46563 48004 46572
rect 47952 46529 47961 46563
rect 47961 46529 47995 46563
rect 47995 46529 48004 46563
rect 47952 46520 48004 46529
rect 3884 46452 3936 46504
rect 3976 46452 4028 46504
rect 14188 46452 14240 46504
rect 14280 46495 14332 46504
rect 14280 46461 14289 46495
rect 14289 46461 14323 46495
rect 14323 46461 14332 46495
rect 19432 46495 19484 46504
rect 14280 46452 14332 46461
rect 19432 46461 19441 46495
rect 19441 46461 19475 46495
rect 19475 46461 19484 46495
rect 19432 46452 19484 46461
rect 20260 46452 20312 46504
rect 20628 46495 20680 46504
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 25136 46495 25188 46504
rect 25136 46461 25145 46495
rect 25145 46461 25179 46495
rect 25179 46461 25188 46495
rect 25136 46452 25188 46461
rect 32404 46495 32456 46504
rect 32404 46461 32413 46495
rect 32413 46461 32447 46495
rect 32447 46461 32456 46495
rect 32404 46452 32456 46461
rect 33324 46452 33376 46504
rect 38384 46495 38436 46504
rect 4620 46384 4672 46436
rect 32220 46384 32272 46436
rect 38384 46461 38393 46495
rect 38393 46461 38427 46495
rect 38427 46461 38436 46495
rect 38384 46452 38436 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 43812 46452 43864 46504
rect 45376 46495 45428 46504
rect 45376 46461 45385 46495
rect 45385 46461 45419 46495
rect 45419 46461 45428 46495
rect 45376 46452 45428 46461
rect 45560 46384 45612 46436
rect 2320 46316 2372 46368
rect 2872 46359 2924 46368
rect 2872 46325 2881 46359
rect 2881 46325 2915 46359
rect 2915 46325 2924 46359
rect 2872 46316 2924 46325
rect 10508 46316 10560 46368
rect 20812 46316 20864 46368
rect 41420 46316 41472 46368
rect 47860 46316 47912 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3884 46155 3936 46164
rect 3884 46121 3893 46155
rect 3893 46121 3927 46155
rect 3927 46121 3936 46155
rect 3884 46112 3936 46121
rect 4620 46155 4672 46164
rect 4620 46121 4629 46155
rect 4629 46121 4663 46155
rect 4663 46121 4672 46155
rect 4620 46112 4672 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 19432 46112 19484 46164
rect 24768 46112 24820 46164
rect 32404 46112 32456 46164
rect 38384 46155 38436 46164
rect 38384 46121 38393 46155
rect 38393 46121 38427 46155
rect 38427 46121 38436 46155
rect 38384 46112 38436 46121
rect 43812 46155 43864 46164
rect 43812 46121 43821 46155
rect 43821 46121 43855 46155
rect 43855 46121 43864 46155
rect 43812 46112 43864 46121
rect 10508 46019 10560 46028
rect 10508 45985 10517 46019
rect 10517 45985 10551 46019
rect 10551 45985 10560 46019
rect 10508 45976 10560 45985
rect 10968 45976 11020 46028
rect 3148 45908 3200 45960
rect 20812 46019 20864 46028
rect 20812 45985 20821 46019
rect 20821 45985 20855 46019
rect 20855 45985 20864 46019
rect 20812 45976 20864 45985
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 25504 45976 25556 46028
rect 41420 46019 41472 46028
rect 24860 45908 24912 45960
rect 10692 45883 10744 45892
rect 2964 45815 3016 45824
rect 2964 45781 2973 45815
rect 2973 45781 3007 45815
rect 3007 45781 3016 45815
rect 2964 45772 3016 45781
rect 10692 45849 10701 45883
rect 10701 45849 10735 45883
rect 10735 45849 10744 45883
rect 10692 45840 10744 45849
rect 20996 45883 21048 45892
rect 20996 45849 21005 45883
rect 21005 45849 21039 45883
rect 21039 45849 21048 45883
rect 20996 45840 21048 45849
rect 25412 45883 25464 45892
rect 25412 45849 25421 45883
rect 25421 45849 25455 45883
rect 25455 45849 25464 45883
rect 25412 45840 25464 45849
rect 10600 45772 10652 45824
rect 25780 45772 25832 45824
rect 41420 45985 41429 46019
rect 41429 45985 41463 46019
rect 41463 45985 41472 46019
rect 41420 45976 41472 45985
rect 42524 46019 42576 46028
rect 42524 45985 42533 46019
rect 42533 45985 42567 46019
rect 42567 45985 42576 46019
rect 42524 45976 42576 45985
rect 40316 45908 40368 45960
rect 45836 45976 45888 46028
rect 46756 45976 46808 46028
rect 48136 46019 48188 46028
rect 48136 45985 48145 46019
rect 48145 45985 48179 46019
rect 48179 45985 48188 46019
rect 48136 45976 48188 45985
rect 45744 45908 45796 45960
rect 41604 45883 41656 45892
rect 41604 45849 41613 45883
rect 41613 45849 41647 45883
rect 41647 45849 41656 45883
rect 41604 45840 41656 45849
rect 46940 45840 46992 45892
rect 27344 45772 27396 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 10692 45611 10744 45620
rect 10692 45577 10701 45611
rect 10701 45577 10735 45611
rect 10735 45577 10744 45611
rect 10692 45568 10744 45577
rect 15936 45568 15988 45620
rect 17408 45568 17460 45620
rect 20260 45568 20312 45620
rect 20996 45611 21048 45620
rect 20996 45577 21005 45611
rect 21005 45577 21039 45611
rect 21039 45577 21048 45611
rect 20996 45568 21048 45577
rect 25412 45611 25464 45620
rect 25412 45577 25421 45611
rect 25421 45577 25455 45611
rect 25455 45577 25464 45611
rect 25412 45568 25464 45577
rect 45100 45568 45152 45620
rect 2964 45500 3016 45552
rect 33324 45543 33376 45552
rect 10600 45475 10652 45484
rect 10600 45441 10609 45475
rect 10609 45441 10643 45475
rect 10643 45441 10652 45475
rect 33324 45509 33333 45543
rect 33333 45509 33367 45543
rect 33367 45509 33376 45543
rect 33324 45500 33376 45509
rect 41604 45500 41656 45552
rect 46848 45543 46900 45552
rect 10600 45432 10652 45441
rect 2872 45364 2924 45416
rect 20812 45432 20864 45484
rect 24860 45432 24912 45484
rect 25320 45475 25372 45484
rect 25320 45441 25329 45475
rect 25329 45441 25363 45475
rect 25363 45441 25372 45475
rect 25320 45432 25372 45441
rect 40960 45475 41012 45484
rect 2780 45296 2832 45348
rect 40960 45441 40969 45475
rect 40969 45441 41003 45475
rect 41003 45441 41012 45475
rect 40960 45432 41012 45441
rect 43812 45475 43864 45484
rect 43812 45441 43821 45475
rect 43821 45441 43855 45475
rect 43855 45441 43864 45475
rect 43812 45432 43864 45441
rect 38660 45407 38712 45416
rect 38660 45373 38669 45407
rect 38669 45373 38703 45407
rect 38703 45373 38712 45407
rect 38660 45364 38712 45373
rect 38844 45407 38896 45416
rect 38844 45373 38853 45407
rect 38853 45373 38887 45407
rect 38887 45373 38896 45407
rect 38844 45364 38896 45373
rect 39856 45407 39908 45416
rect 39856 45373 39865 45407
rect 39865 45373 39899 45407
rect 39899 45373 39908 45407
rect 39856 45364 39908 45373
rect 44456 45407 44508 45416
rect 44456 45373 44465 45407
rect 44465 45373 44499 45407
rect 44499 45373 44508 45407
rect 44456 45364 44508 45373
rect 46848 45509 46857 45543
rect 46857 45509 46891 45543
rect 46891 45509 46900 45543
rect 46848 45500 46900 45509
rect 47492 45432 47544 45484
rect 38752 45296 38804 45348
rect 45468 45296 45520 45348
rect 36268 45228 36320 45280
rect 41420 45228 41472 45280
rect 43444 45228 43496 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 38844 45067 38896 45076
rect 38844 45033 38853 45067
rect 38853 45033 38887 45067
rect 38887 45033 38896 45067
rect 38844 45024 38896 45033
rect 44456 45067 44508 45076
rect 44456 45033 44465 45067
rect 44465 45033 44499 45067
rect 44499 45033 44508 45067
rect 44456 45024 44508 45033
rect 45376 45024 45428 45076
rect 41420 44931 41472 44940
rect 41420 44897 41429 44931
rect 41429 44897 41463 44931
rect 41463 44897 41472 44931
rect 41420 44888 41472 44897
rect 42892 44931 42944 44940
rect 42892 44897 42901 44931
rect 42901 44897 42935 44931
rect 42935 44897 42944 44931
rect 42892 44888 42944 44897
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 28080 44820 28132 44872
rect 38752 44863 38804 44872
rect 38752 44829 38761 44863
rect 38761 44829 38795 44863
rect 38795 44829 38804 44863
rect 38752 44820 38804 44829
rect 45008 44863 45060 44872
rect 45008 44829 45017 44863
rect 45017 44829 45051 44863
rect 45051 44829 45060 44863
rect 45008 44820 45060 44829
rect 45836 44820 45888 44872
rect 46296 44863 46348 44872
rect 46296 44829 46305 44863
rect 46305 44829 46339 44863
rect 46339 44829 46348 44863
rect 46296 44820 46348 44829
rect 41604 44795 41656 44804
rect 41604 44761 41613 44795
rect 41613 44761 41647 44795
rect 41647 44761 41656 44795
rect 41604 44752 41656 44761
rect 38660 44684 38712 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 41604 44523 41656 44532
rect 41604 44489 41613 44523
rect 41613 44489 41647 44523
rect 41647 44489 41656 44523
rect 41604 44480 41656 44489
rect 46940 44523 46992 44532
rect 46940 44489 46949 44523
rect 46949 44489 46983 44523
rect 46983 44489 46992 44523
rect 46940 44480 46992 44489
rect 45560 44344 45612 44396
rect 46296 44344 46348 44396
rect 46848 44387 46900 44396
rect 46848 44353 46857 44387
rect 46857 44353 46891 44387
rect 46891 44353 46900 44387
rect 46848 44344 46900 44353
rect 47492 44344 47544 44396
rect 47308 44276 47360 44328
rect 45836 44140 45888 44192
rect 46572 44140 46624 44192
rect 47676 44183 47728 44192
rect 47676 44149 47685 44183
rect 47685 44149 47719 44183
rect 47719 44149 47728 44183
rect 47676 44140 47728 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 45192 43936 45244 43988
rect 47676 43800 47728 43852
rect 48228 43800 48280 43852
rect 46296 43775 46348 43784
rect 46296 43741 46305 43775
rect 46305 43741 46339 43775
rect 46339 43741 46348 43775
rect 46296 43732 46348 43741
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 46296 43256 46348 43308
rect 1492 43188 1544 43240
rect 46756 43188 46808 43240
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 46296 42687 46348 42696
rect 46296 42653 46305 42687
rect 46305 42653 46339 42687
rect 46339 42653 46348 42687
rect 46296 42644 46348 42653
rect 47676 42576 47728 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 47676 42347 47728 42356
rect 47676 42313 47685 42347
rect 47685 42313 47719 42347
rect 47719 42313 47728 42347
rect 47676 42304 47728 42313
rect 46296 42168 46348 42220
rect 47308 42168 47360 42220
rect 1400 41964 1452 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 47676 41624 47728 41676
rect 48136 41599 48188 41608
rect 48136 41565 48145 41599
rect 48145 41565 48179 41599
rect 48179 41565 48188 41599
rect 48136 41556 48188 41565
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 46940 41488 46992 41540
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 46940 41259 46992 41268
rect 46940 41225 46949 41259
rect 46949 41225 46983 41259
rect 46983 41225 46992 41259
rect 46940 41216 46992 41225
rect 2136 41123 2188 41132
rect 2136 41089 2145 41123
rect 2145 41089 2179 41123
rect 2179 41089 2188 41123
rect 2136 41080 2188 41089
rect 46848 41123 46900 41132
rect 46848 41089 46857 41123
rect 46857 41089 46891 41123
rect 46891 41089 46900 41123
rect 46848 41080 46900 41089
rect 47952 41123 48004 41132
rect 47952 41089 47961 41123
rect 47961 41089 47995 41123
rect 47995 41089 48004 41123
rect 47952 41080 48004 41089
rect 48044 40919 48096 40928
rect 48044 40885 48053 40919
rect 48053 40885 48087 40919
rect 48087 40885 48096 40919
rect 48044 40876 48096 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47676 40715 47728 40724
rect 47676 40681 47685 40715
rect 47685 40681 47719 40715
rect 47719 40681 47728 40715
rect 47676 40672 47728 40681
rect 1400 40511 1452 40520
rect 1400 40477 1409 40511
rect 1409 40477 1443 40511
rect 1443 40477 1452 40511
rect 1400 40468 1452 40477
rect 1676 40332 1728 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 46296 39788 46348 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 40776 39448 40828 39500
rect 40960 39448 41012 39500
rect 46296 39491 46348 39500
rect 46296 39457 46305 39491
rect 46305 39457 46339 39491
rect 46339 39457 46348 39491
rect 46296 39448 46348 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 40132 39380 40184 39432
rect 46940 39312 46992 39364
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 46940 39083 46992 39092
rect 46940 39049 46949 39083
rect 46949 39049 46983 39083
rect 46983 39049 46992 39083
rect 46940 39040 46992 39049
rect 3516 38972 3568 39024
rect 7564 38972 7616 39024
rect 40132 38947 40184 38956
rect 40132 38913 40141 38947
rect 40141 38913 40175 38947
rect 40175 38913 40184 38947
rect 40132 38904 40184 38913
rect 46756 38904 46808 38956
rect 47676 38947 47728 38956
rect 47676 38913 47685 38947
rect 47685 38913 47719 38947
rect 47719 38913 47728 38947
rect 47676 38904 47728 38913
rect 3332 38836 3384 38888
rect 3516 38836 3568 38888
rect 40316 38836 40368 38888
rect 44180 38836 44232 38888
rect 45468 38836 45520 38888
rect 45652 38768 45704 38820
rect 46848 38768 46900 38820
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 41328 38360 41380 38412
rect 45008 38360 45060 38412
rect 44180 38292 44232 38344
rect 46296 38335 46348 38344
rect 46296 38301 46305 38335
rect 46305 38301 46339 38335
rect 46339 38301 46348 38335
rect 46296 38292 46348 38301
rect 40132 38224 40184 38276
rect 47676 38224 47728 38276
rect 48136 38267 48188 38276
rect 48136 38233 48145 38267
rect 48145 38233 48179 38267
rect 48179 38233 48188 38267
rect 48136 38224 48188 38233
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 47676 37995 47728 38004
rect 47676 37961 47685 37995
rect 47685 37961 47719 37995
rect 47719 37961 47728 37995
rect 47676 37952 47728 37961
rect 40132 37859 40184 37868
rect 40132 37825 40141 37859
rect 40141 37825 40175 37859
rect 40175 37825 40184 37859
rect 40132 37816 40184 37825
rect 47584 37859 47636 37868
rect 20720 37748 20772 37800
rect 47584 37825 47593 37859
rect 47593 37825 47627 37859
rect 47627 37825 47636 37859
rect 47584 37816 47636 37825
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 46296 37408 46348 37460
rect 1952 37204 2004 37256
rect 12440 37204 12492 37256
rect 40132 37247 40184 37256
rect 40132 37213 40141 37247
rect 40141 37213 40175 37247
rect 40175 37213 40184 37247
rect 40132 37204 40184 37213
rect 27528 37136 27580 37188
rect 40316 37136 40368 37188
rect 25780 37068 25832 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 27344 36907 27396 36916
rect 27344 36873 27353 36907
rect 27353 36873 27387 36907
rect 27387 36873 27396 36907
rect 27344 36864 27396 36873
rect 25320 36796 25372 36848
rect 40316 36864 40368 36916
rect 40684 36864 40736 36916
rect 1952 36771 2004 36780
rect 1952 36737 1961 36771
rect 1961 36737 1995 36771
rect 1995 36737 2004 36771
rect 1952 36728 2004 36737
rect 2872 36660 2924 36712
rect 2964 36703 3016 36712
rect 2964 36669 2973 36703
rect 2973 36669 3007 36703
rect 3007 36669 3016 36703
rect 2964 36660 3016 36669
rect 25688 36728 25740 36780
rect 26332 36660 26384 36712
rect 27528 36703 27580 36712
rect 27528 36669 27537 36703
rect 27537 36669 27571 36703
rect 27571 36669 27580 36703
rect 27528 36660 27580 36669
rect 22376 36524 22428 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2872 36363 2924 36372
rect 2872 36329 2881 36363
rect 2881 36329 2915 36363
rect 2915 36329 2924 36363
rect 2872 36320 2924 36329
rect 6644 36116 6696 36168
rect 37096 36184 37148 36236
rect 24400 36159 24452 36168
rect 24400 36125 24409 36159
rect 24409 36125 24443 36159
rect 24443 36125 24452 36159
rect 24400 36116 24452 36125
rect 28172 36116 28224 36168
rect 33416 36159 33468 36168
rect 33416 36125 33425 36159
rect 33425 36125 33459 36159
rect 33459 36125 33468 36159
rect 33416 36116 33468 36125
rect 22376 36091 22428 36100
rect 22376 36057 22385 36091
rect 22385 36057 22419 36091
rect 22419 36057 22428 36091
rect 22376 36048 22428 36057
rect 22836 36048 22888 36100
rect 24952 36048 25004 36100
rect 25136 36048 25188 36100
rect 25688 35980 25740 36032
rect 26148 36023 26200 36032
rect 26148 35989 26157 36023
rect 26157 35989 26191 36023
rect 26191 35989 26200 36023
rect 26148 35980 26200 35989
rect 28540 35980 28592 36032
rect 33324 35980 33376 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 22836 35776 22888 35828
rect 24952 35776 25004 35828
rect 22376 35708 22428 35760
rect 29920 35776 29972 35828
rect 33416 35776 33468 35828
rect 33692 35819 33744 35828
rect 33692 35785 33701 35819
rect 33701 35785 33735 35819
rect 33735 35785 33744 35819
rect 33692 35776 33744 35785
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 22008 35640 22060 35692
rect 26148 35708 26200 35760
rect 29276 35708 29328 35760
rect 30656 35708 30708 35760
rect 20536 35572 20588 35624
rect 28540 35640 28592 35692
rect 25780 35615 25832 35624
rect 25780 35581 25789 35615
rect 25789 35581 25823 35615
rect 25823 35581 25832 35615
rect 25780 35572 25832 35581
rect 25596 35504 25648 35556
rect 26240 35572 26292 35624
rect 27160 35615 27212 35624
rect 27160 35581 27169 35615
rect 27169 35581 27203 35615
rect 27203 35581 27212 35615
rect 27160 35572 27212 35581
rect 28448 35572 28500 35624
rect 1400 35479 1452 35488
rect 1400 35445 1409 35479
rect 1409 35445 1443 35479
rect 1443 35445 1452 35479
rect 1400 35436 1452 35445
rect 24584 35479 24636 35488
rect 24584 35445 24593 35479
rect 24593 35445 24627 35479
rect 24627 35445 24636 35479
rect 24584 35436 24636 35445
rect 25872 35436 25924 35488
rect 26056 35436 26108 35488
rect 28172 35436 28224 35488
rect 28540 35436 28592 35488
rect 33508 35572 33560 35624
rect 33416 35504 33468 35556
rect 30380 35436 30432 35488
rect 30840 35436 30892 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 25136 35232 25188 35284
rect 26240 35232 26292 35284
rect 26332 35232 26384 35284
rect 27252 35232 27304 35284
rect 28080 35275 28132 35284
rect 28080 35241 28089 35275
rect 28089 35241 28123 35275
rect 28123 35241 28132 35275
rect 28080 35232 28132 35241
rect 30656 35232 30708 35284
rect 33508 35275 33560 35284
rect 33508 35241 33517 35275
rect 33517 35241 33551 35275
rect 33551 35241 33560 35275
rect 33508 35232 33560 35241
rect 25964 35096 26016 35148
rect 26148 35096 26200 35148
rect 20260 35028 20312 35080
rect 20536 35071 20588 35080
rect 20536 35037 20545 35071
rect 20545 35037 20579 35071
rect 20579 35037 20588 35071
rect 20536 35028 20588 35037
rect 24584 35028 24636 35080
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 25412 35071 25464 35080
rect 25412 35037 25421 35071
rect 25421 35037 25455 35071
rect 25455 35037 25464 35071
rect 25412 35028 25464 35037
rect 25780 35028 25832 35080
rect 25136 34960 25188 35012
rect 31116 35096 31168 35148
rect 28172 35028 28224 35080
rect 28264 35028 28316 35080
rect 34612 35028 34664 35080
rect 48136 35071 48188 35080
rect 48136 35037 48145 35071
rect 48145 35037 48179 35071
rect 48179 35037 48188 35071
rect 48136 35028 48188 35037
rect 27620 34960 27672 35012
rect 20812 34892 20864 34944
rect 27344 34892 27396 34944
rect 31760 34892 31812 34944
rect 47124 34892 47176 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 25688 34688 25740 34740
rect 29000 34731 29052 34740
rect 29000 34697 29009 34731
rect 29009 34697 29043 34731
rect 29043 34697 29052 34731
rect 29000 34688 29052 34697
rect 29276 34731 29328 34740
rect 29276 34697 29285 34731
rect 29285 34697 29319 34731
rect 29319 34697 29328 34731
rect 29276 34688 29328 34697
rect 29460 34731 29512 34740
rect 29460 34697 29469 34731
rect 29469 34697 29503 34731
rect 29503 34697 29512 34731
rect 29460 34688 29512 34697
rect 31116 34731 31168 34740
rect 31116 34697 31125 34731
rect 31125 34697 31159 34731
rect 31159 34697 31168 34731
rect 31116 34688 31168 34697
rect 20812 34552 20864 34604
rect 22008 34552 22060 34604
rect 24860 34552 24912 34604
rect 29552 34552 29604 34604
rect 29920 34595 29972 34604
rect 29920 34561 29929 34595
rect 29929 34561 29963 34595
rect 29963 34561 29972 34595
rect 29920 34552 29972 34561
rect 22192 34527 22244 34536
rect 22192 34493 22201 34527
rect 22201 34493 22235 34527
rect 22235 34493 22244 34527
rect 22192 34484 22244 34493
rect 23480 34527 23532 34536
rect 23480 34493 23489 34527
rect 23489 34493 23523 34527
rect 23523 34493 23532 34527
rect 23480 34484 23532 34493
rect 23756 34527 23808 34536
rect 23756 34493 23765 34527
rect 23765 34493 23799 34527
rect 23799 34493 23808 34527
rect 23756 34484 23808 34493
rect 25228 34527 25280 34536
rect 25228 34493 25237 34527
rect 25237 34493 25271 34527
rect 25271 34493 25280 34527
rect 25228 34484 25280 34493
rect 25412 34484 25464 34536
rect 25780 34527 25832 34536
rect 25780 34493 25789 34527
rect 25789 34493 25823 34527
rect 25823 34493 25832 34527
rect 25780 34484 25832 34493
rect 27620 34484 27672 34536
rect 28080 34484 28132 34536
rect 31300 34620 31352 34672
rect 33324 34663 33376 34672
rect 33324 34629 33333 34663
rect 33333 34629 33367 34663
rect 33367 34629 33376 34663
rect 33324 34620 33376 34629
rect 34796 34620 34848 34672
rect 48136 34595 48188 34604
rect 48136 34561 48145 34595
rect 48145 34561 48179 34595
rect 48179 34561 48188 34595
rect 48136 34552 48188 34561
rect 31668 34484 31720 34536
rect 34612 34484 34664 34536
rect 23480 34348 23532 34400
rect 24400 34348 24452 34400
rect 27160 34416 27212 34468
rect 25964 34391 26016 34400
rect 25964 34357 25973 34391
rect 25973 34357 26007 34391
rect 26007 34357 26016 34391
rect 25964 34348 26016 34357
rect 26148 34391 26200 34400
rect 26148 34357 26157 34391
rect 26157 34357 26191 34391
rect 26191 34357 26200 34391
rect 26148 34348 26200 34357
rect 27252 34348 27304 34400
rect 47860 34348 47912 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 24860 34144 24912 34196
rect 26056 34187 26108 34196
rect 26056 34153 26065 34187
rect 26065 34153 26099 34187
rect 26099 34153 26108 34187
rect 26056 34144 26108 34153
rect 29552 34144 29604 34196
rect 25596 34076 25648 34128
rect 28632 34076 28684 34128
rect 30932 34144 30984 34196
rect 34796 34187 34848 34196
rect 34796 34153 34805 34187
rect 34805 34153 34839 34187
rect 34839 34153 34848 34187
rect 34796 34144 34848 34153
rect 20076 34008 20128 34060
rect 23480 34008 23532 34060
rect 25780 34008 25832 34060
rect 29092 34008 29144 34060
rect 30380 34008 30432 34060
rect 31484 34008 31536 34060
rect 20812 33940 20864 33992
rect 24584 33983 24636 33992
rect 24584 33949 24593 33983
rect 24593 33949 24627 33983
rect 24627 33949 24636 33983
rect 24584 33940 24636 33949
rect 25320 33940 25372 33992
rect 25872 33983 25924 33992
rect 25872 33949 25881 33983
rect 25881 33949 25915 33983
rect 25915 33949 25924 33983
rect 25872 33940 25924 33949
rect 28172 33983 28224 33992
rect 28172 33949 28181 33983
rect 28181 33949 28215 33983
rect 28215 33949 28224 33983
rect 28172 33940 28224 33949
rect 28816 33940 28868 33992
rect 21640 33915 21692 33924
rect 21640 33881 21649 33915
rect 21649 33881 21683 33915
rect 21683 33881 21692 33915
rect 21640 33872 21692 33881
rect 22192 33872 22244 33924
rect 24768 33872 24820 33924
rect 30380 33872 30432 33924
rect 20536 33804 20588 33856
rect 23572 33804 23624 33856
rect 24676 33804 24728 33856
rect 35348 33940 35400 33992
rect 47952 33940 48004 33992
rect 30748 33915 30800 33924
rect 30748 33881 30757 33915
rect 30757 33881 30791 33915
rect 30791 33881 30800 33915
rect 30748 33872 30800 33881
rect 31760 33872 31812 33924
rect 30840 33804 30892 33856
rect 30932 33804 30984 33856
rect 32680 33872 32732 33924
rect 32220 33847 32272 33856
rect 32220 33813 32229 33847
rect 32229 33813 32263 33847
rect 32263 33813 32272 33847
rect 32220 33804 32272 33813
rect 48044 33847 48096 33856
rect 48044 33813 48053 33847
rect 48053 33813 48087 33847
rect 48087 33813 48096 33847
rect 48044 33804 48096 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 21640 33600 21692 33652
rect 23756 33600 23808 33652
rect 28448 33643 28500 33652
rect 28448 33609 28457 33643
rect 28457 33609 28491 33643
rect 28491 33609 28500 33643
rect 28448 33600 28500 33609
rect 29460 33600 29512 33652
rect 15844 33575 15896 33584
rect 15844 33541 15853 33575
rect 15853 33541 15887 33575
rect 15887 33541 15896 33575
rect 15844 33532 15896 33541
rect 1400 33464 1452 33516
rect 20076 33532 20128 33584
rect 20536 33532 20588 33584
rect 22192 33532 22244 33584
rect 21916 33464 21968 33516
rect 23572 33532 23624 33584
rect 26148 33532 26200 33584
rect 22376 33507 22428 33516
rect 22376 33473 22385 33507
rect 22385 33473 22419 33507
rect 22419 33473 22428 33507
rect 22376 33464 22428 33473
rect 22836 33464 22888 33516
rect 24768 33507 24820 33516
rect 24768 33473 24777 33507
rect 24777 33473 24811 33507
rect 24811 33473 24820 33507
rect 24768 33464 24820 33473
rect 25688 33464 25740 33516
rect 28724 33532 28776 33584
rect 32680 33600 32732 33652
rect 48044 33600 48096 33652
rect 30104 33532 30156 33584
rect 46112 33532 46164 33584
rect 27712 33507 27764 33516
rect 27712 33473 27721 33507
rect 27721 33473 27755 33507
rect 27755 33473 27764 33507
rect 27712 33464 27764 33473
rect 3700 33396 3752 33448
rect 4620 33396 4672 33448
rect 13360 33396 13412 33448
rect 14188 33439 14240 33448
rect 14188 33405 14197 33439
rect 14197 33405 14231 33439
rect 14231 33405 14240 33439
rect 14188 33396 14240 33405
rect 20996 33396 21048 33448
rect 24124 33396 24176 33448
rect 25228 33396 25280 33448
rect 28264 33507 28316 33516
rect 28264 33473 28273 33507
rect 28273 33473 28307 33507
rect 28307 33473 28316 33507
rect 28264 33464 28316 33473
rect 29092 33464 29144 33516
rect 30380 33507 30432 33516
rect 27988 33439 28040 33448
rect 16948 33260 17000 33312
rect 22376 33328 22428 33380
rect 25412 33328 25464 33380
rect 27988 33405 27997 33439
rect 27997 33405 28031 33439
rect 28031 33405 28040 33439
rect 27988 33396 28040 33405
rect 28356 33396 28408 33448
rect 30380 33473 30389 33507
rect 30389 33473 30423 33507
rect 30423 33473 30432 33507
rect 30380 33464 30432 33473
rect 30840 33464 30892 33516
rect 30932 33464 30984 33516
rect 32220 33464 32272 33516
rect 32496 33464 32548 33516
rect 35348 33507 35400 33516
rect 35348 33473 35357 33507
rect 35357 33473 35391 33507
rect 35391 33473 35400 33507
rect 35348 33464 35400 33473
rect 21088 33260 21140 33312
rect 22192 33260 22244 33312
rect 22928 33260 22980 33312
rect 25044 33260 25096 33312
rect 28448 33328 28500 33380
rect 33048 33328 33100 33380
rect 30840 33260 30892 33312
rect 33140 33303 33192 33312
rect 33140 33269 33149 33303
rect 33149 33269 33183 33303
rect 33183 33269 33192 33303
rect 33140 33260 33192 33269
rect 33324 33260 33376 33312
rect 35992 33260 36044 33312
rect 47216 33260 47268 33312
rect 47860 33303 47912 33312
rect 47860 33269 47869 33303
rect 47869 33269 47903 33303
rect 47903 33269 47912 33303
rect 47860 33260 47912 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1676 33056 1728 33108
rect 3700 33056 3752 33108
rect 20996 33056 21048 33108
rect 25044 33099 25096 33108
rect 25044 33065 25053 33099
rect 25053 33065 25087 33099
rect 25087 33065 25096 33099
rect 25044 33056 25096 33065
rect 26240 33056 26292 33108
rect 27712 33056 27764 33108
rect 28816 33099 28868 33108
rect 28816 33065 28825 33099
rect 28825 33065 28859 33099
rect 28859 33065 28868 33099
rect 28816 33056 28868 33065
rect 1400 32963 1452 32972
rect 1400 32929 1409 32963
rect 1409 32929 1443 32963
rect 1443 32929 1452 32963
rect 1400 32920 1452 32929
rect 2780 32852 2832 32904
rect 13268 32920 13320 32972
rect 15936 32963 15988 32972
rect 15936 32929 15945 32963
rect 15945 32929 15979 32963
rect 15979 32929 15988 32963
rect 15936 32920 15988 32929
rect 21548 32920 21600 32972
rect 22008 32920 22060 32972
rect 25964 32988 26016 33040
rect 24584 32920 24636 32972
rect 25596 32920 25648 32972
rect 27988 32988 28040 33040
rect 28264 32988 28316 33040
rect 30656 33056 30708 33108
rect 30748 33056 30800 33108
rect 32312 33056 32364 33108
rect 32496 33099 32548 33108
rect 32496 33065 32505 33099
rect 32505 33065 32539 33099
rect 32539 33065 32548 33099
rect 32496 33056 32548 33065
rect 30380 32988 30432 33040
rect 32864 33031 32916 33040
rect 32864 32997 32873 33031
rect 32873 32997 32907 33031
rect 32907 32997 32916 33031
rect 32864 32988 32916 32997
rect 47032 32988 47084 33040
rect 9588 32852 9640 32904
rect 14004 32852 14056 32904
rect 21088 32895 21140 32904
rect 21088 32861 21097 32895
rect 21097 32861 21131 32895
rect 21131 32861 21140 32895
rect 21088 32852 21140 32861
rect 21272 32852 21324 32904
rect 22376 32852 22428 32904
rect 22560 32852 22612 32904
rect 24768 32852 24820 32904
rect 22744 32716 22796 32768
rect 25228 32852 25280 32904
rect 29552 32920 29604 32972
rect 25688 32827 25740 32836
rect 25688 32793 25697 32827
rect 25697 32793 25731 32827
rect 25731 32793 25740 32827
rect 25688 32784 25740 32793
rect 25780 32784 25832 32836
rect 28540 32852 28592 32904
rect 28724 32852 28776 32904
rect 29092 32895 29144 32904
rect 29092 32861 29101 32895
rect 29101 32861 29135 32895
rect 29135 32861 29144 32895
rect 29092 32852 29144 32861
rect 29920 32852 29972 32904
rect 30932 32920 30984 32972
rect 33140 32920 33192 32972
rect 30656 32895 30708 32904
rect 30656 32861 30665 32895
rect 30665 32861 30699 32895
rect 30699 32861 30708 32895
rect 30656 32852 30708 32861
rect 30840 32895 30892 32904
rect 30840 32861 30849 32895
rect 30849 32861 30883 32895
rect 30883 32861 30892 32895
rect 32496 32895 32548 32904
rect 30840 32852 30892 32861
rect 29552 32716 29604 32768
rect 32496 32861 32505 32895
rect 32505 32861 32539 32895
rect 32539 32861 32548 32895
rect 32496 32852 32548 32861
rect 33048 32852 33100 32904
rect 34980 32920 35032 32972
rect 47124 32963 47176 32972
rect 47124 32929 47133 32963
rect 47133 32929 47167 32963
rect 47167 32929 47176 32963
rect 47124 32920 47176 32929
rect 33508 32852 33560 32904
rect 46296 32852 46348 32904
rect 33784 32827 33836 32836
rect 33784 32793 33793 32827
rect 33793 32793 33827 32827
rect 33827 32793 33836 32827
rect 33784 32784 33836 32793
rect 30564 32716 30616 32768
rect 30748 32716 30800 32768
rect 32956 32716 33008 32768
rect 33048 32716 33100 32768
rect 34428 32716 34480 32768
rect 35072 32784 35124 32836
rect 35992 32784 36044 32836
rect 47216 32827 47268 32836
rect 47216 32793 47225 32827
rect 47225 32793 47259 32827
rect 47259 32793 47268 32827
rect 47216 32784 47268 32793
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 3148 32512 3200 32564
rect 41144 32512 41196 32564
rect 2780 32487 2832 32496
rect 2780 32453 2789 32487
rect 2789 32453 2823 32487
rect 2823 32453 2832 32487
rect 2780 32444 2832 32453
rect 8300 32444 8352 32496
rect 2596 32351 2648 32360
rect 2596 32317 2605 32351
rect 2605 32317 2639 32351
rect 2639 32317 2648 32351
rect 2596 32308 2648 32317
rect 4620 32308 4672 32360
rect 2044 32172 2096 32224
rect 9772 32308 9824 32360
rect 12532 32444 12584 32496
rect 14188 32444 14240 32496
rect 20352 32444 20404 32496
rect 21272 32487 21324 32496
rect 21272 32453 21281 32487
rect 21281 32453 21315 32487
rect 21315 32453 21324 32487
rect 21272 32444 21324 32453
rect 21456 32444 21508 32496
rect 22100 32444 22152 32496
rect 25044 32444 25096 32496
rect 25504 32444 25556 32496
rect 25964 32444 26016 32496
rect 27160 32487 27212 32496
rect 27160 32453 27169 32487
rect 27169 32453 27203 32487
rect 27203 32453 27212 32487
rect 27160 32444 27212 32453
rect 14004 32419 14056 32428
rect 14004 32385 14013 32419
rect 14013 32385 14047 32419
rect 14047 32385 14056 32419
rect 14004 32376 14056 32385
rect 21732 32376 21784 32428
rect 21916 32376 21968 32428
rect 24768 32376 24820 32428
rect 25596 32376 25648 32428
rect 29644 32444 29696 32496
rect 29920 32487 29972 32496
rect 29920 32453 29929 32487
rect 29929 32453 29963 32487
rect 29963 32453 29972 32487
rect 29920 32444 29972 32453
rect 10784 32308 10836 32360
rect 11796 32351 11848 32360
rect 11796 32317 11805 32351
rect 11805 32317 11839 32351
rect 11839 32317 11848 32351
rect 11796 32308 11848 32317
rect 13268 32351 13320 32360
rect 13268 32317 13277 32351
rect 13277 32317 13311 32351
rect 13311 32317 13320 32351
rect 13268 32308 13320 32317
rect 13544 32308 13596 32360
rect 27988 32376 28040 32428
rect 28632 32376 28684 32428
rect 29092 32376 29144 32428
rect 30104 32419 30156 32428
rect 30104 32385 30113 32419
rect 30113 32385 30147 32419
rect 30147 32385 30156 32419
rect 30104 32376 30156 32385
rect 30932 32444 30984 32496
rect 32864 32444 32916 32496
rect 27896 32308 27948 32360
rect 28080 32308 28132 32360
rect 28816 32308 28868 32360
rect 30472 32419 30524 32428
rect 30472 32385 30481 32419
rect 30481 32385 30515 32419
rect 30515 32385 30524 32419
rect 30472 32376 30524 32385
rect 32312 32419 32364 32428
rect 32312 32385 32321 32419
rect 32321 32385 32355 32419
rect 32355 32385 32364 32419
rect 32312 32376 32364 32385
rect 33324 32419 33376 32428
rect 33324 32385 33333 32419
rect 33333 32385 33367 32419
rect 33367 32385 33376 32419
rect 33324 32376 33376 32385
rect 35072 32444 35124 32496
rect 34428 32419 34480 32428
rect 34428 32385 34437 32419
rect 34437 32385 34471 32419
rect 34471 32385 34480 32419
rect 34428 32376 34480 32385
rect 34520 32376 34572 32428
rect 34980 32419 35032 32428
rect 34980 32385 34989 32419
rect 34989 32385 35023 32419
rect 35023 32385 35032 32419
rect 34980 32376 35032 32385
rect 35440 32376 35492 32428
rect 30564 32308 30616 32360
rect 32496 32308 32548 32360
rect 47492 32376 47544 32428
rect 46204 32351 46256 32360
rect 46204 32317 46213 32351
rect 46213 32317 46247 32351
rect 46247 32317 46256 32351
rect 46204 32308 46256 32317
rect 22284 32240 22336 32292
rect 25964 32240 26016 32292
rect 12992 32172 13044 32224
rect 14556 32172 14608 32224
rect 22560 32172 22612 32224
rect 23388 32172 23440 32224
rect 26792 32172 26844 32224
rect 34520 32240 34572 32292
rect 30748 32172 30800 32224
rect 31208 32215 31260 32224
rect 31208 32181 31217 32215
rect 31217 32181 31251 32215
rect 31251 32181 31260 32215
rect 31208 32172 31260 32181
rect 31300 32172 31352 32224
rect 46480 32172 46532 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1676 31968 1728 32020
rect 9772 32011 9824 32020
rect 9772 31977 9781 32011
rect 9781 31977 9815 32011
rect 9815 31977 9824 32011
rect 9772 31968 9824 31977
rect 10784 32011 10836 32020
rect 10784 31977 10793 32011
rect 10793 31977 10827 32011
rect 10827 31977 10836 32011
rect 10784 31968 10836 31977
rect 11796 32011 11848 32020
rect 11796 31977 11805 32011
rect 11805 31977 11839 32011
rect 11839 31977 11848 32011
rect 11796 31968 11848 31977
rect 12532 31968 12584 32020
rect 15108 32011 15160 32020
rect 15108 31977 15117 32011
rect 15117 31977 15151 32011
rect 15151 31977 15160 32011
rect 15108 31968 15160 31977
rect 21088 31968 21140 32020
rect 22560 31968 22612 32020
rect 22744 32011 22796 32020
rect 22744 31977 22753 32011
rect 22753 31977 22787 32011
rect 22787 31977 22796 32011
rect 22744 31968 22796 31977
rect 22928 32011 22980 32020
rect 22928 31977 22937 32011
rect 22937 31977 22971 32011
rect 22971 31977 22980 32011
rect 22928 31968 22980 31977
rect 24584 31968 24636 32020
rect 25964 31968 26016 32020
rect 26148 31968 26200 32020
rect 27160 31968 27212 32020
rect 28264 31968 28316 32020
rect 29092 31968 29144 32020
rect 11704 31900 11756 31952
rect 14556 31875 14608 31884
rect 14556 31841 14565 31875
rect 14565 31841 14599 31875
rect 14599 31841 14608 31875
rect 14556 31832 14608 31841
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 3148 31764 3200 31816
rect 9588 31764 9640 31816
rect 10692 31807 10744 31816
rect 10692 31773 10701 31807
rect 10701 31773 10735 31807
rect 10735 31773 10744 31807
rect 10692 31764 10744 31773
rect 12440 31764 12492 31816
rect 13176 31807 13228 31816
rect 12256 31696 12308 31748
rect 13176 31773 13185 31807
rect 13185 31773 13219 31807
rect 13219 31773 13228 31807
rect 13176 31764 13228 31773
rect 13360 31807 13412 31816
rect 13360 31773 13369 31807
rect 13369 31773 13403 31807
rect 13403 31773 13412 31807
rect 13360 31764 13412 31773
rect 14280 31807 14332 31816
rect 14280 31773 14289 31807
rect 14289 31773 14323 31807
rect 14323 31773 14332 31807
rect 14280 31764 14332 31773
rect 14464 31807 14516 31816
rect 14464 31773 14473 31807
rect 14473 31773 14507 31807
rect 14507 31773 14516 31807
rect 14464 31764 14516 31773
rect 20812 31832 20864 31884
rect 20168 31764 20220 31816
rect 21456 31832 21508 31884
rect 22100 31832 22152 31884
rect 21364 31807 21416 31816
rect 21364 31773 21373 31807
rect 21373 31773 21407 31807
rect 21407 31773 21416 31807
rect 22560 31832 22612 31884
rect 25044 31900 25096 31952
rect 25872 31900 25924 31952
rect 31576 31968 31628 32020
rect 29276 31900 29328 31952
rect 31208 31900 31260 31952
rect 31300 31900 31352 31952
rect 32680 31900 32732 31952
rect 33232 31900 33284 31952
rect 21364 31764 21416 31773
rect 22744 31807 22796 31816
rect 22744 31773 22753 31807
rect 22753 31773 22787 31807
rect 22787 31773 22796 31807
rect 22744 31764 22796 31773
rect 16856 31696 16908 31748
rect 25044 31764 25096 31816
rect 25412 31764 25464 31816
rect 25688 31807 25740 31816
rect 25688 31773 25697 31807
rect 25697 31773 25731 31807
rect 25731 31773 25740 31807
rect 25688 31764 25740 31773
rect 25780 31764 25832 31816
rect 26056 31807 26108 31816
rect 26056 31773 26065 31807
rect 26065 31773 26099 31807
rect 26099 31773 26108 31807
rect 26056 31764 26108 31773
rect 2964 31671 3016 31680
rect 2964 31637 2973 31671
rect 2973 31637 3007 31671
rect 3007 31637 3016 31671
rect 2964 31628 3016 31637
rect 12440 31628 12492 31680
rect 13544 31628 13596 31680
rect 14096 31671 14148 31680
rect 14096 31637 14105 31671
rect 14105 31637 14139 31671
rect 14139 31637 14148 31671
rect 14096 31628 14148 31637
rect 21640 31671 21692 31680
rect 21640 31637 21649 31671
rect 21649 31637 21683 31671
rect 21683 31637 21692 31671
rect 21640 31628 21692 31637
rect 24492 31671 24544 31680
rect 24492 31637 24501 31671
rect 24501 31637 24535 31671
rect 24535 31637 24544 31671
rect 24492 31628 24544 31637
rect 26056 31628 26108 31680
rect 27896 31832 27948 31884
rect 28264 31832 28316 31884
rect 28448 31832 28500 31884
rect 30472 31832 30524 31884
rect 26792 31807 26844 31816
rect 26792 31773 26801 31807
rect 26801 31773 26835 31807
rect 26835 31773 26844 31807
rect 26792 31764 26844 31773
rect 27804 31764 27856 31816
rect 27528 31739 27580 31748
rect 27528 31705 27537 31739
rect 27537 31705 27571 31739
rect 27571 31705 27580 31739
rect 27528 31696 27580 31705
rect 31576 31764 31628 31816
rect 32312 31807 32364 31816
rect 32312 31773 32319 31807
rect 32319 31773 32364 31807
rect 32312 31764 32364 31773
rect 32496 31807 32548 31816
rect 32496 31773 32505 31807
rect 32505 31773 32539 31807
rect 32539 31773 32548 31807
rect 32496 31764 32548 31773
rect 32680 31764 32732 31816
rect 35348 31832 35400 31884
rect 46296 31875 46348 31884
rect 46296 31841 46305 31875
rect 46305 31841 46339 31875
rect 46339 31841 46348 31875
rect 46296 31832 46348 31841
rect 46480 31875 46532 31884
rect 46480 31841 46489 31875
rect 46489 31841 46523 31875
rect 46523 31841 46532 31875
rect 46480 31832 46532 31841
rect 48136 31875 48188 31884
rect 48136 31841 48145 31875
rect 48145 31841 48179 31875
rect 48179 31841 48188 31875
rect 48136 31832 48188 31841
rect 34796 31807 34848 31816
rect 34796 31773 34805 31807
rect 34805 31773 34839 31807
rect 34839 31773 34848 31807
rect 34796 31764 34848 31773
rect 33784 31628 33836 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 14648 31424 14700 31476
rect 20904 31424 20956 31476
rect 21456 31424 21508 31476
rect 21732 31424 21784 31476
rect 27160 31424 27212 31476
rect 27528 31424 27580 31476
rect 31208 31424 31260 31476
rect 31576 31424 31628 31476
rect 32312 31424 32364 31476
rect 2964 31356 3016 31408
rect 14096 31356 14148 31408
rect 20168 31356 20220 31408
rect 23480 31356 23532 31408
rect 2044 31331 2096 31340
rect 2044 31297 2053 31331
rect 2053 31297 2087 31331
rect 2087 31297 2096 31331
rect 2044 31288 2096 31297
rect 10692 31288 10744 31340
rect 10876 31331 10928 31340
rect 10876 31297 10885 31331
rect 10885 31297 10919 31331
rect 10919 31297 10928 31331
rect 10876 31288 10928 31297
rect 12256 31331 12308 31340
rect 12256 31297 12265 31331
rect 12265 31297 12299 31331
rect 12299 31297 12308 31331
rect 12256 31288 12308 31297
rect 15108 31288 15160 31340
rect 15292 31288 15344 31340
rect 16856 31288 16908 31340
rect 20812 31288 20864 31340
rect 21272 31288 21324 31340
rect 22284 31288 22336 31340
rect 22928 31288 22980 31340
rect 24676 31356 24728 31408
rect 2780 31263 2832 31272
rect 2780 31229 2789 31263
rect 2789 31229 2823 31263
rect 2823 31229 2832 31263
rect 2780 31220 2832 31229
rect 18880 31263 18932 31272
rect 18880 31229 18889 31263
rect 18889 31229 18923 31263
rect 18923 31229 18932 31263
rect 18880 31220 18932 31229
rect 20628 31220 20680 31272
rect 22468 31220 22520 31272
rect 26332 31288 26384 31340
rect 31576 31288 31628 31340
rect 33508 31356 33560 31408
rect 34796 31356 34848 31408
rect 46112 31399 46164 31408
rect 46112 31365 46121 31399
rect 46121 31365 46155 31399
rect 46155 31365 46164 31399
rect 46112 31356 46164 31365
rect 24492 31220 24544 31272
rect 33232 31263 33284 31272
rect 33232 31229 33241 31263
rect 33241 31229 33275 31263
rect 33275 31229 33284 31263
rect 33232 31220 33284 31229
rect 46020 31263 46072 31272
rect 46020 31229 46029 31263
rect 46029 31229 46063 31263
rect 46063 31229 46072 31263
rect 46020 31220 46072 31229
rect 47032 31220 47084 31272
rect 22284 31152 22336 31204
rect 22744 31152 22796 31204
rect 10784 31084 10836 31136
rect 12348 31127 12400 31136
rect 12348 31093 12357 31127
rect 12357 31093 12391 31127
rect 12391 31093 12400 31127
rect 12348 31084 12400 31093
rect 16672 31084 16724 31136
rect 21180 31127 21232 31136
rect 21180 31093 21189 31127
rect 21189 31093 21223 31127
rect 21223 31093 21232 31127
rect 21180 31084 21232 31093
rect 21732 31084 21784 31136
rect 24952 31084 25004 31136
rect 26056 31084 26108 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 21364 30880 21416 30932
rect 25688 30923 25740 30932
rect 25688 30889 25697 30923
rect 25697 30889 25731 30923
rect 25731 30889 25740 30923
rect 25688 30880 25740 30889
rect 26332 30923 26384 30932
rect 26332 30889 26341 30923
rect 26341 30889 26375 30923
rect 26375 30889 26384 30923
rect 26332 30880 26384 30889
rect 26792 30880 26844 30932
rect 29000 30880 29052 30932
rect 29644 30880 29696 30932
rect 12992 30855 13044 30864
rect 12992 30821 13001 30855
rect 13001 30821 13035 30855
rect 13035 30821 13044 30855
rect 12992 30812 13044 30821
rect 21548 30812 21600 30864
rect 10784 30787 10836 30796
rect 10784 30753 10793 30787
rect 10793 30753 10827 30787
rect 10827 30753 10836 30787
rect 10784 30744 10836 30753
rect 14280 30744 14332 30796
rect 13544 30676 13596 30728
rect 14372 30676 14424 30728
rect 18880 30744 18932 30796
rect 20076 30744 20128 30796
rect 26148 30744 26200 30796
rect 28540 30744 28592 30796
rect 15660 30719 15712 30728
rect 15660 30685 15669 30719
rect 15669 30685 15703 30719
rect 15703 30685 15712 30719
rect 15660 30676 15712 30685
rect 21180 30676 21232 30728
rect 22284 30719 22336 30728
rect 11060 30651 11112 30660
rect 11060 30617 11069 30651
rect 11069 30617 11103 30651
rect 11103 30617 11112 30651
rect 11060 30608 11112 30617
rect 12348 30608 12400 30660
rect 13360 30651 13412 30660
rect 13360 30617 13369 30651
rect 13369 30617 13403 30651
rect 13403 30617 13412 30651
rect 13360 30608 13412 30617
rect 12624 30540 12676 30592
rect 14188 30540 14240 30592
rect 16672 30608 16724 30660
rect 21364 30608 21416 30660
rect 22284 30685 22293 30719
rect 22293 30685 22327 30719
rect 22327 30685 22336 30719
rect 22284 30676 22336 30685
rect 22376 30676 22428 30728
rect 23388 30719 23440 30728
rect 23388 30685 23397 30719
rect 23397 30685 23431 30719
rect 23431 30685 23440 30719
rect 23388 30676 23440 30685
rect 26056 30676 26108 30728
rect 26240 30719 26292 30728
rect 26240 30685 26249 30719
rect 26249 30685 26283 30719
rect 26283 30685 26292 30719
rect 26240 30676 26292 30685
rect 28724 30676 28776 30728
rect 31392 30744 31444 30796
rect 35808 30812 35860 30864
rect 30472 30676 30524 30728
rect 31024 30676 31076 30728
rect 31300 30676 31352 30728
rect 34520 30744 34572 30796
rect 33784 30719 33836 30728
rect 33784 30685 33793 30719
rect 33793 30685 33827 30719
rect 33827 30685 33836 30719
rect 33784 30676 33836 30685
rect 44364 30744 44416 30796
rect 35164 30719 35216 30728
rect 35164 30685 35173 30719
rect 35173 30685 35207 30719
rect 35207 30685 35216 30719
rect 35440 30719 35492 30728
rect 35164 30676 35216 30685
rect 35440 30685 35449 30719
rect 35449 30685 35483 30719
rect 35483 30685 35492 30719
rect 35440 30676 35492 30685
rect 22560 30608 22612 30660
rect 24860 30608 24912 30660
rect 28632 30608 28684 30660
rect 31116 30608 31168 30660
rect 32312 30608 32364 30660
rect 21916 30540 21968 30592
rect 24676 30583 24728 30592
rect 24676 30549 24685 30583
rect 24685 30549 24719 30583
rect 24719 30549 24728 30583
rect 24676 30540 24728 30549
rect 30656 30583 30708 30592
rect 30656 30549 30665 30583
rect 30665 30549 30699 30583
rect 30699 30549 30708 30583
rect 30656 30540 30708 30549
rect 31576 30583 31628 30592
rect 31576 30549 31585 30583
rect 31585 30549 31619 30583
rect 31619 30549 31628 30583
rect 31576 30540 31628 30549
rect 32220 30583 32272 30592
rect 32220 30549 32229 30583
rect 32229 30549 32263 30583
rect 32263 30549 32272 30583
rect 32220 30540 32272 30549
rect 34520 30608 34572 30660
rect 34152 30540 34204 30592
rect 35256 30540 35308 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 11060 30336 11112 30388
rect 12624 30336 12676 30388
rect 14280 30379 14332 30388
rect 14280 30345 14289 30379
rect 14289 30345 14323 30379
rect 14323 30345 14332 30379
rect 14280 30336 14332 30345
rect 15660 30336 15712 30388
rect 21456 30336 21508 30388
rect 22376 30336 22428 30388
rect 12716 30268 12768 30320
rect 13360 30268 13412 30320
rect 20628 30268 20680 30320
rect 21824 30268 21876 30320
rect 10600 30243 10652 30252
rect 10600 30209 10609 30243
rect 10609 30209 10643 30243
rect 10643 30209 10652 30243
rect 10600 30200 10652 30209
rect 10692 30243 10744 30252
rect 10692 30209 10701 30243
rect 10701 30209 10735 30243
rect 10735 30209 10744 30243
rect 10968 30243 11020 30252
rect 10692 30200 10744 30209
rect 10968 30209 10977 30243
rect 10977 30209 11011 30243
rect 11011 30209 11020 30243
rect 10968 30200 11020 30209
rect 12440 30243 12492 30252
rect 12440 30209 12449 30243
rect 12449 30209 12483 30243
rect 12483 30209 12492 30243
rect 12440 30200 12492 30209
rect 13176 30200 13228 30252
rect 14188 30200 14240 30252
rect 15292 30200 15344 30252
rect 20904 30243 20956 30252
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 21732 30200 21784 30252
rect 21916 30243 21968 30252
rect 21916 30209 21925 30243
rect 21925 30209 21959 30243
rect 21959 30209 21968 30243
rect 21916 30200 21968 30209
rect 23020 30268 23072 30320
rect 22376 30200 22428 30252
rect 22652 30200 22704 30252
rect 14464 30132 14516 30184
rect 20536 30175 20588 30184
rect 20536 30141 20545 30175
rect 20545 30141 20579 30175
rect 20579 30141 20588 30175
rect 20536 30132 20588 30141
rect 22284 30175 22336 30184
rect 22284 30141 22293 30175
rect 22293 30141 22327 30175
rect 22327 30141 22336 30175
rect 22284 30132 22336 30141
rect 17132 30064 17184 30116
rect 12440 29996 12492 30048
rect 21364 30064 21416 30116
rect 24216 30243 24268 30252
rect 25688 30268 25740 30320
rect 25964 30268 26016 30320
rect 27712 30268 27764 30320
rect 28172 30268 28224 30320
rect 31576 30336 31628 30388
rect 35164 30336 35216 30388
rect 24216 30209 24258 30243
rect 24258 30209 24268 30243
rect 24216 30200 24268 30209
rect 25412 30243 25464 30252
rect 25412 30209 25421 30243
rect 25421 30209 25455 30243
rect 25455 30209 25464 30243
rect 25412 30200 25464 30209
rect 26056 30243 26108 30252
rect 26056 30209 26065 30243
rect 26065 30209 26099 30243
rect 26099 30209 26108 30243
rect 26056 30200 26108 30209
rect 27528 30243 27580 30252
rect 27528 30209 27537 30243
rect 27537 30209 27571 30243
rect 27571 30209 27580 30243
rect 27528 30200 27580 30209
rect 24768 30175 24820 30184
rect 24768 30141 24777 30175
rect 24777 30141 24811 30175
rect 24811 30141 24820 30175
rect 24768 30132 24820 30141
rect 25044 30132 25096 30184
rect 28172 30132 28224 30184
rect 29000 30200 29052 30252
rect 32220 30268 32272 30320
rect 33324 30243 33376 30252
rect 33324 30209 33333 30243
rect 33333 30209 33367 30243
rect 33367 30209 33376 30243
rect 33324 30200 33376 30209
rect 33508 30268 33560 30320
rect 35256 30311 35308 30320
rect 34152 30243 34204 30252
rect 34152 30209 34161 30243
rect 34161 30209 34195 30243
rect 34195 30209 34204 30243
rect 34152 30200 34204 30209
rect 35256 30277 35265 30311
rect 35265 30277 35299 30311
rect 35299 30277 35308 30311
rect 35256 30268 35308 30277
rect 35900 30268 35952 30320
rect 30564 30132 30616 30184
rect 31300 30132 31352 30184
rect 34244 30132 34296 30184
rect 24124 30107 24176 30116
rect 24124 30073 24133 30107
rect 24133 30073 24167 30107
rect 24167 30073 24176 30107
rect 24124 30064 24176 30073
rect 24860 29996 24912 30048
rect 28540 30064 28592 30116
rect 31116 30064 31168 30116
rect 34796 30064 34848 30116
rect 26608 29996 26660 30048
rect 27620 29996 27672 30048
rect 31392 29996 31444 30048
rect 31668 29996 31720 30048
rect 34152 29996 34204 30048
rect 34428 29996 34480 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 9312 29792 9364 29844
rect 17132 29792 17184 29844
rect 20536 29792 20588 29844
rect 21548 29792 21600 29844
rect 24768 29792 24820 29844
rect 24952 29835 25004 29844
rect 24952 29801 24961 29835
rect 24961 29801 24995 29835
rect 24995 29801 25004 29835
rect 24952 29792 25004 29801
rect 29000 29835 29052 29844
rect 10968 29656 11020 29708
rect 23020 29724 23072 29776
rect 29000 29801 29009 29835
rect 29009 29801 29043 29835
rect 29043 29801 29052 29835
rect 29000 29792 29052 29801
rect 30564 29835 30616 29844
rect 30564 29801 30573 29835
rect 30573 29801 30607 29835
rect 30607 29801 30616 29835
rect 30564 29792 30616 29801
rect 30748 29792 30800 29844
rect 29552 29724 29604 29776
rect 15292 29588 15344 29640
rect 9680 29520 9732 29572
rect 9036 29452 9088 29504
rect 15752 29520 15804 29572
rect 16948 29520 17000 29572
rect 22100 29588 22152 29640
rect 24676 29656 24728 29708
rect 28816 29656 28868 29708
rect 25044 29588 25096 29640
rect 25964 29631 26016 29640
rect 25964 29597 25973 29631
rect 25973 29597 26007 29631
rect 26007 29597 26016 29631
rect 25964 29588 26016 29597
rect 26148 29631 26200 29640
rect 26148 29597 26157 29631
rect 26157 29597 26191 29631
rect 26191 29597 26200 29631
rect 26148 29588 26200 29597
rect 29828 29631 29880 29640
rect 24216 29520 24268 29572
rect 24492 29520 24544 29572
rect 26056 29520 26108 29572
rect 29828 29597 29837 29631
rect 29837 29597 29871 29631
rect 29871 29597 29880 29631
rect 29828 29588 29880 29597
rect 30656 29656 30708 29708
rect 30380 29631 30432 29640
rect 27804 29520 27856 29572
rect 29276 29520 29328 29572
rect 29736 29520 29788 29572
rect 30380 29597 30389 29631
rect 30389 29597 30423 29631
rect 30423 29597 30432 29631
rect 30380 29588 30432 29597
rect 30656 29520 30708 29572
rect 17868 29495 17920 29504
rect 17868 29461 17877 29495
rect 17877 29461 17911 29495
rect 17911 29461 17920 29495
rect 17868 29452 17920 29461
rect 21456 29495 21508 29504
rect 21456 29461 21465 29495
rect 21465 29461 21499 29495
rect 21499 29461 21508 29495
rect 21456 29452 21508 29461
rect 24768 29452 24820 29504
rect 26608 29452 26660 29504
rect 34704 29835 34756 29844
rect 34704 29801 34713 29835
rect 34713 29801 34747 29835
rect 34747 29801 34756 29835
rect 34704 29792 34756 29801
rect 34796 29792 34848 29844
rect 35900 29835 35952 29844
rect 35900 29801 35909 29835
rect 35909 29801 35943 29835
rect 35943 29801 35952 29835
rect 35900 29792 35952 29801
rect 31576 29656 31628 29708
rect 31392 29588 31444 29640
rect 33324 29699 33376 29708
rect 33324 29665 33333 29699
rect 33333 29665 33367 29699
rect 33367 29665 33376 29699
rect 34888 29699 34940 29708
rect 33324 29656 33376 29665
rect 34888 29665 34897 29699
rect 34897 29665 34931 29699
rect 34931 29665 34940 29699
rect 34888 29656 34940 29665
rect 47216 29656 47268 29708
rect 32036 29631 32088 29640
rect 32036 29597 32045 29631
rect 32045 29597 32079 29631
rect 32079 29597 32088 29631
rect 32036 29588 32088 29597
rect 32404 29631 32456 29640
rect 32404 29597 32413 29631
rect 32413 29597 32447 29631
rect 32447 29597 32456 29631
rect 32404 29588 32456 29597
rect 33140 29588 33192 29640
rect 33324 29520 33376 29572
rect 34520 29588 34572 29640
rect 34612 29588 34664 29640
rect 35808 29631 35860 29640
rect 35808 29597 35817 29631
rect 35817 29597 35851 29631
rect 35851 29597 35860 29631
rect 35808 29588 35860 29597
rect 47400 29588 47452 29640
rect 34428 29520 34480 29572
rect 34520 29452 34572 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 9680 29291 9732 29300
rect 9680 29257 9689 29291
rect 9689 29257 9723 29291
rect 9723 29257 9732 29291
rect 9680 29248 9732 29257
rect 16948 29291 17000 29300
rect 16948 29257 16957 29291
rect 16957 29257 16991 29291
rect 16991 29257 17000 29291
rect 16948 29248 17000 29257
rect 25412 29248 25464 29300
rect 32312 29291 32364 29300
rect 13176 29180 13228 29232
rect 14464 29180 14516 29232
rect 21640 29180 21692 29232
rect 25596 29180 25648 29232
rect 32312 29257 32321 29291
rect 32321 29257 32355 29291
rect 32355 29257 32364 29291
rect 32312 29248 32364 29257
rect 32404 29248 32456 29300
rect 9588 29155 9640 29164
rect 9588 29121 9597 29155
rect 9597 29121 9631 29155
rect 9631 29121 9640 29155
rect 9588 29112 9640 29121
rect 13544 29112 13596 29164
rect 15200 29112 15252 29164
rect 15660 29112 15712 29164
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 16856 29112 16908 29121
rect 22468 29112 22520 29164
rect 23296 29112 23348 29164
rect 27896 29155 27948 29164
rect 15476 29087 15528 29096
rect 15476 29053 15485 29087
rect 15485 29053 15519 29087
rect 15519 29053 15528 29087
rect 15476 29044 15528 29053
rect 15752 29087 15804 29096
rect 15752 29053 15761 29087
rect 15761 29053 15795 29087
rect 15795 29053 15804 29087
rect 15752 29044 15804 29053
rect 13636 29019 13688 29028
rect 13636 28985 13645 29019
rect 13645 28985 13679 29019
rect 13679 28985 13688 29019
rect 13636 28976 13688 28985
rect 27896 29121 27905 29155
rect 27905 29121 27939 29155
rect 27939 29121 27948 29155
rect 27896 29112 27948 29121
rect 30656 29155 30708 29164
rect 30656 29121 30665 29155
rect 30665 29121 30699 29155
rect 30699 29121 30708 29155
rect 30656 29112 30708 29121
rect 31392 29112 31444 29164
rect 34888 29248 34940 29300
rect 34520 29223 34572 29232
rect 34520 29189 34529 29223
rect 34529 29189 34563 29223
rect 34563 29189 34572 29223
rect 34520 29180 34572 29189
rect 35532 29180 35584 29232
rect 34244 29155 34296 29164
rect 34244 29121 34253 29155
rect 34253 29121 34287 29155
rect 34287 29121 34296 29155
rect 34244 29112 34296 29121
rect 24952 29044 25004 29096
rect 30380 29044 30432 29096
rect 10140 28908 10192 28960
rect 10692 28908 10744 28960
rect 12716 28908 12768 28960
rect 14740 28908 14792 28960
rect 21824 28976 21876 29028
rect 26056 29019 26108 29028
rect 26056 28985 26065 29019
rect 26065 28985 26099 29019
rect 26099 28985 26108 29019
rect 26056 28976 26108 28985
rect 27528 28976 27580 29028
rect 30564 28976 30616 29028
rect 21088 28908 21140 28960
rect 22560 28908 22612 28960
rect 25320 28908 25372 28960
rect 30748 28976 30800 29028
rect 31024 29019 31076 29028
rect 31024 28985 31033 29019
rect 31033 28985 31067 29019
rect 31067 28985 31076 29019
rect 34152 29044 34204 29096
rect 31024 28976 31076 28985
rect 33508 28908 33560 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 14464 28747 14516 28756
rect 14464 28713 14473 28747
rect 14473 28713 14507 28747
rect 14507 28713 14516 28747
rect 14464 28704 14516 28713
rect 10600 28636 10652 28688
rect 10876 28636 10928 28688
rect 14096 28636 14148 28688
rect 12716 28568 12768 28620
rect 14188 28568 14240 28620
rect 10140 28543 10192 28552
rect 10140 28509 10149 28543
rect 10149 28509 10183 28543
rect 10183 28509 10192 28543
rect 10140 28500 10192 28509
rect 10968 28543 11020 28552
rect 10968 28509 10977 28543
rect 10977 28509 11011 28543
rect 11011 28509 11020 28543
rect 10968 28500 11020 28509
rect 11980 28432 12032 28484
rect 14740 28500 14792 28552
rect 15200 28500 15252 28552
rect 16672 28568 16724 28620
rect 21640 28568 21692 28620
rect 26240 28704 26292 28756
rect 27804 28704 27856 28756
rect 28816 28704 28868 28756
rect 29828 28704 29880 28756
rect 30472 28704 30524 28756
rect 31484 28704 31536 28756
rect 33508 28747 33560 28756
rect 33508 28713 33517 28747
rect 33517 28713 33551 28747
rect 33551 28713 33560 28747
rect 33508 28704 33560 28713
rect 33968 28704 34020 28756
rect 35348 28704 35400 28756
rect 35532 28747 35584 28756
rect 35532 28713 35541 28747
rect 35541 28713 35575 28747
rect 35575 28713 35584 28747
rect 35532 28704 35584 28713
rect 22744 28636 22796 28688
rect 22928 28636 22980 28688
rect 15936 28500 15988 28552
rect 17776 28500 17828 28552
rect 14556 28432 14608 28484
rect 15568 28432 15620 28484
rect 16304 28475 16356 28484
rect 16304 28441 16313 28475
rect 16313 28441 16347 28475
rect 16347 28441 16356 28475
rect 16304 28432 16356 28441
rect 17316 28432 17368 28484
rect 20996 28500 21048 28552
rect 21824 28543 21876 28552
rect 21824 28509 21833 28543
rect 21833 28509 21867 28543
rect 21867 28509 21876 28543
rect 21824 28500 21876 28509
rect 22744 28500 22796 28552
rect 24584 28543 24636 28552
rect 19432 28432 19484 28484
rect 20536 28432 20588 28484
rect 21180 28432 21232 28484
rect 21732 28475 21784 28484
rect 21732 28441 21741 28475
rect 21741 28441 21775 28475
rect 21775 28441 21784 28475
rect 21732 28432 21784 28441
rect 22560 28432 22612 28484
rect 24584 28509 24593 28543
rect 24593 28509 24627 28543
rect 24627 28509 24636 28543
rect 24584 28500 24636 28509
rect 26056 28568 26108 28620
rect 24768 28432 24820 28484
rect 14372 28364 14424 28416
rect 18052 28364 18104 28416
rect 18236 28364 18288 28416
rect 21364 28364 21416 28416
rect 22008 28407 22060 28416
rect 22008 28373 22017 28407
rect 22017 28373 22051 28407
rect 22051 28373 22060 28407
rect 22008 28364 22060 28373
rect 22284 28364 22336 28416
rect 25320 28432 25372 28484
rect 25412 28432 25464 28484
rect 26332 28500 26384 28552
rect 27528 28543 27580 28552
rect 27528 28509 27535 28543
rect 27535 28509 27580 28543
rect 27528 28500 27580 28509
rect 26976 28432 27028 28484
rect 27712 28636 27764 28688
rect 28172 28636 28224 28688
rect 30656 28679 30708 28688
rect 30656 28645 30665 28679
rect 30665 28645 30699 28679
rect 30699 28645 30708 28679
rect 30656 28636 30708 28645
rect 27988 28568 28040 28620
rect 28632 28611 28684 28620
rect 27804 28543 27856 28552
rect 27804 28509 27818 28543
rect 27818 28509 27852 28543
rect 27852 28509 27856 28543
rect 27804 28500 27856 28509
rect 28172 28500 28224 28552
rect 28632 28577 28641 28611
rect 28641 28577 28675 28611
rect 28675 28577 28684 28611
rect 28632 28568 28684 28577
rect 28540 28543 28592 28552
rect 28540 28509 28549 28543
rect 28549 28509 28583 28543
rect 28583 28509 28592 28543
rect 28540 28500 28592 28509
rect 28724 28500 28776 28552
rect 31392 28568 31444 28620
rect 30564 28543 30616 28552
rect 30564 28509 30573 28543
rect 30573 28509 30607 28543
rect 30607 28509 30616 28543
rect 30564 28500 30616 28509
rect 31576 28543 31628 28552
rect 31576 28509 31585 28543
rect 31585 28509 31619 28543
rect 31619 28509 31628 28543
rect 31576 28500 31628 28509
rect 32036 28500 32088 28552
rect 34612 28500 34664 28552
rect 33416 28475 33468 28484
rect 33416 28441 33425 28475
rect 33425 28441 33459 28475
rect 33459 28441 33468 28475
rect 33416 28432 33468 28441
rect 33508 28432 33560 28484
rect 35348 28500 35400 28552
rect 46940 28500 46992 28552
rect 30380 28364 30432 28416
rect 31392 28364 31444 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 1768 28160 1820 28212
rect 14096 28160 14148 28212
rect 14188 28160 14240 28212
rect 16304 28160 16356 28212
rect 20536 28203 20588 28212
rect 20536 28169 20545 28203
rect 20545 28169 20579 28203
rect 20579 28169 20588 28203
rect 20536 28160 20588 28169
rect 21180 28203 21232 28212
rect 21180 28169 21189 28203
rect 21189 28169 21223 28203
rect 21223 28169 21232 28203
rect 21180 28160 21232 28169
rect 21364 28160 21416 28212
rect 22376 28160 22428 28212
rect 25412 28160 25464 28212
rect 25596 28203 25648 28212
rect 25596 28169 25605 28203
rect 25605 28169 25639 28203
rect 25639 28169 25648 28203
rect 25596 28160 25648 28169
rect 26332 28203 26384 28212
rect 26332 28169 26341 28203
rect 26341 28169 26375 28203
rect 26375 28169 26384 28203
rect 26332 28160 26384 28169
rect 27160 28203 27212 28212
rect 27160 28169 27169 28203
rect 27169 28169 27203 28203
rect 27203 28169 27212 28203
rect 27160 28160 27212 28169
rect 27436 28160 27488 28212
rect 28724 28160 28776 28212
rect 10968 28092 11020 28144
rect 15476 28092 15528 28144
rect 11336 28024 11388 28076
rect 14556 28067 14608 28076
rect 9680 27956 9732 28008
rect 7564 27888 7616 27940
rect 10784 27956 10836 28008
rect 14556 28033 14565 28067
rect 14565 28033 14599 28067
rect 14599 28033 14608 28067
rect 14556 28024 14608 28033
rect 14740 28067 14792 28076
rect 14740 28033 14749 28067
rect 14749 28033 14783 28067
rect 14783 28033 14792 28067
rect 15568 28067 15620 28076
rect 14740 28024 14792 28033
rect 15568 28033 15577 28067
rect 15577 28033 15611 28067
rect 15611 28033 15620 28067
rect 15568 28024 15620 28033
rect 15752 28067 15804 28076
rect 15752 28033 15761 28067
rect 15761 28033 15795 28067
rect 15795 28033 15804 28067
rect 15752 28024 15804 28033
rect 15936 28092 15988 28144
rect 18236 28135 18288 28144
rect 18236 28101 18245 28135
rect 18245 28101 18279 28135
rect 18279 28101 18288 28135
rect 18236 28092 18288 28101
rect 21640 28092 21692 28144
rect 16488 28024 16540 28076
rect 18052 28067 18104 28076
rect 18052 28033 18061 28067
rect 18061 28033 18095 28067
rect 18095 28033 18104 28067
rect 18052 28024 18104 28033
rect 14372 27931 14424 27940
rect 14372 27897 14381 27931
rect 14381 27897 14415 27931
rect 14415 27897 14424 27931
rect 14372 27888 14424 27897
rect 20260 28024 20312 28076
rect 20628 28024 20680 28076
rect 21088 28067 21140 28076
rect 21088 28033 21097 28067
rect 21097 28033 21131 28067
rect 21131 28033 21140 28067
rect 21088 28024 21140 28033
rect 21364 28024 21416 28076
rect 22008 28024 22060 28076
rect 22284 28067 22336 28076
rect 22284 28033 22293 28067
rect 22293 28033 22327 28067
rect 22327 28033 22336 28067
rect 27620 28092 27672 28144
rect 22284 28024 22336 28033
rect 26424 28067 26476 28076
rect 26424 28033 26433 28067
rect 26433 28033 26467 28067
rect 26467 28033 26476 28067
rect 26424 28024 26476 28033
rect 27436 28024 27488 28076
rect 27804 28092 27856 28144
rect 28080 28024 28132 28076
rect 29092 28067 29144 28076
rect 29092 28033 29101 28067
rect 29101 28033 29135 28067
rect 29135 28033 29144 28067
rect 29092 28024 29144 28033
rect 26332 27956 26384 28008
rect 27160 27956 27212 28008
rect 32312 28092 32364 28144
rect 31208 28067 31260 28076
rect 31208 28033 31217 28067
rect 31217 28033 31251 28067
rect 31251 28033 31260 28067
rect 31208 28024 31260 28033
rect 31392 28067 31444 28076
rect 31392 28033 31401 28067
rect 31401 28033 31435 28067
rect 31435 28033 31444 28067
rect 31392 28024 31444 28033
rect 31484 28067 31536 28076
rect 31484 28033 31493 28067
rect 31493 28033 31527 28067
rect 31527 28033 31536 28067
rect 31484 28024 31536 28033
rect 35348 28024 35400 28076
rect 13544 27820 13596 27872
rect 31484 27888 31536 27940
rect 33232 27999 33284 28008
rect 33232 27965 33241 27999
rect 33241 27965 33275 27999
rect 33275 27965 33284 27999
rect 33232 27956 33284 27965
rect 34704 27999 34756 28008
rect 34704 27965 34713 27999
rect 34713 27965 34747 27999
rect 34747 27965 34756 27999
rect 34704 27956 34756 27965
rect 47584 28067 47636 28076
rect 47584 28033 47593 28067
rect 47593 28033 47627 28067
rect 47627 28033 47636 28067
rect 47584 28024 47636 28033
rect 46388 27956 46440 28008
rect 23112 27863 23164 27872
rect 23112 27829 23121 27863
rect 23121 27829 23155 27863
rect 23155 27829 23164 27863
rect 23112 27820 23164 27829
rect 25688 27820 25740 27872
rect 27068 27820 27120 27872
rect 28172 27820 28224 27872
rect 30748 27820 30800 27872
rect 31024 27863 31076 27872
rect 31024 27829 31033 27863
rect 31033 27829 31067 27863
rect 31067 27829 31076 27863
rect 31024 27820 31076 27829
rect 47676 27863 47728 27872
rect 47676 27829 47685 27863
rect 47685 27829 47719 27863
rect 47719 27829 47728 27863
rect 47676 27820 47728 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3976 27616 4028 27668
rect 9680 27591 9732 27600
rect 9680 27557 9689 27591
rect 9689 27557 9723 27591
rect 9723 27557 9732 27591
rect 9680 27548 9732 27557
rect 11980 27548 12032 27600
rect 15752 27548 15804 27600
rect 17868 27548 17920 27600
rect 21180 27616 21232 27668
rect 21548 27659 21600 27668
rect 21548 27625 21557 27659
rect 21557 27625 21591 27659
rect 21591 27625 21600 27659
rect 21548 27616 21600 27625
rect 26424 27616 26476 27668
rect 28448 27616 28500 27668
rect 28540 27616 28592 27668
rect 33508 27616 33560 27668
rect 33876 27616 33928 27668
rect 16672 27523 16724 27532
rect 16672 27489 16681 27523
rect 16681 27489 16715 27523
rect 16715 27489 16724 27523
rect 16672 27480 16724 27489
rect 24216 27548 24268 27600
rect 27252 27548 27304 27600
rect 20996 27480 21048 27532
rect 23296 27523 23348 27532
rect 9588 27455 9640 27464
rect 9588 27421 9597 27455
rect 9597 27421 9631 27455
rect 9631 27421 9640 27455
rect 9588 27412 9640 27421
rect 10968 27412 11020 27464
rect 12624 27412 12676 27464
rect 13360 27455 13412 27464
rect 13360 27421 13369 27455
rect 13369 27421 13403 27455
rect 13403 27421 13412 27455
rect 13360 27412 13412 27421
rect 14096 27455 14148 27464
rect 14096 27421 14105 27455
rect 14105 27421 14139 27455
rect 14139 27421 14148 27455
rect 14096 27412 14148 27421
rect 16396 27455 16448 27464
rect 16396 27421 16405 27455
rect 16405 27421 16439 27455
rect 16439 27421 16448 27455
rect 16396 27412 16448 27421
rect 17776 27412 17828 27464
rect 11520 27344 11572 27396
rect 21088 27412 21140 27464
rect 21272 27412 21324 27464
rect 22376 27455 22428 27464
rect 22376 27421 22385 27455
rect 22385 27421 22419 27455
rect 22419 27421 22428 27455
rect 22376 27412 22428 27421
rect 23296 27489 23305 27523
rect 23305 27489 23339 27523
rect 23339 27489 23348 27523
rect 23296 27480 23348 27489
rect 10876 27276 10928 27328
rect 13636 27276 13688 27328
rect 15384 27276 15436 27328
rect 16488 27276 16540 27328
rect 18052 27276 18104 27328
rect 20904 27319 20956 27328
rect 20904 27285 20913 27319
rect 20913 27285 20947 27319
rect 20947 27285 20956 27319
rect 20904 27276 20956 27285
rect 21364 27387 21416 27396
rect 21364 27353 21373 27387
rect 21373 27353 21407 27387
rect 21407 27353 21416 27387
rect 21364 27344 21416 27353
rect 24860 27455 24912 27464
rect 24860 27421 24869 27455
rect 24869 27421 24903 27455
rect 24903 27421 24912 27455
rect 24860 27412 24912 27421
rect 26148 27455 26200 27464
rect 26148 27421 26157 27455
rect 26157 27421 26191 27455
rect 26191 27421 26200 27455
rect 26148 27412 26200 27421
rect 27068 27412 27120 27464
rect 29092 27548 29144 27600
rect 30748 27591 30800 27600
rect 27620 27480 27672 27532
rect 28264 27412 28316 27464
rect 28540 27412 28592 27464
rect 30748 27557 30757 27591
rect 30757 27557 30791 27591
rect 30791 27557 30800 27591
rect 30748 27548 30800 27557
rect 33232 27548 33284 27600
rect 29828 27412 29880 27464
rect 21640 27276 21692 27328
rect 21824 27319 21876 27328
rect 21824 27285 21833 27319
rect 21833 27285 21867 27319
rect 21867 27285 21876 27319
rect 21824 27276 21876 27285
rect 22100 27276 22152 27328
rect 24952 27344 25004 27396
rect 25136 27344 25188 27396
rect 26700 27344 26752 27396
rect 27988 27344 28040 27396
rect 28172 27387 28224 27396
rect 28172 27353 28181 27387
rect 28181 27353 28215 27387
rect 28215 27353 28224 27387
rect 28172 27344 28224 27353
rect 28724 27387 28776 27396
rect 28724 27353 28733 27387
rect 28733 27353 28767 27387
rect 28767 27353 28776 27387
rect 28724 27344 28776 27353
rect 31116 27480 31168 27532
rect 46940 27548 46992 27600
rect 47676 27480 47728 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 26240 27319 26292 27328
rect 26240 27285 26249 27319
rect 26249 27285 26283 27319
rect 26283 27285 26292 27319
rect 26240 27276 26292 27285
rect 28448 27276 28500 27328
rect 31024 27412 31076 27464
rect 31668 27455 31720 27464
rect 31668 27421 31675 27455
rect 31675 27421 31720 27455
rect 31668 27412 31720 27421
rect 31944 27455 31996 27464
rect 31944 27421 31958 27455
rect 31958 27421 31992 27455
rect 31992 27421 31996 27455
rect 31944 27412 31996 27421
rect 30748 27344 30800 27396
rect 31300 27344 31352 27396
rect 31852 27387 31904 27396
rect 31852 27353 31861 27387
rect 31861 27353 31895 27387
rect 31895 27353 31904 27387
rect 31852 27344 31904 27353
rect 30656 27276 30708 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 10968 27072 11020 27124
rect 13636 27072 13688 27124
rect 15292 27115 15344 27124
rect 15292 27081 15301 27115
rect 15301 27081 15335 27115
rect 15335 27081 15344 27115
rect 15292 27072 15344 27081
rect 15936 27072 15988 27124
rect 17316 27072 17368 27124
rect 19248 27072 19300 27124
rect 21824 27072 21876 27124
rect 24492 27072 24544 27124
rect 26148 27072 26200 27124
rect 27252 27072 27304 27124
rect 28540 27072 28592 27124
rect 28724 27072 28776 27124
rect 29276 27115 29328 27124
rect 29276 27081 29285 27115
rect 29285 27081 29319 27115
rect 29319 27081 29328 27115
rect 29276 27072 29328 27081
rect 31300 27072 31352 27124
rect 7472 27004 7524 27056
rect 18052 27047 18104 27056
rect 10784 26936 10836 26988
rect 10968 26936 11020 26988
rect 12624 26936 12676 26988
rect 13912 26979 13964 26988
rect 13912 26945 13921 26979
rect 13921 26945 13955 26979
rect 13955 26945 13964 26979
rect 13912 26936 13964 26945
rect 14096 26936 14148 26988
rect 14924 26936 14976 26988
rect 15384 26979 15436 26988
rect 15384 26945 15393 26979
rect 15393 26945 15427 26979
rect 15427 26945 15436 26979
rect 15384 26936 15436 26945
rect 15200 26868 15252 26920
rect 16396 26936 16448 26988
rect 16672 26936 16724 26988
rect 18052 27013 18061 27047
rect 18061 27013 18095 27047
rect 18095 27013 18104 27047
rect 18052 27004 18104 27013
rect 20628 27004 20680 27056
rect 17868 26979 17920 26988
rect 17868 26945 17877 26979
rect 17877 26945 17911 26979
rect 17911 26945 17920 26979
rect 17868 26936 17920 26945
rect 23112 27004 23164 27056
rect 27620 27047 27672 27056
rect 20076 26868 20128 26920
rect 20904 26936 20956 26988
rect 22008 26979 22060 26988
rect 22008 26945 22017 26979
rect 22017 26945 22051 26979
rect 22051 26945 22060 26979
rect 22008 26936 22060 26945
rect 22100 26979 22152 26988
rect 22100 26945 22109 26979
rect 22109 26945 22143 26979
rect 22143 26945 22152 26979
rect 22100 26936 22152 26945
rect 22652 26936 22704 26988
rect 24308 26979 24360 26988
rect 24308 26945 24317 26979
rect 24317 26945 24351 26979
rect 24351 26945 24360 26979
rect 24308 26936 24360 26945
rect 25688 26979 25740 26988
rect 25688 26945 25697 26979
rect 25697 26945 25731 26979
rect 25731 26945 25740 26979
rect 25688 26936 25740 26945
rect 24860 26868 24912 26920
rect 9588 26800 9640 26852
rect 10600 26732 10652 26784
rect 11612 26732 11664 26784
rect 14556 26800 14608 26852
rect 15660 26732 15712 26784
rect 15844 26775 15896 26784
rect 15844 26741 15853 26775
rect 15853 26741 15887 26775
rect 15887 26741 15896 26775
rect 15844 26732 15896 26741
rect 20628 26732 20680 26784
rect 20812 26775 20864 26784
rect 20812 26741 20821 26775
rect 20821 26741 20855 26775
rect 20855 26741 20864 26775
rect 20812 26732 20864 26741
rect 22560 26775 22612 26784
rect 22560 26741 22569 26775
rect 22569 26741 22603 26775
rect 22603 26741 22612 26775
rect 22560 26732 22612 26741
rect 23848 26775 23900 26784
rect 23848 26741 23857 26775
rect 23857 26741 23891 26775
rect 23891 26741 23900 26775
rect 23848 26732 23900 26741
rect 24216 26843 24268 26852
rect 24216 26809 24225 26843
rect 24225 26809 24259 26843
rect 24259 26809 24268 26843
rect 24216 26800 24268 26809
rect 24676 26800 24728 26852
rect 24584 26732 24636 26784
rect 27620 27013 27629 27047
rect 27629 27013 27663 27047
rect 27663 27013 27672 27047
rect 27620 27004 27672 27013
rect 27988 27004 28040 27056
rect 31024 27004 31076 27056
rect 31116 27004 31168 27056
rect 27252 26868 27304 26920
rect 29184 26979 29236 26988
rect 29184 26945 29193 26979
rect 29193 26945 29227 26979
rect 29227 26945 29236 26979
rect 29184 26936 29236 26945
rect 27988 26868 28040 26920
rect 28632 26868 28684 26920
rect 31208 26936 31260 26988
rect 31576 26868 31628 26920
rect 33140 27004 33192 27056
rect 33508 27004 33560 27056
rect 32496 26936 32548 26988
rect 33416 26979 33468 26988
rect 26240 26800 26292 26852
rect 33416 26945 33425 26979
rect 33425 26945 33459 26979
rect 33459 26945 33468 26979
rect 33416 26936 33468 26945
rect 33968 26979 34020 26988
rect 33968 26945 33977 26979
rect 33977 26945 34011 26979
rect 34011 26945 34020 26979
rect 33968 26936 34020 26945
rect 32956 26868 33008 26920
rect 40408 26868 40460 26920
rect 27344 26732 27396 26784
rect 27804 26775 27856 26784
rect 27804 26741 27813 26775
rect 27813 26741 27847 26775
rect 27847 26741 27856 26775
rect 27804 26732 27856 26741
rect 27988 26775 28040 26784
rect 27988 26741 27997 26775
rect 27997 26741 28031 26775
rect 28031 26741 28040 26775
rect 27988 26732 28040 26741
rect 29920 26732 29972 26784
rect 31024 26732 31076 26784
rect 33324 26732 33376 26784
rect 34704 26732 34756 26784
rect 46296 26732 46348 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 11336 26528 11388 26580
rect 12348 26571 12400 26580
rect 12348 26537 12357 26571
rect 12357 26537 12391 26571
rect 12391 26537 12400 26571
rect 12348 26528 12400 26537
rect 14740 26528 14792 26580
rect 14924 26528 14976 26580
rect 22560 26528 22612 26580
rect 27068 26571 27120 26580
rect 10600 26435 10652 26444
rect 10600 26401 10609 26435
rect 10609 26401 10643 26435
rect 10643 26401 10652 26435
rect 10600 26392 10652 26401
rect 10876 26435 10928 26444
rect 10876 26401 10885 26435
rect 10885 26401 10919 26435
rect 10919 26401 10928 26435
rect 10876 26392 10928 26401
rect 15844 26392 15896 26444
rect 19432 26392 19484 26444
rect 22284 26460 22336 26512
rect 24584 26460 24636 26512
rect 27068 26537 27077 26571
rect 27077 26537 27111 26571
rect 27111 26537 27120 26571
rect 27068 26528 27120 26537
rect 27252 26571 27304 26580
rect 27252 26537 27261 26571
rect 27261 26537 27295 26571
rect 27295 26537 27304 26571
rect 27252 26528 27304 26537
rect 27988 26528 28040 26580
rect 31392 26528 31444 26580
rect 31576 26528 31628 26580
rect 27160 26460 27212 26512
rect 27344 26460 27396 26512
rect 14188 26367 14240 26376
rect 14188 26333 14197 26367
rect 14197 26333 14231 26367
rect 14231 26333 14240 26367
rect 14188 26324 14240 26333
rect 14740 26324 14792 26376
rect 21640 26392 21692 26444
rect 21916 26392 21968 26444
rect 22008 26324 22060 26376
rect 24676 26367 24728 26376
rect 24676 26333 24685 26367
rect 24685 26333 24719 26367
rect 24719 26333 24728 26367
rect 24676 26324 24728 26333
rect 24860 26367 24912 26376
rect 24860 26333 24869 26367
rect 24869 26333 24903 26367
rect 24903 26333 24912 26367
rect 24860 26324 24912 26333
rect 26700 26367 26752 26376
rect 26700 26333 26709 26367
rect 26709 26333 26743 26367
rect 26743 26333 26752 26367
rect 26700 26324 26752 26333
rect 27160 26324 27212 26376
rect 28540 26392 28592 26444
rect 28724 26324 28776 26376
rect 30380 26460 30432 26512
rect 32496 26460 32548 26512
rect 29644 26392 29696 26444
rect 31024 26392 31076 26444
rect 31392 26392 31444 26444
rect 33416 26392 33468 26444
rect 33692 26435 33744 26444
rect 33692 26401 33701 26435
rect 33701 26401 33735 26435
rect 33735 26401 33744 26435
rect 46296 26435 46348 26444
rect 33692 26392 33744 26401
rect 46296 26401 46305 26435
rect 46305 26401 46339 26435
rect 46339 26401 46348 26435
rect 46296 26392 46348 26401
rect 11612 26256 11664 26308
rect 15384 26299 15436 26308
rect 15384 26265 15393 26299
rect 15393 26265 15427 26299
rect 15427 26265 15436 26299
rect 15384 26256 15436 26265
rect 16028 26256 16080 26308
rect 20812 26256 20864 26308
rect 21088 26256 21140 26308
rect 13360 26188 13412 26240
rect 17776 26188 17828 26240
rect 21364 26256 21416 26308
rect 21916 26256 21968 26308
rect 23664 26299 23716 26308
rect 23664 26265 23673 26299
rect 23673 26265 23707 26299
rect 23707 26265 23716 26299
rect 23664 26256 23716 26265
rect 24308 26256 24360 26308
rect 25504 26256 25556 26308
rect 26332 26256 26384 26308
rect 29184 26256 29236 26308
rect 25044 26231 25096 26240
rect 25044 26197 25053 26231
rect 25053 26197 25087 26231
rect 25087 26197 25096 26231
rect 25044 26188 25096 26197
rect 29920 26367 29972 26376
rect 29920 26333 29929 26367
rect 29929 26333 29963 26367
rect 29963 26333 29972 26367
rect 30196 26367 30248 26376
rect 29920 26324 29972 26333
rect 30196 26333 30221 26367
rect 30221 26333 30248 26367
rect 30196 26324 30248 26333
rect 33324 26367 33376 26376
rect 33324 26333 33333 26367
rect 33333 26333 33367 26367
rect 33367 26333 33376 26367
rect 33324 26324 33376 26333
rect 33508 26367 33560 26376
rect 33508 26333 33517 26367
rect 33517 26333 33551 26367
rect 33551 26333 33560 26367
rect 33508 26324 33560 26333
rect 33600 26367 33652 26376
rect 33600 26333 33609 26367
rect 33609 26333 33643 26367
rect 33643 26333 33652 26367
rect 33600 26324 33652 26333
rect 33968 26324 34020 26376
rect 32588 26256 32640 26308
rect 46848 26256 46900 26308
rect 48228 26256 48280 26308
rect 30196 26188 30248 26240
rect 34060 26231 34112 26240
rect 34060 26197 34069 26231
rect 34069 26197 34103 26231
rect 34103 26197 34112 26231
rect 34060 26188 34112 26197
rect 46388 26188 46440 26240
rect 46756 26188 46808 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 14188 25984 14240 26036
rect 15292 26027 15344 26036
rect 15292 25993 15301 26027
rect 15301 25993 15335 26027
rect 15335 25993 15344 26027
rect 15292 25984 15344 25993
rect 16028 26027 16080 26036
rect 16028 25993 16037 26027
rect 16037 25993 16071 26027
rect 16071 25993 16080 26027
rect 16028 25984 16080 25993
rect 17776 25984 17828 26036
rect 23848 26027 23900 26036
rect 23848 25993 23857 26027
rect 23857 25993 23891 26027
rect 23891 25993 23900 26027
rect 23848 25984 23900 25993
rect 25504 25984 25556 26036
rect 29644 25984 29696 26036
rect 31300 26027 31352 26036
rect 31300 25993 31309 26027
rect 31309 25993 31343 26027
rect 31343 25993 31352 26027
rect 31300 25984 31352 25993
rect 32588 26027 32640 26036
rect 32588 25993 32597 26027
rect 32597 25993 32631 26027
rect 32631 25993 32640 26027
rect 32588 25984 32640 25993
rect 33600 25984 33652 26036
rect 47768 25984 47820 26036
rect 11428 25916 11480 25968
rect 12348 25916 12400 25968
rect 14280 25916 14332 25968
rect 14924 25959 14976 25968
rect 14924 25925 14933 25959
rect 14933 25925 14967 25959
rect 14967 25925 14976 25959
rect 14924 25916 14976 25925
rect 10968 25848 11020 25900
rect 11336 25848 11388 25900
rect 11888 25848 11940 25900
rect 14188 25891 14240 25900
rect 14188 25857 14197 25891
rect 14197 25857 14231 25891
rect 14231 25857 14240 25891
rect 14188 25848 14240 25857
rect 14740 25848 14792 25900
rect 16672 25848 16724 25900
rect 17224 25891 17276 25900
rect 17224 25857 17233 25891
rect 17233 25857 17267 25891
rect 17267 25857 17276 25891
rect 17224 25848 17276 25857
rect 20996 25891 21048 25900
rect 20996 25857 21005 25891
rect 21005 25857 21039 25891
rect 21039 25857 21048 25891
rect 20996 25848 21048 25857
rect 21272 25891 21324 25900
rect 21272 25857 21281 25891
rect 21281 25857 21315 25891
rect 21315 25857 21324 25891
rect 21272 25848 21324 25857
rect 21364 25780 21416 25832
rect 11520 25755 11572 25764
rect 11520 25721 11529 25755
rect 11529 25721 11563 25755
rect 11563 25721 11572 25755
rect 11520 25712 11572 25721
rect 14188 25712 14240 25764
rect 19248 25712 19300 25764
rect 21548 25712 21600 25764
rect 24216 25848 24268 25900
rect 24584 25891 24636 25900
rect 24584 25857 24593 25891
rect 24593 25857 24627 25891
rect 24627 25857 24636 25891
rect 24584 25848 24636 25857
rect 24676 25891 24728 25900
rect 24676 25857 24685 25891
rect 24685 25857 24719 25891
rect 24719 25857 24728 25891
rect 24676 25848 24728 25857
rect 24860 25823 24912 25832
rect 24860 25789 24869 25823
rect 24869 25789 24903 25823
rect 24903 25789 24912 25823
rect 24860 25780 24912 25789
rect 25688 25712 25740 25764
rect 27252 25848 27304 25900
rect 28632 25891 28684 25900
rect 28632 25857 28641 25891
rect 28641 25857 28675 25891
rect 28675 25857 28684 25891
rect 28632 25848 28684 25857
rect 31392 25916 31444 25968
rect 34060 25916 34112 25968
rect 34612 25916 34664 25968
rect 31576 25848 31628 25900
rect 33784 25848 33836 25900
rect 46664 25848 46716 25900
rect 31484 25780 31536 25832
rect 33876 25823 33928 25832
rect 33876 25789 33885 25823
rect 33885 25789 33919 25823
rect 33919 25789 33928 25823
rect 33876 25780 33928 25789
rect 45836 25780 45888 25832
rect 46388 25780 46440 25832
rect 33048 25712 33100 25764
rect 46296 25712 46348 25764
rect 9680 25644 9732 25696
rect 11428 25644 11480 25696
rect 14556 25644 14608 25696
rect 20536 25687 20588 25696
rect 20536 25653 20545 25687
rect 20545 25653 20579 25687
rect 20579 25653 20588 25687
rect 20536 25644 20588 25653
rect 22376 25644 22428 25696
rect 24768 25687 24820 25696
rect 24768 25653 24777 25687
rect 24777 25653 24811 25687
rect 24811 25653 24820 25687
rect 24768 25644 24820 25653
rect 26608 25644 26660 25696
rect 27160 25687 27212 25696
rect 27160 25653 27169 25687
rect 27169 25653 27203 25687
rect 27203 25653 27212 25687
rect 27160 25644 27212 25653
rect 31024 25644 31076 25696
rect 31484 25644 31536 25696
rect 46480 25644 46532 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 14280 25483 14332 25492
rect 2320 25304 2372 25356
rect 10968 25372 11020 25424
rect 14280 25449 14289 25483
rect 14289 25449 14323 25483
rect 14323 25449 14332 25483
rect 14280 25440 14332 25449
rect 15200 25440 15252 25492
rect 15384 25440 15436 25492
rect 25688 25440 25740 25492
rect 27436 25440 27488 25492
rect 31576 25483 31628 25492
rect 31576 25449 31585 25483
rect 31585 25449 31619 25483
rect 31619 25449 31628 25483
rect 31576 25440 31628 25449
rect 34244 25440 34296 25492
rect 43352 25440 43404 25492
rect 23664 25372 23716 25424
rect 24676 25372 24728 25424
rect 9680 25347 9732 25356
rect 9680 25313 9689 25347
rect 9689 25313 9723 25347
rect 9723 25313 9732 25347
rect 9680 25304 9732 25313
rect 1860 25279 1912 25288
rect 1860 25245 1869 25279
rect 1869 25245 1903 25279
rect 1903 25245 1912 25279
rect 1860 25236 1912 25245
rect 12348 25304 12400 25356
rect 12624 25279 12676 25288
rect 12624 25245 12633 25279
rect 12633 25245 12667 25279
rect 12667 25245 12676 25279
rect 12624 25236 12676 25245
rect 13268 25236 13320 25288
rect 13452 25236 13504 25288
rect 13544 25236 13596 25288
rect 20536 25304 20588 25356
rect 22376 25347 22428 25356
rect 22376 25313 22385 25347
rect 22385 25313 22419 25347
rect 22419 25313 22428 25347
rect 22376 25304 22428 25313
rect 9956 25211 10008 25220
rect 9956 25177 9965 25211
rect 9965 25177 9999 25211
rect 9999 25177 10008 25211
rect 9956 25168 10008 25177
rect 14188 25168 14240 25220
rect 14740 25168 14792 25220
rect 15660 25279 15712 25288
rect 15660 25245 15669 25279
rect 15669 25245 15703 25279
rect 15703 25245 15712 25279
rect 15660 25236 15712 25245
rect 15844 25279 15896 25288
rect 15844 25245 15853 25279
rect 15853 25245 15887 25279
rect 15887 25245 15896 25279
rect 15844 25236 15896 25245
rect 23480 25236 23532 25288
rect 24768 25304 24820 25356
rect 25044 25236 25096 25288
rect 25780 25304 25832 25356
rect 28172 25304 28224 25356
rect 34612 25372 34664 25424
rect 25688 25236 25740 25288
rect 28540 25236 28592 25288
rect 29276 25236 29328 25288
rect 29644 25236 29696 25288
rect 29920 25279 29972 25288
rect 29920 25245 29929 25279
rect 29929 25245 29963 25279
rect 29963 25245 29972 25279
rect 31208 25304 31260 25356
rect 33876 25304 33928 25356
rect 46480 25347 46532 25356
rect 46480 25313 46489 25347
rect 46489 25313 46523 25347
rect 46523 25313 46532 25347
rect 46480 25304 46532 25313
rect 48136 25347 48188 25356
rect 48136 25313 48145 25347
rect 48145 25313 48179 25347
rect 48179 25313 48188 25347
rect 48136 25304 48188 25313
rect 29920 25236 29972 25245
rect 30288 25236 30340 25288
rect 32496 25236 32548 25288
rect 33784 25236 33836 25288
rect 45468 25279 45520 25288
rect 45468 25245 45477 25279
rect 45477 25245 45511 25279
rect 45511 25245 45520 25279
rect 45468 25236 45520 25245
rect 22284 25168 22336 25220
rect 1860 25100 1912 25152
rect 10876 25100 10928 25152
rect 13636 25100 13688 25152
rect 14464 25143 14516 25152
rect 14464 25109 14473 25143
rect 14473 25109 14507 25143
rect 14507 25109 14516 25143
rect 14464 25100 14516 25109
rect 16672 25143 16724 25152
rect 16672 25109 16681 25143
rect 16681 25109 16715 25143
rect 16715 25109 16724 25143
rect 16672 25100 16724 25109
rect 17960 25100 18012 25152
rect 21732 25100 21784 25152
rect 28816 25168 28868 25220
rect 29368 25168 29420 25220
rect 30656 25168 30708 25220
rect 31576 25168 31628 25220
rect 34704 25168 34756 25220
rect 35992 25168 36044 25220
rect 46480 25168 46532 25220
rect 25412 25143 25464 25152
rect 25412 25109 25421 25143
rect 25421 25109 25455 25143
rect 25455 25109 25464 25143
rect 25412 25100 25464 25109
rect 25872 25100 25924 25152
rect 29644 25143 29696 25152
rect 29644 25109 29653 25143
rect 29653 25109 29687 25143
rect 29687 25109 29696 25143
rect 29644 25100 29696 25109
rect 31852 25143 31904 25152
rect 31852 25109 31861 25143
rect 31861 25109 31895 25143
rect 31895 25109 31904 25143
rect 31852 25100 31904 25109
rect 32956 25100 33008 25152
rect 45560 25143 45612 25152
rect 45560 25109 45569 25143
rect 45569 25109 45603 25143
rect 45603 25109 45612 25143
rect 45560 25100 45612 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 25872 24896 25924 24948
rect 10876 24828 10928 24880
rect 13636 24871 13688 24880
rect 13636 24837 13645 24871
rect 13645 24837 13679 24871
rect 13679 24837 13688 24871
rect 13636 24828 13688 24837
rect 17960 24828 18012 24880
rect 21272 24871 21324 24880
rect 21272 24837 21281 24871
rect 21281 24837 21315 24871
rect 21315 24837 21324 24871
rect 21272 24828 21324 24837
rect 25780 24828 25832 24880
rect 26148 24871 26200 24880
rect 26148 24837 26157 24871
rect 26157 24837 26191 24871
rect 26191 24837 26200 24871
rect 29920 24896 29972 24948
rect 30012 24896 30064 24948
rect 30288 24896 30340 24948
rect 26148 24828 26200 24837
rect 23020 24803 23072 24812
rect 8392 24735 8444 24744
rect 8392 24701 8401 24735
rect 8401 24701 8435 24735
rect 8435 24701 8444 24735
rect 8392 24692 8444 24701
rect 8760 24692 8812 24744
rect 3608 24556 3660 24608
rect 11796 24692 11848 24744
rect 11428 24624 11480 24676
rect 23020 24769 23029 24803
rect 23029 24769 23063 24803
rect 23063 24769 23072 24803
rect 23020 24760 23072 24769
rect 23480 24760 23532 24812
rect 24676 24803 24728 24812
rect 24676 24769 24685 24803
rect 24685 24769 24719 24803
rect 24719 24769 24728 24803
rect 24676 24760 24728 24769
rect 24952 24803 25004 24812
rect 24952 24769 24961 24803
rect 24961 24769 24995 24803
rect 24995 24769 25004 24803
rect 24952 24760 25004 24769
rect 25688 24760 25740 24812
rect 26424 24760 26476 24812
rect 29644 24828 29696 24880
rect 27988 24803 28040 24812
rect 27988 24769 27997 24803
rect 27997 24769 28031 24803
rect 28031 24769 28040 24803
rect 27988 24760 28040 24769
rect 28540 24760 28592 24812
rect 14372 24692 14424 24744
rect 14556 24735 14608 24744
rect 14556 24701 14565 24735
rect 14565 24701 14599 24735
rect 14599 24701 14608 24735
rect 14556 24692 14608 24701
rect 17040 24692 17092 24744
rect 18052 24692 18104 24744
rect 18972 24735 19024 24744
rect 18972 24701 18981 24735
rect 18981 24701 19015 24735
rect 19015 24701 19024 24735
rect 18972 24692 19024 24701
rect 19616 24735 19668 24744
rect 19616 24701 19625 24735
rect 19625 24701 19659 24735
rect 19659 24701 19668 24735
rect 19616 24692 19668 24701
rect 28264 24692 28316 24744
rect 29276 24803 29328 24812
rect 29276 24769 29285 24803
rect 29285 24769 29319 24803
rect 29319 24769 29328 24803
rect 29276 24760 29328 24769
rect 29920 24760 29972 24812
rect 32956 24896 33008 24948
rect 30564 24828 30616 24880
rect 31208 24871 31260 24880
rect 31208 24837 31217 24871
rect 31217 24837 31251 24871
rect 31251 24837 31260 24871
rect 31208 24828 31260 24837
rect 35716 24871 35768 24880
rect 35716 24837 35725 24871
rect 35725 24837 35759 24871
rect 35759 24837 35768 24871
rect 35716 24828 35768 24837
rect 31300 24760 31352 24812
rect 33784 24760 33836 24812
rect 35992 24760 36044 24812
rect 30564 24735 30616 24744
rect 30564 24701 30573 24735
rect 30573 24701 30607 24735
rect 30607 24701 30616 24735
rect 30564 24692 30616 24701
rect 40040 24735 40092 24744
rect 12624 24624 12676 24676
rect 14464 24624 14516 24676
rect 25872 24624 25924 24676
rect 27896 24624 27948 24676
rect 11612 24556 11664 24608
rect 11980 24556 12032 24608
rect 23020 24556 23072 24608
rect 25964 24556 26016 24608
rect 28080 24556 28132 24608
rect 30380 24556 30432 24608
rect 30472 24599 30524 24608
rect 30472 24565 30481 24599
rect 30481 24565 30515 24599
rect 30515 24565 30524 24599
rect 33048 24624 33100 24676
rect 35716 24624 35768 24676
rect 40040 24701 40049 24735
rect 40049 24701 40083 24735
rect 40083 24701 40092 24735
rect 40040 24692 40092 24701
rect 40316 24692 40368 24744
rect 40408 24692 40460 24744
rect 42892 24760 42944 24812
rect 43628 24803 43680 24812
rect 43628 24769 43637 24803
rect 43637 24769 43671 24803
rect 43671 24769 43680 24803
rect 43628 24760 43680 24769
rect 45468 24828 45520 24880
rect 44548 24760 44600 24812
rect 45560 24760 45612 24812
rect 44272 24692 44324 24744
rect 46848 24760 46900 24812
rect 47124 24760 47176 24812
rect 46848 24624 46900 24676
rect 31392 24599 31444 24608
rect 30472 24556 30524 24565
rect 31392 24565 31401 24599
rect 31401 24565 31435 24599
rect 31435 24565 31444 24599
rect 31392 24556 31444 24565
rect 36360 24599 36412 24608
rect 36360 24565 36369 24599
rect 36369 24565 36403 24599
rect 36403 24565 36412 24599
rect 36360 24556 36412 24565
rect 43904 24556 43956 24608
rect 46388 24556 46440 24608
rect 46572 24599 46624 24608
rect 46572 24565 46581 24599
rect 46581 24565 46615 24599
rect 46615 24565 46624 24599
rect 46572 24556 46624 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 9956 24352 10008 24404
rect 11796 24352 11848 24404
rect 17040 24395 17092 24404
rect 17040 24361 17049 24395
rect 17049 24361 17083 24395
rect 17083 24361 17092 24395
rect 17040 24352 17092 24361
rect 8392 24216 8444 24268
rect 10876 24259 10928 24268
rect 10876 24225 10885 24259
rect 10885 24225 10919 24259
rect 10919 24225 10928 24259
rect 10876 24216 10928 24225
rect 12440 24216 12492 24268
rect 15844 24284 15896 24336
rect 15384 24216 15436 24268
rect 11428 24148 11480 24200
rect 11612 24191 11664 24200
rect 11612 24157 11621 24191
rect 11621 24157 11655 24191
rect 11655 24157 11664 24191
rect 11612 24148 11664 24157
rect 11888 24191 11940 24200
rect 11888 24157 11897 24191
rect 11897 24157 11931 24191
rect 11931 24157 11940 24191
rect 11888 24148 11940 24157
rect 13084 24148 13136 24200
rect 13544 24148 13596 24200
rect 13636 24148 13688 24200
rect 12624 24080 12676 24132
rect 16856 24148 16908 24200
rect 19064 24352 19116 24404
rect 19616 24352 19668 24404
rect 26976 24352 27028 24404
rect 28264 24352 28316 24404
rect 28448 24352 28500 24404
rect 28632 24395 28684 24404
rect 28632 24361 28641 24395
rect 28641 24361 28675 24395
rect 28675 24361 28684 24395
rect 28632 24352 28684 24361
rect 30196 24395 30248 24404
rect 30196 24361 30205 24395
rect 30205 24361 30239 24395
rect 30239 24361 30248 24395
rect 30196 24352 30248 24361
rect 18144 24284 18196 24336
rect 18788 24216 18840 24268
rect 25504 24216 25556 24268
rect 16580 24080 16632 24132
rect 18972 24080 19024 24132
rect 11060 24012 11112 24064
rect 11428 24055 11480 24064
rect 11428 24021 11437 24055
rect 11437 24021 11471 24055
rect 11471 24021 11480 24055
rect 11428 24012 11480 24021
rect 11796 24055 11848 24064
rect 11796 24021 11805 24055
rect 11805 24021 11839 24055
rect 11839 24021 11848 24055
rect 11796 24012 11848 24021
rect 13360 24055 13412 24064
rect 13360 24021 13369 24055
rect 13369 24021 13403 24055
rect 13403 24021 13412 24055
rect 13360 24012 13412 24021
rect 15200 24012 15252 24064
rect 17684 24055 17736 24064
rect 17684 24021 17699 24055
rect 17699 24021 17733 24055
rect 17733 24021 17736 24055
rect 17684 24012 17736 24021
rect 19892 24148 19944 24200
rect 23112 24148 23164 24200
rect 25964 24191 26016 24200
rect 25964 24157 25973 24191
rect 25973 24157 26007 24191
rect 26007 24157 26016 24191
rect 25964 24148 26016 24157
rect 29552 24284 29604 24336
rect 30472 24352 30524 24404
rect 30564 24352 30616 24404
rect 36268 24352 36320 24404
rect 44272 24352 44324 24404
rect 30380 24284 30432 24336
rect 28080 24216 28132 24268
rect 40040 24284 40092 24336
rect 40868 24284 40920 24336
rect 45928 24284 45980 24336
rect 28172 24191 28224 24200
rect 20168 24123 20220 24132
rect 20168 24089 20177 24123
rect 20177 24089 20211 24123
rect 20211 24089 20220 24123
rect 20168 24080 20220 24089
rect 21824 24123 21876 24132
rect 21824 24089 21833 24123
rect 21833 24089 21867 24123
rect 21867 24089 21876 24123
rect 21824 24080 21876 24089
rect 25688 24080 25740 24132
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 26976 24080 27028 24132
rect 28540 24148 28592 24200
rect 29552 24191 29604 24200
rect 29552 24157 29561 24191
rect 29561 24157 29595 24191
rect 29595 24157 29604 24191
rect 29552 24148 29604 24157
rect 20536 24012 20588 24064
rect 23480 24055 23532 24064
rect 23480 24021 23489 24055
rect 23489 24021 23523 24055
rect 23523 24021 23532 24055
rect 23480 24012 23532 24021
rect 25504 24012 25556 24064
rect 28448 24012 28500 24064
rect 29920 24148 29972 24200
rect 30196 24191 30248 24200
rect 30196 24157 30205 24191
rect 30205 24157 30239 24191
rect 30239 24157 30248 24191
rect 30196 24148 30248 24157
rect 37096 24259 37148 24268
rect 37096 24225 37105 24259
rect 37105 24225 37139 24259
rect 37139 24225 37148 24259
rect 37096 24216 37148 24225
rect 31484 24191 31536 24200
rect 31484 24157 31493 24191
rect 31493 24157 31527 24191
rect 31527 24157 31536 24191
rect 31484 24148 31536 24157
rect 32864 24148 32916 24200
rect 36360 24191 36412 24200
rect 36360 24157 36369 24191
rect 36369 24157 36403 24191
rect 36403 24157 36412 24191
rect 36360 24148 36412 24157
rect 38752 24148 38804 24200
rect 31392 24080 31444 24132
rect 40316 24191 40368 24200
rect 40316 24157 40325 24191
rect 40325 24157 40359 24191
rect 40359 24157 40368 24191
rect 40960 24216 41012 24268
rect 43812 24216 43864 24268
rect 45560 24216 45612 24268
rect 46388 24259 46440 24268
rect 46388 24225 46397 24259
rect 46397 24225 46431 24259
rect 46431 24225 46440 24259
rect 46388 24216 46440 24225
rect 40316 24148 40368 24157
rect 43168 24148 43220 24200
rect 43444 24148 43496 24200
rect 43536 24191 43588 24200
rect 43536 24157 43545 24191
rect 43545 24157 43579 24191
rect 43579 24157 43588 24191
rect 43536 24148 43588 24157
rect 45744 24148 45796 24200
rect 46204 24191 46256 24200
rect 46204 24157 46213 24191
rect 46213 24157 46247 24191
rect 46247 24157 46256 24191
rect 46204 24148 46256 24157
rect 44548 24080 44600 24132
rect 45836 24080 45888 24132
rect 30564 24012 30616 24064
rect 36176 24012 36228 24064
rect 42524 24012 42576 24064
rect 43628 24012 43680 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 8760 23851 8812 23860
rect 8760 23817 8769 23851
rect 8769 23817 8803 23851
rect 8803 23817 8812 23851
rect 8760 23808 8812 23817
rect 11060 23808 11112 23860
rect 11888 23808 11940 23860
rect 18052 23851 18104 23860
rect 18052 23817 18061 23851
rect 18061 23817 18095 23851
rect 18095 23817 18104 23851
rect 18052 23808 18104 23817
rect 18972 23851 19024 23860
rect 18972 23817 18981 23851
rect 18981 23817 19015 23851
rect 19015 23817 19024 23851
rect 18972 23808 19024 23817
rect 19064 23851 19116 23860
rect 19064 23817 19073 23851
rect 19073 23817 19107 23851
rect 19107 23817 19116 23851
rect 19064 23808 19116 23817
rect 20168 23808 20220 23860
rect 22284 23808 22336 23860
rect 12440 23740 12492 23792
rect 18788 23740 18840 23792
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 8944 23672 8996 23724
rect 13636 23715 13688 23724
rect 13636 23681 13645 23715
rect 13645 23681 13679 23715
rect 13679 23681 13688 23715
rect 13636 23672 13688 23681
rect 16672 23715 16724 23724
rect 16672 23681 16681 23715
rect 16681 23681 16715 23715
rect 16715 23681 16724 23715
rect 16672 23672 16724 23681
rect 17684 23672 17736 23724
rect 18144 23715 18196 23724
rect 18144 23681 18153 23715
rect 18153 23681 18187 23715
rect 18187 23681 18196 23715
rect 18144 23672 18196 23681
rect 18880 23715 18932 23724
rect 18880 23681 18889 23715
rect 18889 23681 18923 23715
rect 18923 23681 18932 23715
rect 18880 23672 18932 23681
rect 19984 23715 20036 23724
rect 19984 23681 19993 23715
rect 19993 23681 20027 23715
rect 20027 23681 20036 23715
rect 19984 23672 20036 23681
rect 25136 23808 25188 23860
rect 28172 23808 28224 23860
rect 29552 23808 29604 23860
rect 31300 23808 31352 23860
rect 32864 23851 32916 23860
rect 32864 23817 32873 23851
rect 32873 23817 32907 23851
rect 32907 23817 32916 23851
rect 32864 23808 32916 23817
rect 23020 23783 23072 23792
rect 23020 23749 23029 23783
rect 23029 23749 23063 23783
rect 23063 23749 23072 23783
rect 23020 23740 23072 23749
rect 23480 23740 23532 23792
rect 13820 23647 13872 23656
rect 13820 23613 13829 23647
rect 13829 23613 13863 23647
rect 13863 23613 13872 23647
rect 13820 23604 13872 23613
rect 14096 23647 14148 23656
rect 14096 23613 14105 23647
rect 14105 23613 14139 23647
rect 14139 23613 14148 23647
rect 14096 23604 14148 23613
rect 28448 23672 28500 23724
rect 28632 23672 28684 23724
rect 29644 23672 29696 23724
rect 30104 23672 30156 23724
rect 30472 23672 30524 23724
rect 31024 23672 31076 23724
rect 33232 23740 33284 23792
rect 33784 23808 33836 23860
rect 40960 23851 41012 23860
rect 40960 23817 40969 23851
rect 40969 23817 41003 23851
rect 41003 23817 41012 23851
rect 40960 23808 41012 23817
rect 42524 23851 42576 23860
rect 42524 23817 42533 23851
rect 42533 23817 42567 23851
rect 42567 23817 42576 23851
rect 42524 23808 42576 23817
rect 43168 23851 43220 23860
rect 43168 23817 43177 23851
rect 43177 23817 43211 23851
rect 43211 23817 43220 23851
rect 43168 23808 43220 23817
rect 36268 23783 36320 23792
rect 36268 23749 36277 23783
rect 36277 23749 36311 23783
rect 36311 23749 36320 23783
rect 36268 23740 36320 23749
rect 37648 23740 37700 23792
rect 47492 23808 47544 23860
rect 23112 23604 23164 23656
rect 24860 23604 24912 23656
rect 28080 23604 28132 23656
rect 33968 23672 34020 23724
rect 36360 23672 36412 23724
rect 40592 23715 40644 23724
rect 40592 23681 40601 23715
rect 40601 23681 40635 23715
rect 40635 23681 40644 23715
rect 40592 23672 40644 23681
rect 43352 23672 43404 23724
rect 43904 23715 43956 23724
rect 43904 23681 43913 23715
rect 43913 23681 43947 23715
rect 43947 23681 43956 23715
rect 43904 23672 43956 23681
rect 46204 23740 46256 23792
rect 47768 23783 47820 23792
rect 47768 23749 47777 23783
rect 47777 23749 47811 23783
rect 47811 23749 47820 23783
rect 47768 23740 47820 23749
rect 47584 23715 47636 23724
rect 47584 23681 47593 23715
rect 47593 23681 47627 23715
rect 47627 23681 47636 23715
rect 47584 23672 47636 23681
rect 42892 23647 42944 23656
rect 1584 23579 1636 23588
rect 1584 23545 1593 23579
rect 1593 23545 1627 23579
rect 1627 23545 1636 23579
rect 1584 23536 1636 23545
rect 11428 23536 11480 23588
rect 24400 23536 24452 23588
rect 25228 23536 25280 23588
rect 26516 23536 26568 23588
rect 40408 23536 40460 23588
rect 42892 23613 42901 23647
rect 42901 23613 42935 23647
rect 42935 23613 42944 23647
rect 42892 23604 42944 23613
rect 45376 23647 45428 23656
rect 45376 23613 45385 23647
rect 45385 23613 45419 23647
rect 45419 23613 45428 23647
rect 45376 23604 45428 23613
rect 45560 23604 45612 23656
rect 48044 23536 48096 23588
rect 11704 23468 11756 23520
rect 16764 23511 16816 23520
rect 16764 23477 16773 23511
rect 16773 23477 16807 23511
rect 16807 23477 16816 23511
rect 16764 23468 16816 23477
rect 19432 23468 19484 23520
rect 22284 23468 22336 23520
rect 27160 23468 27212 23520
rect 31024 23468 31076 23520
rect 31392 23468 31444 23520
rect 44732 23468 44784 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 3884 23264 3936 23316
rect 12072 23264 12124 23316
rect 13084 23264 13136 23316
rect 13820 23264 13872 23316
rect 16580 23264 16632 23316
rect 26976 23307 27028 23316
rect 26976 23273 26985 23307
rect 26985 23273 27019 23307
rect 27019 23273 27028 23307
rect 26976 23264 27028 23273
rect 30380 23264 30432 23316
rect 31576 23264 31628 23316
rect 28816 23196 28868 23248
rect 11704 23171 11756 23180
rect 11704 23137 11713 23171
rect 11713 23137 11747 23171
rect 11747 23137 11756 23171
rect 11704 23128 11756 23137
rect 12072 23128 12124 23180
rect 23480 23128 23532 23180
rect 25504 23171 25556 23180
rect 25504 23137 25513 23171
rect 25513 23137 25547 23171
rect 25547 23137 25556 23171
rect 25504 23128 25556 23137
rect 30196 23128 30248 23180
rect 11428 23103 11480 23112
rect 11428 23069 11437 23103
rect 11437 23069 11471 23103
rect 11471 23069 11480 23103
rect 11428 23060 11480 23069
rect 13452 23060 13504 23112
rect 15108 23103 15160 23112
rect 15108 23069 15117 23103
rect 15117 23069 15151 23103
rect 15151 23069 15160 23103
rect 15108 23060 15160 23069
rect 16672 23060 16724 23112
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 20536 23060 20588 23112
rect 20904 23103 20956 23112
rect 20904 23069 20913 23103
rect 20913 23069 20947 23103
rect 20947 23069 20956 23103
rect 20904 23060 20956 23069
rect 22284 23060 22336 23112
rect 25136 23060 25188 23112
rect 27160 23060 27212 23112
rect 28264 23060 28316 23112
rect 30380 23103 30432 23112
rect 30380 23069 30389 23103
rect 30389 23069 30423 23103
rect 30423 23069 30432 23103
rect 30380 23060 30432 23069
rect 31484 23128 31536 23180
rect 36176 23171 36228 23180
rect 36176 23137 36185 23171
rect 36185 23137 36219 23171
rect 36219 23137 36228 23171
rect 36176 23128 36228 23137
rect 42892 23264 42944 23316
rect 45376 23264 45428 23316
rect 45284 23196 45336 23248
rect 40868 23171 40920 23180
rect 40868 23137 40877 23171
rect 40877 23137 40911 23171
rect 40911 23137 40920 23171
rect 40868 23128 40920 23137
rect 42064 23171 42116 23180
rect 42064 23137 42073 23171
rect 42073 23137 42107 23171
rect 42107 23137 42116 23171
rect 42064 23128 42116 23137
rect 45560 23128 45612 23180
rect 45744 23128 45796 23180
rect 46296 23171 46348 23180
rect 46296 23137 46305 23171
rect 46305 23137 46339 23171
rect 46339 23137 46348 23171
rect 46296 23128 46348 23137
rect 48136 23171 48188 23180
rect 48136 23137 48145 23171
rect 48145 23137 48179 23171
rect 48179 23137 48188 23171
rect 48136 23128 48188 23137
rect 30932 23060 30984 23112
rect 31576 23060 31628 23112
rect 35992 23103 36044 23112
rect 35992 23069 36001 23103
rect 36001 23069 36035 23103
rect 36035 23069 36044 23103
rect 35992 23060 36044 23069
rect 40408 23103 40460 23112
rect 40408 23069 40417 23103
rect 40417 23069 40451 23103
rect 40451 23069 40460 23103
rect 40408 23060 40460 23069
rect 43444 23060 43496 23112
rect 12440 22992 12492 23044
rect 15384 23035 15436 23044
rect 15384 23001 15393 23035
rect 15393 23001 15427 23035
rect 15427 23001 15436 23035
rect 15384 22992 15436 23001
rect 16764 22992 16816 23044
rect 21180 23035 21232 23044
rect 21180 23001 21189 23035
rect 21189 23001 21223 23035
rect 21223 23001 21232 23035
rect 21180 22992 21232 23001
rect 27068 22992 27120 23044
rect 30564 23035 30616 23044
rect 30564 23001 30573 23035
rect 30573 23001 30607 23035
rect 30607 23001 30616 23035
rect 30564 22992 30616 23001
rect 17500 22967 17552 22976
rect 17500 22933 17509 22967
rect 17509 22933 17543 22967
rect 17543 22933 17552 22967
rect 17500 22924 17552 22933
rect 19340 22924 19392 22976
rect 22100 22924 22152 22976
rect 28080 22924 28132 22976
rect 31208 22924 31260 22976
rect 33416 22992 33468 23044
rect 43628 22992 43680 23044
rect 45560 23035 45612 23044
rect 45560 23001 45569 23035
rect 45569 23001 45603 23035
rect 45603 23001 45612 23035
rect 45560 22992 45612 23001
rect 46940 22992 46992 23044
rect 48136 22924 48188 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 12440 22763 12492 22772
rect 12440 22729 12449 22763
rect 12449 22729 12483 22763
rect 12483 22729 12492 22763
rect 12440 22720 12492 22729
rect 17960 22720 18012 22772
rect 18880 22720 18932 22772
rect 19156 22763 19208 22772
rect 19156 22729 19165 22763
rect 19165 22729 19199 22763
rect 19199 22729 19208 22763
rect 19156 22720 19208 22729
rect 21180 22763 21232 22772
rect 21180 22729 21189 22763
rect 21189 22729 21223 22763
rect 21223 22729 21232 22763
rect 21180 22720 21232 22729
rect 27068 22763 27120 22772
rect 27068 22729 27077 22763
rect 27077 22729 27111 22763
rect 27111 22729 27120 22763
rect 27068 22720 27120 22729
rect 28264 22763 28316 22772
rect 28264 22729 28273 22763
rect 28273 22729 28307 22763
rect 28307 22729 28316 22763
rect 28264 22720 28316 22729
rect 17224 22652 17276 22704
rect 17500 22652 17552 22704
rect 18236 22652 18288 22704
rect 8944 22627 8996 22636
rect 8944 22593 8953 22627
rect 8953 22593 8987 22627
rect 8987 22593 8996 22627
rect 8944 22584 8996 22593
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 9772 22584 9824 22593
rect 11336 22584 11388 22636
rect 13360 22584 13412 22636
rect 13912 22627 13964 22636
rect 13912 22593 13921 22627
rect 13921 22593 13955 22627
rect 13955 22593 13964 22627
rect 13912 22584 13964 22593
rect 16580 22584 16632 22636
rect 18788 22584 18840 22636
rect 20904 22652 20956 22704
rect 26884 22652 26936 22704
rect 30564 22720 30616 22772
rect 31576 22763 31628 22772
rect 31576 22729 31585 22763
rect 31585 22729 31619 22763
rect 31619 22729 31628 22763
rect 31576 22720 31628 22729
rect 33416 22720 33468 22772
rect 40408 22720 40460 22772
rect 46940 22763 46992 22772
rect 46940 22729 46949 22763
rect 46949 22729 46983 22763
rect 46983 22729 46992 22763
rect 46940 22720 46992 22729
rect 48136 22763 48188 22772
rect 48136 22729 48145 22763
rect 48145 22729 48179 22763
rect 48179 22729 48188 22763
rect 48136 22720 48188 22729
rect 31208 22695 31260 22704
rect 31208 22661 31217 22695
rect 31217 22661 31251 22695
rect 31251 22661 31260 22695
rect 31208 22652 31260 22661
rect 31392 22695 31444 22704
rect 31392 22661 31401 22695
rect 31401 22661 31435 22695
rect 31435 22661 31444 22695
rect 31392 22652 31444 22661
rect 45744 22652 45796 22704
rect 47308 22652 47360 22704
rect 11060 22516 11112 22568
rect 11888 22516 11940 22568
rect 16672 22559 16724 22568
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 16948 22559 17000 22568
rect 16948 22525 16957 22559
rect 16957 22525 16991 22559
rect 16991 22525 17000 22559
rect 16948 22516 17000 22525
rect 19064 22516 19116 22568
rect 19984 22516 20036 22568
rect 22192 22584 22244 22636
rect 27344 22584 27396 22636
rect 28172 22584 28224 22636
rect 28448 22584 28500 22636
rect 28908 22627 28960 22636
rect 28908 22593 28917 22627
rect 28917 22593 28951 22627
rect 28951 22593 28960 22627
rect 28908 22584 28960 22593
rect 30196 22627 30248 22636
rect 23112 22559 23164 22568
rect 23112 22525 23121 22559
rect 23121 22525 23155 22559
rect 23155 22525 23164 22559
rect 23112 22516 23164 22525
rect 23480 22559 23532 22568
rect 23480 22525 23489 22559
rect 23489 22525 23523 22559
rect 23523 22525 23532 22559
rect 23480 22516 23532 22525
rect 9128 22380 9180 22432
rect 10140 22423 10192 22432
rect 10140 22389 10149 22423
rect 10149 22389 10183 22423
rect 10183 22389 10192 22423
rect 10140 22380 10192 22389
rect 10692 22423 10744 22432
rect 10692 22389 10701 22423
rect 10701 22389 10735 22423
rect 10735 22389 10744 22423
rect 10692 22380 10744 22389
rect 11612 22423 11664 22432
rect 11612 22389 11621 22423
rect 11621 22389 11655 22423
rect 11655 22389 11664 22423
rect 11612 22380 11664 22389
rect 14004 22380 14056 22432
rect 18512 22380 18564 22432
rect 20996 22380 21048 22432
rect 22008 22423 22060 22432
rect 22008 22389 22017 22423
rect 22017 22389 22051 22423
rect 22051 22389 22060 22423
rect 22008 22380 22060 22389
rect 23848 22448 23900 22500
rect 30196 22593 30205 22627
rect 30205 22593 30239 22627
rect 30239 22593 30248 22627
rect 30196 22584 30248 22593
rect 33232 22627 33284 22636
rect 33232 22593 33241 22627
rect 33241 22593 33275 22627
rect 33275 22593 33284 22627
rect 33232 22584 33284 22593
rect 36360 22584 36412 22636
rect 40316 22627 40368 22636
rect 40316 22593 40325 22627
rect 40325 22593 40359 22627
rect 40359 22593 40368 22627
rect 40316 22584 40368 22593
rect 29828 22516 29880 22568
rect 36636 22559 36688 22568
rect 36636 22525 36645 22559
rect 36645 22525 36679 22559
rect 36679 22525 36688 22559
rect 36636 22516 36688 22525
rect 42800 22516 42852 22568
rect 42892 22448 42944 22500
rect 43536 22448 43588 22500
rect 45560 22584 45612 22636
rect 47768 22584 47820 22636
rect 47216 22516 47268 22568
rect 47860 22559 47912 22568
rect 47860 22525 47869 22559
rect 47869 22525 47903 22559
rect 47903 22525 47912 22559
rect 47860 22516 47912 22525
rect 47952 22448 48004 22500
rect 23480 22380 23532 22432
rect 29460 22423 29512 22432
rect 29460 22389 29469 22423
rect 29469 22389 29503 22423
rect 29503 22389 29512 22423
rect 29460 22380 29512 22389
rect 40500 22423 40552 22432
rect 40500 22389 40509 22423
rect 40509 22389 40543 22423
rect 40543 22389 40552 22423
rect 40500 22380 40552 22389
rect 43720 22380 43772 22432
rect 47584 22380 47636 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 10140 22176 10192 22228
rect 16948 22176 17000 22228
rect 23112 22176 23164 22228
rect 25412 22219 25464 22228
rect 25412 22185 25442 22219
rect 25442 22185 25464 22219
rect 25412 22176 25464 22185
rect 26884 22176 26936 22228
rect 31944 22176 31996 22228
rect 10692 22040 10744 22092
rect 11060 22040 11112 22092
rect 11796 22083 11848 22092
rect 11796 22049 11805 22083
rect 11805 22049 11839 22083
rect 11839 22049 11848 22083
rect 11796 22040 11848 22049
rect 13176 22040 13228 22092
rect 42892 22108 42944 22160
rect 8944 22015 8996 22024
rect 8944 21981 8953 22015
rect 8953 21981 8987 22015
rect 8987 21981 8996 22015
rect 8944 21972 8996 21981
rect 12348 22015 12400 22024
rect 12348 21981 12357 22015
rect 12357 21981 12391 22015
rect 12391 21981 12400 22015
rect 12348 21972 12400 21981
rect 13360 22015 13412 22024
rect 13360 21981 13369 22015
rect 13369 21981 13403 22015
rect 13403 21981 13412 22015
rect 13360 21972 13412 21981
rect 14004 21972 14056 22024
rect 18144 22040 18196 22092
rect 20996 22083 21048 22092
rect 20996 22049 21005 22083
rect 21005 22049 21039 22083
rect 21039 22049 21048 22083
rect 20996 22040 21048 22049
rect 20 21904 72 21956
rect 8852 21904 8904 21956
rect 11612 21904 11664 21956
rect 8760 21836 8812 21888
rect 9772 21836 9824 21888
rect 11060 21836 11112 21888
rect 11336 21836 11388 21888
rect 13636 21904 13688 21956
rect 16212 21904 16264 21956
rect 17960 21972 18012 22024
rect 18512 21972 18564 22024
rect 19340 21972 19392 22024
rect 20812 22015 20864 22024
rect 20812 21981 20821 22015
rect 20821 21981 20855 22015
rect 20855 21981 20864 22015
rect 20812 21972 20864 21981
rect 22192 21972 22244 22024
rect 26792 22040 26844 22092
rect 28080 22040 28132 22092
rect 25136 22015 25188 22024
rect 25136 21981 25145 22015
rect 25145 21981 25179 22015
rect 25179 21981 25188 22015
rect 25136 21972 25188 21981
rect 27344 22015 27396 22024
rect 25688 21904 25740 21956
rect 27344 21981 27353 22015
rect 27353 21981 27387 22015
rect 27387 21981 27396 22015
rect 27344 21972 27396 21981
rect 42800 22083 42852 22092
rect 42800 22049 42809 22083
rect 42809 22049 42843 22083
rect 42843 22049 42852 22083
rect 42800 22040 42852 22049
rect 28816 22015 28868 22024
rect 28816 21981 28825 22015
rect 28825 21981 28859 22015
rect 28859 21981 28868 22015
rect 28816 21972 28868 21981
rect 34152 21972 34204 22024
rect 40316 22015 40368 22024
rect 40316 21981 40325 22015
rect 40325 21981 40359 22015
rect 40359 21981 40368 22015
rect 40316 21972 40368 21981
rect 40500 22015 40552 22024
rect 40500 21981 40509 22015
rect 40509 21981 40543 22015
rect 40543 21981 40552 22015
rect 40500 21972 40552 21981
rect 42616 21972 42668 22024
rect 42984 21972 43036 22024
rect 43536 22015 43588 22024
rect 14372 21836 14424 21888
rect 16856 21836 16908 21888
rect 18144 21836 18196 21888
rect 20904 21836 20956 21888
rect 22100 21836 22152 21888
rect 26792 21836 26844 21888
rect 27988 21879 28040 21888
rect 27988 21845 27997 21879
rect 27997 21845 28031 21879
rect 28031 21845 28040 21879
rect 27988 21836 28040 21845
rect 29460 21904 29512 21956
rect 43536 21981 43545 22015
rect 43545 21981 43579 22015
rect 43579 21981 43588 22015
rect 43536 21972 43588 21981
rect 46020 22015 46072 22024
rect 43812 21904 43864 21956
rect 46020 21981 46029 22015
rect 46029 21981 46063 22015
rect 46063 21981 46072 22015
rect 46020 21972 46072 21981
rect 46204 21972 46256 22024
rect 47308 22015 47360 22024
rect 47308 21981 47317 22015
rect 47317 21981 47351 22015
rect 47351 21981 47360 22015
rect 47308 21972 47360 21981
rect 48044 21904 48096 21956
rect 29276 21836 29328 21888
rect 34704 21879 34756 21888
rect 34704 21845 34713 21879
rect 34713 21845 34747 21879
rect 34747 21845 34756 21879
rect 34704 21836 34756 21845
rect 40500 21836 40552 21888
rect 43352 21836 43404 21888
rect 46388 21836 46440 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 3056 21632 3108 21684
rect 34152 21675 34204 21684
rect 8760 21607 8812 21616
rect 8760 21573 8769 21607
rect 8769 21573 8803 21607
rect 8803 21573 8812 21607
rect 8760 21564 8812 21573
rect 8944 21564 8996 21616
rect 13360 21564 13412 21616
rect 13636 21607 13688 21616
rect 11336 21496 11388 21548
rect 13636 21573 13645 21607
rect 13645 21573 13679 21607
rect 13679 21573 13688 21607
rect 13636 21564 13688 21573
rect 14372 21607 14424 21616
rect 14372 21573 14381 21607
rect 14381 21573 14415 21607
rect 14415 21573 14424 21607
rect 14372 21564 14424 21573
rect 18144 21607 18196 21616
rect 18144 21573 18153 21607
rect 18153 21573 18187 21607
rect 18187 21573 18196 21607
rect 18144 21564 18196 21573
rect 22008 21607 22060 21616
rect 22008 21573 22017 21607
rect 22017 21573 22051 21607
rect 22051 21573 22060 21607
rect 22008 21564 22060 21573
rect 27988 21564 28040 21616
rect 28172 21564 28224 21616
rect 16028 21539 16080 21548
rect 16028 21505 16037 21539
rect 16037 21505 16071 21539
rect 16071 21505 16080 21539
rect 16028 21496 16080 21505
rect 16856 21539 16908 21548
rect 16856 21505 16865 21539
rect 16865 21505 16899 21539
rect 16899 21505 16908 21539
rect 16856 21496 16908 21505
rect 19248 21496 19300 21548
rect 20904 21496 20956 21548
rect 21732 21496 21784 21548
rect 25136 21496 25188 21548
rect 32312 21539 32364 21548
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 8852 21428 8904 21480
rect 14188 21471 14240 21480
rect 14188 21437 14197 21471
rect 14197 21437 14231 21471
rect 14231 21437 14240 21471
rect 14188 21428 14240 21437
rect 17224 21428 17276 21480
rect 18788 21428 18840 21480
rect 10968 21360 11020 21412
rect 11428 21360 11480 21412
rect 16672 21403 16724 21412
rect 16672 21369 16681 21403
rect 16681 21369 16715 21403
rect 16715 21369 16724 21403
rect 16672 21360 16724 21369
rect 28908 21428 28960 21480
rect 17040 21292 17092 21344
rect 20904 21335 20956 21344
rect 20904 21301 20913 21335
rect 20913 21301 20947 21335
rect 20947 21301 20956 21335
rect 20904 21292 20956 21301
rect 31852 21292 31904 21344
rect 34152 21641 34161 21675
rect 34161 21641 34195 21675
rect 34195 21641 34204 21675
rect 34152 21632 34204 21641
rect 43536 21632 43588 21684
rect 47768 21675 47820 21684
rect 47768 21641 47777 21675
rect 47777 21641 47811 21675
rect 47811 21641 47820 21675
rect 47768 21632 47820 21641
rect 47952 21675 48004 21684
rect 47952 21641 47961 21675
rect 47961 21641 47995 21675
rect 47995 21641 48004 21675
rect 47952 21632 48004 21641
rect 34704 21564 34756 21616
rect 42984 21564 43036 21616
rect 33784 21496 33836 21548
rect 42616 21496 42668 21548
rect 47032 21564 47084 21616
rect 47492 21564 47544 21616
rect 47860 21607 47912 21616
rect 47860 21573 47869 21607
rect 47869 21573 47903 21607
rect 47903 21573 47912 21607
rect 47860 21564 47912 21573
rect 43720 21539 43772 21548
rect 43720 21505 43729 21539
rect 43729 21505 43763 21539
rect 43763 21505 43772 21539
rect 43720 21496 43772 21505
rect 44732 21539 44784 21548
rect 44732 21505 44741 21539
rect 44741 21505 44775 21539
rect 44775 21505 44784 21539
rect 44732 21496 44784 21505
rect 47216 21496 47268 21548
rect 34520 21428 34572 21480
rect 43812 21471 43864 21480
rect 43812 21437 43821 21471
rect 43821 21437 43855 21471
rect 43855 21437 43864 21471
rect 43812 21428 43864 21437
rect 35900 21360 35952 21412
rect 42708 21360 42760 21412
rect 44640 21428 44692 21480
rect 46848 21471 46900 21480
rect 46848 21437 46857 21471
rect 46857 21437 46891 21471
rect 46891 21437 46900 21471
rect 46848 21428 46900 21437
rect 40316 21292 40368 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 3424 21088 3476 21140
rect 17040 21088 17092 21140
rect 17224 21131 17276 21140
rect 17224 21097 17233 21131
rect 17233 21097 17267 21131
rect 17267 21097 17276 21131
rect 17224 21088 17276 21097
rect 19248 21088 19300 21140
rect 23848 21131 23900 21140
rect 23848 21097 23857 21131
rect 23857 21097 23891 21131
rect 23891 21097 23900 21131
rect 23848 21088 23900 21097
rect 27344 21088 27396 21140
rect 28172 21088 28224 21140
rect 2596 21020 2648 21072
rect 25688 21020 25740 21072
rect 46756 21088 46808 21140
rect 30196 20995 30248 21004
rect 30196 20961 30205 20995
rect 30205 20961 30239 20995
rect 30239 20961 30248 20995
rect 30196 20952 30248 20961
rect 31208 20995 31260 21004
rect 31208 20961 31217 20995
rect 31217 20961 31251 20995
rect 31251 20961 31260 20995
rect 31208 20952 31260 20961
rect 46204 21020 46256 21072
rect 32128 20995 32180 21004
rect 32128 20961 32137 20995
rect 32137 20961 32171 20995
rect 32171 20961 32180 20995
rect 32128 20952 32180 20961
rect 16856 20884 16908 20936
rect 19248 20927 19300 20936
rect 19248 20893 19257 20927
rect 19257 20893 19291 20927
rect 19291 20893 19300 20927
rect 19248 20884 19300 20893
rect 20904 20884 20956 20936
rect 26700 20927 26752 20936
rect 26700 20893 26709 20927
rect 26709 20893 26743 20927
rect 26743 20893 26752 20927
rect 26700 20884 26752 20893
rect 27344 20884 27396 20936
rect 9128 20859 9180 20868
rect 9128 20825 9137 20859
rect 9137 20825 9171 20859
rect 9171 20825 9180 20859
rect 9128 20816 9180 20825
rect 10784 20859 10836 20868
rect 10784 20825 10793 20859
rect 10793 20825 10827 20859
rect 10827 20825 10836 20859
rect 10784 20816 10836 20825
rect 22652 20816 22704 20868
rect 23388 20816 23440 20868
rect 30288 20859 30340 20868
rect 30288 20825 30297 20859
rect 30297 20825 30331 20859
rect 30331 20825 30340 20859
rect 30288 20816 30340 20825
rect 31852 20859 31904 20868
rect 31852 20825 31861 20859
rect 31861 20825 31895 20859
rect 31895 20825 31904 20859
rect 31852 20816 31904 20825
rect 9772 20748 9824 20800
rect 30196 20748 30248 20800
rect 35900 20927 35952 20936
rect 35900 20893 35909 20927
rect 35909 20893 35943 20927
rect 35943 20893 35952 20927
rect 35900 20884 35952 20893
rect 33784 20816 33836 20868
rect 36360 20816 36412 20868
rect 42708 20952 42760 21004
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 42340 20884 42392 20936
rect 43904 20927 43956 20936
rect 43904 20893 43913 20927
rect 43913 20893 43947 20927
rect 43947 20893 43956 20927
rect 43904 20884 43956 20893
rect 44088 20927 44140 20936
rect 44088 20893 44097 20927
rect 44097 20893 44131 20927
rect 44131 20893 44140 20927
rect 44088 20884 44140 20893
rect 45652 20927 45704 20936
rect 45652 20893 45661 20927
rect 45661 20893 45695 20927
rect 45695 20893 45704 20927
rect 45652 20884 45704 20893
rect 43996 20791 44048 20800
rect 43996 20757 44005 20791
rect 44005 20757 44039 20791
rect 44039 20757 44048 20791
rect 43996 20748 44048 20757
rect 45928 20748 45980 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 3056 20544 3108 20596
rect 10968 20544 11020 20596
rect 12808 20476 12860 20528
rect 13820 20544 13872 20596
rect 14188 20544 14240 20596
rect 14280 20587 14332 20596
rect 14280 20553 14289 20587
rect 14289 20553 14323 20587
rect 14323 20553 14332 20587
rect 14280 20544 14332 20553
rect 19340 20544 19392 20596
rect 21272 20544 21324 20596
rect 23388 20544 23440 20596
rect 22100 20476 22152 20528
rect 11336 20408 11388 20460
rect 14004 20451 14056 20460
rect 14004 20417 14013 20451
rect 14013 20417 14047 20451
rect 14047 20417 14056 20451
rect 14004 20408 14056 20417
rect 14464 20408 14516 20460
rect 11796 20383 11848 20392
rect 11796 20349 11805 20383
rect 11805 20349 11839 20383
rect 11839 20349 11848 20383
rect 11796 20340 11848 20349
rect 13544 20340 13596 20392
rect 16856 20408 16908 20460
rect 14096 20272 14148 20324
rect 19248 20408 19300 20460
rect 13084 20204 13136 20256
rect 15660 20204 15712 20256
rect 16856 20204 16908 20256
rect 18144 20247 18196 20256
rect 18144 20213 18153 20247
rect 18153 20213 18187 20247
rect 18187 20213 18196 20247
rect 18144 20204 18196 20213
rect 18604 20204 18656 20256
rect 20812 20408 20864 20460
rect 21180 20408 21232 20460
rect 23848 20476 23900 20528
rect 22652 20340 22704 20392
rect 21732 20272 21784 20324
rect 21824 20272 21876 20324
rect 23480 20408 23532 20460
rect 24492 20408 24544 20460
rect 25780 20451 25832 20460
rect 25780 20417 25789 20451
rect 25789 20417 25823 20451
rect 25823 20417 25832 20451
rect 25780 20408 25832 20417
rect 27344 20408 27396 20460
rect 27620 20408 27672 20460
rect 30288 20476 30340 20528
rect 32312 20544 32364 20596
rect 44088 20544 44140 20596
rect 46480 20544 46532 20596
rect 48044 20587 48096 20596
rect 48044 20553 48053 20587
rect 48053 20553 48087 20587
rect 48087 20553 48096 20587
rect 48044 20544 48096 20553
rect 31208 20451 31260 20460
rect 31208 20417 31217 20451
rect 31217 20417 31251 20451
rect 31251 20417 31260 20451
rect 31208 20408 31260 20417
rect 45560 20476 45612 20528
rect 42340 20408 42392 20460
rect 42708 20408 42760 20460
rect 43352 20408 43404 20460
rect 43996 20408 44048 20460
rect 44640 20451 44692 20460
rect 44640 20417 44649 20451
rect 44649 20417 44683 20451
rect 44683 20417 44692 20451
rect 44640 20408 44692 20417
rect 47952 20408 48004 20460
rect 29920 20340 29972 20392
rect 30012 20383 30064 20392
rect 30012 20349 30021 20383
rect 30021 20349 30055 20383
rect 30055 20349 30064 20383
rect 30012 20340 30064 20349
rect 41052 20340 41104 20392
rect 43536 20383 43588 20392
rect 43536 20349 43545 20383
rect 43545 20349 43579 20383
rect 43579 20349 43588 20383
rect 43536 20340 43588 20349
rect 45192 20340 45244 20392
rect 46020 20383 46072 20392
rect 46020 20349 46029 20383
rect 46029 20349 46063 20383
rect 46063 20349 46072 20383
rect 46020 20340 46072 20349
rect 24584 20272 24636 20324
rect 27160 20272 27212 20324
rect 20260 20247 20312 20256
rect 20260 20213 20269 20247
rect 20269 20213 20303 20247
rect 20303 20213 20312 20247
rect 20260 20204 20312 20213
rect 25228 20204 25280 20256
rect 25504 20204 25556 20256
rect 26240 20204 26292 20256
rect 27068 20247 27120 20256
rect 27068 20213 27077 20247
rect 27077 20213 27111 20247
rect 27111 20213 27120 20247
rect 27068 20204 27120 20213
rect 30196 20204 30248 20256
rect 32312 20247 32364 20256
rect 32312 20213 32321 20247
rect 32321 20213 32355 20247
rect 32355 20213 32364 20247
rect 32312 20204 32364 20213
rect 47216 20204 47268 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3516 20000 3568 20052
rect 30012 20000 30064 20052
rect 45192 20043 45244 20052
rect 45192 20009 45201 20043
rect 45201 20009 45235 20043
rect 45235 20009 45244 20043
rect 45192 20000 45244 20009
rect 11796 19932 11848 19984
rect 12808 19975 12860 19984
rect 12808 19941 12817 19975
rect 12817 19941 12851 19975
rect 12851 19941 12860 19975
rect 12808 19932 12860 19941
rect 21732 19975 21784 19984
rect 21732 19941 21741 19975
rect 21741 19941 21775 19975
rect 21775 19941 21784 19975
rect 21732 19932 21784 19941
rect 43812 19975 43864 19984
rect 43812 19941 43821 19975
rect 43821 19941 43855 19975
rect 43855 19941 43864 19975
rect 43812 19932 43864 19941
rect 10968 19864 11020 19916
rect 11888 19796 11940 19848
rect 12348 19864 12400 19916
rect 16856 19907 16908 19916
rect 13084 19796 13136 19848
rect 16856 19873 16865 19907
rect 16865 19873 16899 19907
rect 16899 19873 16908 19907
rect 16856 19864 16908 19873
rect 18328 19864 18380 19916
rect 19432 19864 19484 19916
rect 20996 19864 21048 19916
rect 25228 19907 25280 19916
rect 25228 19873 25237 19907
rect 25237 19873 25271 19907
rect 25271 19873 25280 19907
rect 25228 19864 25280 19873
rect 25504 19907 25556 19916
rect 25504 19873 25513 19907
rect 25513 19873 25547 19907
rect 25547 19873 25556 19907
rect 25504 19864 25556 19873
rect 30196 19907 30248 19916
rect 30196 19873 30205 19907
rect 30205 19873 30239 19907
rect 30239 19873 30248 19907
rect 30196 19864 30248 19873
rect 31668 19907 31720 19916
rect 31668 19873 31677 19907
rect 31677 19873 31711 19907
rect 31711 19873 31720 19907
rect 31668 19864 31720 19873
rect 43352 19907 43404 19916
rect 43352 19873 43361 19907
rect 43361 19873 43395 19907
rect 43395 19873 43404 19907
rect 43352 19864 43404 19873
rect 43904 19907 43956 19916
rect 43904 19873 43913 19907
rect 43913 19873 43947 19907
rect 43947 19873 43956 19907
rect 43904 19864 43956 19873
rect 46480 19932 46532 19984
rect 46388 19907 46440 19916
rect 46388 19873 46397 19907
rect 46397 19873 46431 19907
rect 46431 19873 46440 19907
rect 46388 19864 46440 19873
rect 46848 19864 46900 19916
rect 19984 19839 20036 19848
rect 19984 19805 19993 19839
rect 19993 19805 20027 19839
rect 20027 19805 20036 19839
rect 19984 19796 20036 19805
rect 24492 19839 24544 19848
rect 24492 19805 24501 19839
rect 24501 19805 24535 19839
rect 24535 19805 24544 19839
rect 24492 19796 24544 19805
rect 27160 19796 27212 19848
rect 42432 19796 42484 19848
rect 44824 19796 44876 19848
rect 45836 19796 45888 19848
rect 13728 19728 13780 19780
rect 14096 19728 14148 19780
rect 15752 19728 15804 19780
rect 18144 19728 18196 19780
rect 20536 19728 20588 19780
rect 21916 19728 21968 19780
rect 25412 19728 25464 19780
rect 26240 19728 26292 19780
rect 43904 19728 43956 19780
rect 14004 19660 14056 19712
rect 14832 19660 14884 19712
rect 16304 19660 16356 19712
rect 18604 19703 18656 19712
rect 18604 19669 18613 19703
rect 18613 19669 18647 19703
rect 18647 19669 18656 19703
rect 18604 19660 18656 19669
rect 19248 19660 19300 19712
rect 21824 19660 21876 19712
rect 23296 19660 23348 19712
rect 35992 19660 36044 19712
rect 45928 19660 45980 19712
rect 47676 19660 47728 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1676 19456 1728 19508
rect 3056 19388 3108 19440
rect 13820 19431 13872 19440
rect 13820 19397 13829 19431
rect 13829 19397 13863 19431
rect 13863 19397 13872 19431
rect 13820 19388 13872 19397
rect 14004 19431 14056 19440
rect 14004 19397 14013 19431
rect 14013 19397 14047 19431
rect 14047 19397 14056 19431
rect 14004 19388 14056 19397
rect 14464 19388 14516 19440
rect 14832 19431 14884 19440
rect 14832 19397 14841 19431
rect 14841 19397 14875 19431
rect 14875 19397 14884 19431
rect 14832 19388 14884 19397
rect 15016 19431 15068 19440
rect 15016 19397 15041 19431
rect 15041 19397 15068 19431
rect 15752 19431 15804 19440
rect 15016 19388 15068 19397
rect 15752 19397 15761 19431
rect 15761 19397 15795 19431
rect 15795 19397 15804 19431
rect 15752 19388 15804 19397
rect 18512 19388 18564 19440
rect 19064 19388 19116 19440
rect 19984 19388 20036 19440
rect 11336 19320 11388 19372
rect 12348 19320 12400 19372
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 16580 19320 16632 19372
rect 18604 19320 18656 19372
rect 19432 19363 19484 19372
rect 19432 19329 19441 19363
rect 19441 19329 19475 19363
rect 19475 19329 19484 19363
rect 19432 19320 19484 19329
rect 21732 19388 21784 19440
rect 21916 19431 21968 19440
rect 21916 19397 21925 19431
rect 21925 19397 21959 19431
rect 21959 19397 21968 19431
rect 21916 19388 21968 19397
rect 25780 19456 25832 19508
rect 28264 19456 28316 19508
rect 28724 19456 28776 19508
rect 29920 19499 29972 19508
rect 29920 19465 29929 19499
rect 29929 19465 29963 19499
rect 29963 19465 29972 19499
rect 29920 19456 29972 19465
rect 43536 19499 43588 19508
rect 43536 19465 43545 19499
rect 43545 19465 43579 19499
rect 43579 19465 43588 19499
rect 43536 19456 43588 19465
rect 45560 19388 45612 19440
rect 21180 19363 21232 19372
rect 2044 19295 2096 19304
rect 2044 19261 2053 19295
rect 2053 19261 2087 19295
rect 2087 19261 2096 19295
rect 2044 19252 2096 19261
rect 2780 19295 2832 19304
rect 2780 19261 2789 19295
rect 2789 19261 2823 19295
rect 2823 19261 2832 19295
rect 2780 19252 2832 19261
rect 14280 19252 14332 19304
rect 18328 19295 18380 19304
rect 18328 19261 18337 19295
rect 18337 19261 18371 19295
rect 18371 19261 18380 19295
rect 18328 19252 18380 19261
rect 20260 19295 20312 19304
rect 20260 19261 20269 19295
rect 20269 19261 20303 19295
rect 20303 19261 20312 19295
rect 20260 19252 20312 19261
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 21180 19329 21189 19363
rect 21189 19329 21223 19363
rect 21223 19329 21232 19363
rect 21180 19320 21232 19329
rect 21272 19363 21324 19372
rect 21272 19329 21281 19363
rect 21281 19329 21315 19363
rect 21315 19329 21324 19363
rect 21824 19363 21876 19372
rect 21272 19320 21324 19329
rect 21824 19329 21833 19363
rect 21833 19329 21867 19363
rect 21867 19329 21876 19363
rect 21824 19320 21876 19329
rect 23756 19363 23808 19372
rect 23756 19329 23765 19363
rect 23765 19329 23799 19363
rect 23799 19329 23808 19363
rect 23756 19320 23808 19329
rect 24584 19363 24636 19372
rect 24584 19329 24593 19363
rect 24593 19329 24627 19363
rect 24627 19329 24636 19363
rect 24584 19320 24636 19329
rect 25596 19363 25648 19372
rect 22100 19252 22152 19304
rect 22560 19252 22612 19304
rect 25044 19252 25096 19304
rect 19340 19184 19392 19236
rect 24400 19184 24452 19236
rect 25596 19329 25605 19363
rect 25605 19329 25639 19363
rect 25639 19329 25648 19363
rect 25596 19320 25648 19329
rect 28264 19363 28316 19372
rect 28264 19329 28273 19363
rect 28273 19329 28307 19363
rect 28307 19329 28316 19363
rect 28264 19320 28316 19329
rect 28908 19320 28960 19372
rect 42432 19320 42484 19372
rect 43904 19320 43956 19372
rect 45928 19363 45980 19372
rect 45928 19329 45937 19363
rect 45937 19329 45971 19363
rect 45971 19329 45980 19363
rect 45928 19320 45980 19329
rect 47952 19456 48004 19508
rect 48044 19456 48096 19508
rect 29092 19295 29144 19304
rect 29092 19261 29101 19295
rect 29101 19261 29135 19295
rect 29135 19261 29144 19295
rect 29092 19252 29144 19261
rect 47676 19320 47728 19372
rect 47860 19184 47912 19236
rect 11796 19116 11848 19168
rect 12072 19116 12124 19168
rect 13728 19116 13780 19168
rect 14464 19116 14516 19168
rect 15108 19116 15160 19168
rect 20720 19116 20772 19168
rect 22376 19116 22428 19168
rect 24860 19159 24912 19168
rect 24860 19125 24869 19159
rect 24869 19125 24903 19159
rect 24903 19125 24912 19159
rect 24860 19116 24912 19125
rect 25044 19116 25096 19168
rect 45468 19159 45520 19168
rect 45468 19125 45477 19159
rect 45477 19125 45511 19159
rect 45511 19125 45520 19159
rect 45468 19116 45520 19125
rect 46204 19159 46256 19168
rect 46204 19125 46213 19159
rect 46213 19125 46247 19159
rect 46247 19125 46256 19159
rect 46204 19116 46256 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2044 18912 2096 18964
rect 3056 18955 3108 18964
rect 3056 18921 3065 18955
rect 3065 18921 3099 18955
rect 3099 18921 3108 18955
rect 3056 18912 3108 18921
rect 13820 18912 13872 18964
rect 14096 18955 14148 18964
rect 14096 18921 14105 18955
rect 14105 18921 14139 18955
rect 14139 18921 14148 18955
rect 14096 18912 14148 18921
rect 13728 18844 13780 18896
rect 36268 18912 36320 18964
rect 11796 18819 11848 18828
rect 11796 18785 11805 18819
rect 11805 18785 11839 18819
rect 11839 18785 11848 18819
rect 11796 18776 11848 18785
rect 12072 18819 12124 18828
rect 12072 18785 12081 18819
rect 12081 18785 12115 18819
rect 12115 18785 12124 18819
rect 12072 18776 12124 18785
rect 2964 18751 3016 18760
rect 2964 18717 2973 18751
rect 2973 18717 3007 18751
rect 3007 18717 3016 18751
rect 2964 18708 3016 18717
rect 13176 18708 13228 18760
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 14832 18708 14884 18760
rect 15016 18751 15068 18760
rect 15016 18717 15025 18751
rect 15025 18717 15059 18751
rect 15059 18717 15068 18751
rect 15016 18708 15068 18717
rect 16580 18708 16632 18760
rect 20720 18844 20772 18896
rect 23756 18844 23808 18896
rect 27160 18887 27212 18896
rect 27160 18853 27169 18887
rect 27169 18853 27203 18887
rect 27203 18853 27212 18887
rect 27160 18844 27212 18853
rect 20260 18776 20312 18828
rect 24860 18776 24912 18828
rect 27804 18776 27856 18828
rect 20812 18751 20864 18760
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 24400 18751 24452 18760
rect 24400 18717 24409 18751
rect 24409 18717 24443 18751
rect 24443 18717 24452 18751
rect 24400 18708 24452 18717
rect 24768 18708 24820 18760
rect 25412 18751 25464 18760
rect 25412 18717 25421 18751
rect 25421 18717 25455 18751
rect 25455 18717 25464 18751
rect 25412 18708 25464 18717
rect 29092 18844 29144 18896
rect 29920 18776 29972 18828
rect 28724 18708 28776 18760
rect 29000 18751 29052 18760
rect 29000 18717 29009 18751
rect 29009 18717 29043 18751
rect 29043 18717 29052 18751
rect 29000 18708 29052 18717
rect 43260 18708 43312 18760
rect 43904 18751 43956 18760
rect 22376 18640 22428 18692
rect 27068 18640 27120 18692
rect 30012 18640 30064 18692
rect 30288 18640 30340 18692
rect 31116 18640 31168 18692
rect 31944 18640 31996 18692
rect 32128 18683 32180 18692
rect 32128 18649 32137 18683
rect 32137 18649 32171 18683
rect 32171 18649 32180 18683
rect 32128 18640 32180 18649
rect 42064 18640 42116 18692
rect 43904 18717 43913 18751
rect 43913 18717 43947 18751
rect 43947 18717 43956 18751
rect 43904 18708 43956 18717
rect 44916 18708 44968 18760
rect 45468 18776 45520 18828
rect 48136 18819 48188 18828
rect 48136 18785 48145 18819
rect 48145 18785 48179 18819
rect 48179 18785 48188 18819
rect 48136 18776 48188 18785
rect 45100 18708 45152 18760
rect 45836 18751 45888 18760
rect 45836 18717 45845 18751
rect 45845 18717 45879 18751
rect 45879 18717 45888 18751
rect 45836 18708 45888 18717
rect 15108 18572 15160 18624
rect 17316 18615 17368 18624
rect 17316 18581 17325 18615
rect 17325 18581 17359 18615
rect 17359 18581 17368 18615
rect 17316 18572 17368 18581
rect 22560 18615 22612 18624
rect 22560 18581 22569 18615
rect 22569 18581 22603 18615
rect 22603 18581 22612 18615
rect 22560 18572 22612 18581
rect 23112 18572 23164 18624
rect 28172 18572 28224 18624
rect 30196 18572 30248 18624
rect 43812 18615 43864 18624
rect 43812 18581 43821 18615
rect 43821 18581 43855 18615
rect 43855 18581 43864 18615
rect 43812 18572 43864 18581
rect 47676 18640 47728 18692
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2964 18368 3016 18420
rect 12992 18368 13044 18420
rect 13176 18411 13228 18420
rect 13176 18377 13185 18411
rect 13185 18377 13219 18411
rect 13219 18377 13228 18411
rect 13176 18368 13228 18377
rect 20812 18368 20864 18420
rect 24492 18368 24544 18420
rect 29736 18368 29788 18420
rect 47676 18411 47728 18420
rect 47676 18377 47685 18411
rect 47685 18377 47719 18411
rect 47719 18377 47728 18411
rect 47676 18368 47728 18377
rect 4620 18300 4672 18352
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 16304 18232 16356 18284
rect 20996 18232 21048 18284
rect 22192 18232 22244 18284
rect 23296 18275 23348 18284
rect 23296 18241 23305 18275
rect 23305 18241 23339 18275
rect 23339 18241 23348 18275
rect 23296 18232 23348 18241
rect 24860 18232 24912 18284
rect 27528 18275 27580 18284
rect 27528 18241 27537 18275
rect 27537 18241 27571 18275
rect 27571 18241 27580 18275
rect 27528 18232 27580 18241
rect 28172 18275 28224 18284
rect 28172 18241 28181 18275
rect 28181 18241 28215 18275
rect 28215 18241 28224 18275
rect 28172 18232 28224 18241
rect 31116 18275 31168 18284
rect 12992 18164 13044 18216
rect 13728 18164 13780 18216
rect 17132 18207 17184 18216
rect 17132 18173 17141 18207
rect 17141 18173 17175 18207
rect 17175 18173 17184 18207
rect 17132 18164 17184 18173
rect 18788 18207 18840 18216
rect 18788 18173 18797 18207
rect 18797 18173 18831 18207
rect 18831 18173 18840 18207
rect 18788 18164 18840 18173
rect 23480 18164 23532 18216
rect 24676 18164 24728 18216
rect 31116 18241 31125 18275
rect 31125 18241 31159 18275
rect 31159 18241 31168 18275
rect 31116 18232 31168 18241
rect 40132 18232 40184 18284
rect 40776 18275 40828 18284
rect 40776 18241 40785 18275
rect 40785 18241 40819 18275
rect 40819 18241 40828 18275
rect 40776 18232 40828 18241
rect 42524 18232 42576 18284
rect 46204 18300 46256 18352
rect 43812 18275 43864 18284
rect 43812 18241 43821 18275
rect 43821 18241 43855 18275
rect 43855 18241 43864 18275
rect 43812 18232 43864 18241
rect 47032 18232 47084 18284
rect 47400 18232 47452 18284
rect 3332 18096 3384 18148
rect 24492 18028 24544 18080
rect 24768 18028 24820 18080
rect 42156 18164 42208 18216
rect 45008 18164 45060 18216
rect 46848 18207 46900 18216
rect 46848 18173 46857 18207
rect 46857 18173 46891 18207
rect 46891 18173 46900 18207
rect 46848 18164 46900 18173
rect 30380 18028 30432 18080
rect 40040 18096 40092 18148
rect 42064 18096 42116 18148
rect 44180 18096 44232 18148
rect 40960 18028 41012 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 17132 17824 17184 17876
rect 23572 17824 23624 17876
rect 23756 17824 23808 17876
rect 14832 17756 14884 17808
rect 22744 17756 22796 17808
rect 24584 17756 24636 17808
rect 42524 17824 42576 17876
rect 42708 17824 42760 17876
rect 43904 17824 43956 17876
rect 14648 17731 14700 17740
rect 14648 17697 14657 17731
rect 14657 17697 14691 17731
rect 14691 17697 14700 17731
rect 14648 17688 14700 17697
rect 23388 17688 23440 17740
rect 24676 17731 24728 17740
rect 24676 17697 24685 17731
rect 24685 17697 24719 17731
rect 24719 17697 24728 17731
rect 24676 17688 24728 17697
rect 42156 17756 42208 17808
rect 42432 17799 42484 17808
rect 42432 17765 42441 17799
rect 42441 17765 42475 17799
rect 42475 17765 42484 17799
rect 42432 17756 42484 17765
rect 1768 17620 1820 17672
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 14832 17663 14884 17672
rect 14832 17629 14841 17663
rect 14841 17629 14875 17663
rect 14875 17629 14884 17663
rect 14832 17620 14884 17629
rect 17316 17620 17368 17672
rect 18512 17663 18564 17672
rect 18512 17629 18521 17663
rect 18521 17629 18555 17663
rect 18555 17629 18564 17663
rect 18512 17620 18564 17629
rect 19156 17620 19208 17672
rect 20996 17620 21048 17672
rect 23480 17620 23532 17672
rect 24400 17620 24452 17672
rect 3516 17552 3568 17604
rect 9036 17552 9088 17604
rect 21088 17595 21140 17604
rect 21088 17561 21097 17595
rect 21097 17561 21131 17595
rect 21131 17561 21140 17595
rect 21088 17552 21140 17561
rect 23296 17595 23348 17604
rect 23296 17561 23305 17595
rect 23305 17561 23339 17595
rect 23339 17561 23348 17595
rect 23296 17552 23348 17561
rect 25136 17620 25188 17672
rect 26700 17620 26752 17672
rect 27804 17663 27856 17672
rect 27804 17629 27813 17663
rect 27813 17629 27847 17663
rect 27847 17629 27856 17663
rect 27804 17620 27856 17629
rect 28724 17688 28776 17740
rect 30196 17731 30248 17740
rect 30196 17697 30205 17731
rect 30205 17697 30239 17731
rect 30239 17697 30248 17731
rect 30196 17688 30248 17697
rect 30380 17731 30432 17740
rect 30380 17697 30389 17731
rect 30389 17697 30423 17731
rect 30423 17697 30432 17731
rect 30380 17688 30432 17697
rect 32128 17688 32180 17740
rect 40960 17731 41012 17740
rect 40960 17697 40969 17731
rect 40969 17697 41003 17731
rect 41003 17697 41012 17731
rect 40960 17688 41012 17697
rect 28632 17663 28684 17672
rect 28632 17629 28641 17663
rect 28641 17629 28675 17663
rect 28675 17629 28684 17663
rect 28632 17620 28684 17629
rect 42156 17663 42208 17672
rect 1952 17484 2004 17536
rect 15016 17527 15068 17536
rect 15016 17493 15025 17527
rect 15025 17493 15059 17527
rect 15059 17493 15068 17527
rect 15016 17484 15068 17493
rect 29000 17552 29052 17604
rect 42156 17629 42165 17663
rect 42165 17629 42199 17663
rect 42199 17629 42208 17663
rect 42156 17620 42208 17629
rect 43260 17620 43312 17672
rect 45560 17756 45612 17808
rect 43444 17663 43496 17672
rect 43444 17629 43453 17663
rect 43453 17629 43487 17663
rect 43487 17629 43496 17663
rect 47952 17688 48004 17740
rect 43444 17620 43496 17629
rect 42708 17595 42760 17604
rect 42708 17561 42717 17595
rect 42717 17561 42751 17595
rect 42751 17561 42760 17595
rect 42708 17552 42760 17561
rect 43168 17552 43220 17604
rect 44916 17620 44968 17672
rect 46296 17663 46348 17672
rect 46296 17629 46305 17663
rect 46305 17629 46339 17663
rect 46339 17629 46348 17663
rect 46296 17620 46348 17629
rect 43720 17552 43772 17604
rect 45100 17552 45152 17604
rect 47676 17552 47728 17604
rect 48136 17595 48188 17604
rect 48136 17561 48145 17595
rect 48145 17561 48179 17595
rect 48179 17561 48188 17595
rect 48136 17552 48188 17561
rect 23664 17484 23716 17536
rect 23848 17527 23900 17536
rect 23848 17493 23857 17527
rect 23857 17493 23891 17527
rect 23891 17493 23900 17527
rect 23848 17484 23900 17493
rect 24676 17484 24728 17536
rect 25596 17527 25648 17536
rect 25596 17493 25605 17527
rect 25605 17493 25639 17527
rect 25639 17493 25648 17527
rect 25596 17484 25648 17493
rect 42524 17484 42576 17536
rect 43444 17484 43496 17536
rect 47860 17484 47912 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 2136 17280 2188 17332
rect 37648 17280 37700 17332
rect 40040 17280 40092 17332
rect 43444 17280 43496 17332
rect 47676 17323 47728 17332
rect 1952 17255 2004 17264
rect 1952 17221 1961 17255
rect 1961 17221 1995 17255
rect 1995 17221 2004 17255
rect 1952 17212 2004 17221
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 15660 17144 15712 17196
rect 20996 17212 21048 17264
rect 22192 17212 22244 17264
rect 22744 17255 22796 17264
rect 22744 17221 22753 17255
rect 22753 17221 22787 17255
rect 22787 17221 22796 17255
rect 22744 17212 22796 17221
rect 23388 17212 23440 17264
rect 24768 17255 24820 17264
rect 24768 17221 24777 17255
rect 24777 17221 24811 17255
rect 24811 17221 24820 17255
rect 24768 17212 24820 17221
rect 25504 17212 25556 17264
rect 27804 17255 27856 17264
rect 27804 17221 27813 17255
rect 27813 17221 27847 17255
rect 27847 17221 27856 17255
rect 27804 17212 27856 17221
rect 40132 17212 40184 17264
rect 43168 17212 43220 17264
rect 14924 17076 14976 17128
rect 22468 17187 22520 17196
rect 22468 17153 22477 17187
rect 22477 17153 22511 17187
rect 22511 17153 22520 17187
rect 22468 17144 22520 17153
rect 23480 17187 23532 17196
rect 20996 17076 21048 17128
rect 23480 17153 23489 17187
rect 23489 17153 23523 17187
rect 23523 17153 23532 17187
rect 23480 17144 23532 17153
rect 26884 17144 26936 17196
rect 27160 17144 27212 17196
rect 42708 17144 42760 17196
rect 43720 17255 43772 17264
rect 43720 17221 43729 17255
rect 43729 17221 43763 17255
rect 43763 17221 43772 17255
rect 43720 17212 43772 17221
rect 24492 17119 24544 17128
rect 20444 17051 20496 17060
rect 20444 17017 20453 17051
rect 20453 17017 20487 17051
rect 20487 17017 20496 17051
rect 20444 17008 20496 17017
rect 21824 17008 21876 17060
rect 14372 16940 14424 16992
rect 15384 16940 15436 16992
rect 17960 16940 18012 16992
rect 22468 17008 22520 17060
rect 24492 17085 24501 17119
rect 24501 17085 24535 17119
rect 24535 17085 24544 17119
rect 24492 17076 24544 17085
rect 23296 17051 23348 17060
rect 23296 17017 23305 17051
rect 23305 17017 23339 17051
rect 23339 17017 23348 17051
rect 25136 17076 25188 17128
rect 29460 17119 29512 17128
rect 23296 17008 23348 17017
rect 25780 17008 25832 17060
rect 29460 17085 29469 17119
rect 29469 17085 29503 17119
rect 29503 17085 29512 17119
rect 29460 17076 29512 17085
rect 31116 17119 31168 17128
rect 31116 17085 31125 17119
rect 31125 17085 31159 17119
rect 31159 17085 31168 17119
rect 31116 17076 31168 17085
rect 42524 17119 42576 17128
rect 42524 17085 42533 17119
rect 42533 17085 42567 17119
rect 42567 17085 42576 17119
rect 42524 17076 42576 17085
rect 40684 17008 40736 17060
rect 46296 17144 46348 17196
rect 47676 17289 47685 17323
rect 47685 17289 47719 17323
rect 47719 17289 47728 17323
rect 47676 17280 47728 17289
rect 43904 17076 43956 17128
rect 44180 17119 44232 17128
rect 44180 17085 44189 17119
rect 44189 17085 44223 17119
rect 44223 17085 44232 17119
rect 44180 17076 44232 17085
rect 46756 17076 46808 17128
rect 44272 17008 44324 17060
rect 47584 17008 47636 17060
rect 23480 16940 23532 16992
rect 46940 16983 46992 16992
rect 46940 16949 46949 16983
rect 46949 16949 46983 16983
rect 46983 16949 46992 16983
rect 46940 16940 46992 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 22560 16736 22612 16788
rect 23112 16736 23164 16788
rect 25780 16736 25832 16788
rect 28632 16736 28684 16788
rect 29460 16736 29512 16788
rect 14372 16643 14424 16652
rect 14372 16609 14381 16643
rect 14381 16609 14415 16643
rect 14415 16609 14424 16643
rect 14372 16600 14424 16609
rect 15660 16600 15712 16652
rect 17592 16643 17644 16652
rect 17592 16609 17601 16643
rect 17601 16609 17635 16643
rect 17635 16609 17644 16643
rect 17592 16600 17644 16609
rect 18236 16600 18288 16652
rect 19984 16600 20036 16652
rect 22468 16668 22520 16720
rect 24676 16711 24728 16720
rect 18144 16532 18196 16584
rect 23848 16600 23900 16652
rect 24676 16677 24685 16711
rect 24685 16677 24719 16711
rect 24719 16677 24728 16711
rect 24676 16668 24728 16677
rect 25228 16600 25280 16652
rect 25596 16600 25648 16652
rect 26884 16643 26936 16652
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 14648 16507 14700 16516
rect 14648 16473 14657 16507
rect 14657 16473 14691 16507
rect 14691 16473 14700 16507
rect 14648 16464 14700 16473
rect 15384 16464 15436 16516
rect 16580 16464 16632 16516
rect 18788 16464 18840 16516
rect 22100 16464 22152 16516
rect 23664 16464 23716 16516
rect 25504 16575 25556 16584
rect 25504 16541 25513 16575
rect 25513 16541 25547 16575
rect 25547 16541 25556 16575
rect 27160 16600 27212 16652
rect 29276 16600 29328 16652
rect 44916 16600 44968 16652
rect 25504 16532 25556 16541
rect 29552 16575 29604 16584
rect 29552 16541 29561 16575
rect 29561 16541 29595 16575
rect 29595 16541 29604 16575
rect 29552 16532 29604 16541
rect 47768 16600 47820 16652
rect 46296 16464 46348 16516
rect 46940 16464 46992 16516
rect 48136 16507 48188 16516
rect 48136 16473 48145 16507
rect 48145 16473 48179 16507
rect 48179 16473 48188 16507
rect 48136 16464 48188 16473
rect 16948 16439 17000 16448
rect 16948 16405 16957 16439
rect 16957 16405 16991 16439
rect 16991 16405 17000 16439
rect 16948 16396 17000 16405
rect 19340 16396 19392 16448
rect 21916 16439 21968 16448
rect 21916 16405 21925 16439
rect 21925 16405 21959 16439
rect 21959 16405 21968 16439
rect 21916 16396 21968 16405
rect 24860 16439 24912 16448
rect 24860 16405 24869 16439
rect 24869 16405 24903 16439
rect 24903 16405 24912 16439
rect 24860 16396 24912 16405
rect 45192 16396 45244 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 15108 16192 15160 16244
rect 16580 16192 16632 16244
rect 20996 16192 21048 16244
rect 24492 16192 24544 16244
rect 15016 16124 15068 16176
rect 14924 16099 14976 16108
rect 14924 16065 14933 16099
rect 14933 16065 14967 16099
rect 14967 16065 14976 16099
rect 14924 16056 14976 16065
rect 14648 15988 14700 16040
rect 16028 16056 16080 16108
rect 17868 16124 17920 16176
rect 18236 16167 18288 16176
rect 18236 16133 18245 16167
rect 18245 16133 18279 16167
rect 18279 16133 18288 16167
rect 18236 16124 18288 16133
rect 17960 16099 18012 16108
rect 17960 16065 17969 16099
rect 17969 16065 18003 16099
rect 18003 16065 18012 16099
rect 17960 16056 18012 16065
rect 19340 16056 19392 16108
rect 19800 16056 19852 16108
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 22100 16056 22152 16108
rect 22560 16099 22612 16108
rect 22560 16065 22569 16099
rect 22569 16065 22603 16099
rect 22603 16065 22612 16099
rect 22560 16056 22612 16065
rect 23848 16124 23900 16176
rect 17776 15988 17828 16040
rect 23480 16056 23532 16108
rect 23756 16099 23808 16108
rect 23756 16065 23765 16099
rect 23765 16065 23799 16099
rect 23799 16065 23808 16099
rect 23756 16056 23808 16065
rect 43904 16099 43956 16108
rect 43904 16065 43913 16099
rect 43913 16065 43947 16099
rect 43947 16065 43956 16099
rect 43904 16056 43956 16065
rect 47768 16099 47820 16108
rect 47768 16065 47777 16099
rect 47777 16065 47811 16099
rect 47811 16065 47820 16099
rect 47768 16056 47820 16065
rect 44088 16031 44140 16040
rect 44088 15997 44097 16031
rect 44097 15997 44131 16031
rect 44131 15997 44140 16031
rect 44088 15988 44140 15997
rect 45468 16031 45520 16040
rect 45468 15997 45477 16031
rect 45477 15997 45511 16031
rect 45511 15997 45520 16031
rect 45468 15988 45520 15997
rect 14924 15895 14976 15904
rect 14924 15861 14933 15895
rect 14933 15861 14967 15895
rect 14967 15861 14976 15895
rect 14924 15852 14976 15861
rect 15200 15852 15252 15904
rect 17960 15852 18012 15904
rect 18604 15852 18656 15904
rect 20904 15852 20956 15904
rect 23112 15895 23164 15904
rect 23112 15861 23121 15895
rect 23121 15861 23155 15895
rect 23155 15861 23164 15895
rect 23112 15852 23164 15861
rect 24400 15852 24452 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 17776 15691 17828 15700
rect 17776 15657 17785 15691
rect 17785 15657 17819 15691
rect 17819 15657 17828 15691
rect 17776 15648 17828 15657
rect 18144 15580 18196 15632
rect 14924 15555 14976 15564
rect 14924 15521 14933 15555
rect 14933 15521 14967 15555
rect 14967 15521 14976 15555
rect 14924 15512 14976 15521
rect 15200 15555 15252 15564
rect 15200 15521 15209 15555
rect 15209 15521 15243 15555
rect 15243 15521 15252 15555
rect 15200 15512 15252 15521
rect 1768 15444 1820 15496
rect 16948 15444 17000 15496
rect 18604 15487 18656 15496
rect 17960 15376 18012 15428
rect 18604 15453 18613 15487
rect 18613 15453 18647 15487
rect 18647 15453 18656 15487
rect 18604 15444 18656 15453
rect 23480 15648 23532 15700
rect 44088 15691 44140 15700
rect 44088 15657 44097 15691
rect 44097 15657 44131 15691
rect 44131 15657 44140 15691
rect 44088 15648 44140 15657
rect 20904 15555 20956 15564
rect 20904 15521 20913 15555
rect 20913 15521 20947 15555
rect 20947 15521 20956 15555
rect 20904 15512 20956 15521
rect 23112 15512 23164 15564
rect 23756 15512 23808 15564
rect 19800 15444 19852 15496
rect 19984 15487 20036 15496
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 22560 15444 22612 15496
rect 24400 15487 24452 15496
rect 15936 15308 15988 15360
rect 17592 15351 17644 15360
rect 17592 15317 17627 15351
rect 17627 15317 17644 15351
rect 21916 15376 21968 15428
rect 17592 15308 17644 15317
rect 18144 15308 18196 15360
rect 19432 15351 19484 15360
rect 19432 15317 19441 15351
rect 19441 15317 19475 15351
rect 19475 15317 19484 15351
rect 19432 15308 19484 15317
rect 20168 15308 20220 15360
rect 22100 15308 22152 15360
rect 24400 15453 24409 15487
rect 24409 15453 24443 15487
rect 24443 15453 24452 15487
rect 24400 15444 24452 15453
rect 40868 15444 40920 15496
rect 47308 15580 47360 15632
rect 45008 15555 45060 15564
rect 45008 15521 45017 15555
rect 45017 15521 45051 15555
rect 45051 15521 45060 15555
rect 45008 15512 45060 15521
rect 45192 15555 45244 15564
rect 45192 15521 45201 15555
rect 45201 15521 45235 15555
rect 45235 15521 45244 15555
rect 45192 15512 45244 15521
rect 46664 15555 46716 15564
rect 46664 15521 46673 15555
rect 46673 15521 46707 15555
rect 46707 15521 46716 15555
rect 46664 15512 46716 15521
rect 25320 15376 25372 15428
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 25320 15147 25372 15156
rect 25320 15113 25329 15147
rect 25329 15113 25363 15147
rect 25363 15113 25372 15147
rect 25320 15104 25372 15113
rect 20168 15036 20220 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 16764 14968 16816 15020
rect 17316 14968 17368 15020
rect 17960 14968 18012 15020
rect 25228 15011 25280 15020
rect 25228 14977 25237 15011
rect 25237 14977 25271 15011
rect 25271 14977 25280 15011
rect 25228 14968 25280 14977
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 18144 14943 18196 14952
rect 18144 14909 18153 14943
rect 18153 14909 18187 14943
rect 18187 14909 18196 14943
rect 18144 14900 18196 14909
rect 19524 14900 19576 14952
rect 22100 14943 22152 14952
rect 22100 14909 22109 14943
rect 22109 14909 22143 14943
rect 22143 14909 22152 14943
rect 22284 14943 22336 14952
rect 22100 14900 22152 14909
rect 22284 14909 22293 14943
rect 22293 14909 22327 14943
rect 22327 14909 22336 14943
rect 22284 14900 22336 14909
rect 23940 14943 23992 14952
rect 23940 14909 23949 14943
rect 23949 14909 23983 14943
rect 23983 14909 23992 14943
rect 23940 14900 23992 14909
rect 16120 14764 16172 14816
rect 17960 14764 18012 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 27528 14560 27580 14612
rect 2136 14356 2188 14365
rect 3332 14220 3384 14272
rect 15936 14467 15988 14476
rect 15936 14433 15945 14467
rect 15945 14433 15979 14467
rect 15979 14433 15988 14467
rect 15936 14424 15988 14433
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 22284 14492 22336 14544
rect 31208 14492 31260 14544
rect 22468 14424 22520 14476
rect 23572 14467 23624 14476
rect 23572 14433 23581 14467
rect 23581 14433 23615 14467
rect 23615 14433 23624 14467
rect 23572 14424 23624 14433
rect 22008 14220 22060 14272
rect 22192 14331 22244 14340
rect 22192 14297 22201 14331
rect 22201 14297 22235 14331
rect 22235 14297 22244 14331
rect 22192 14288 22244 14297
rect 22560 14220 22612 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 22008 13991 22060 14000
rect 22008 13957 22017 13991
rect 22017 13957 22051 13991
rect 22051 13957 22060 13991
rect 22008 13948 22060 13957
rect 16764 13923 16816 13932
rect 16764 13889 16773 13923
rect 16773 13889 16807 13923
rect 16807 13889 16816 13923
rect 16764 13880 16816 13889
rect 18604 13880 18656 13932
rect 21824 13923 21876 13932
rect 21824 13889 21833 13923
rect 21833 13889 21867 13923
rect 21867 13889 21876 13923
rect 21824 13880 21876 13889
rect 44548 13880 44600 13932
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 22836 13855 22888 13864
rect 22836 13821 22845 13855
rect 22845 13821 22879 13855
rect 22879 13821 22888 13855
rect 22836 13812 22888 13821
rect 3424 13744 3476 13796
rect 14556 13744 14608 13796
rect 16764 13676 16816 13728
rect 16948 13676 17000 13728
rect 46480 13676 46532 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 22192 13472 22244 13524
rect 14832 13404 14884 13456
rect 16764 13379 16816 13388
rect 16764 13345 16773 13379
rect 16773 13345 16807 13379
rect 16807 13345 16816 13379
rect 16764 13336 16816 13345
rect 46480 13379 46532 13388
rect 46480 13345 46489 13379
rect 46489 13345 46523 13379
rect 46523 13345 46532 13379
rect 46480 13336 46532 13345
rect 22468 13268 22520 13320
rect 46296 13311 46348 13320
rect 46296 13277 46305 13311
rect 46305 13277 46339 13311
rect 46339 13277 46348 13311
rect 46296 13268 46348 13277
rect 17960 13200 18012 13252
rect 48136 13243 48188 13252
rect 48136 13209 48145 13243
rect 48145 13209 48179 13243
rect 48179 13209 48188 13243
rect 48136 13200 48188 13209
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 16948 12903 17000 12912
rect 16948 12869 16957 12903
rect 16957 12869 16991 12903
rect 16991 12869 17000 12903
rect 16948 12860 17000 12869
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 16580 12792 16632 12844
rect 46296 12792 46348 12844
rect 18604 12767 18656 12776
rect 18604 12733 18613 12767
rect 18613 12733 18647 12767
rect 18647 12733 18656 12767
rect 18604 12724 18656 12733
rect 26424 12588 26476 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 46296 11500 46348 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 46296 11203 46348 11212
rect 46296 11169 46305 11203
rect 46305 11169 46339 11203
rect 46339 11169 46348 11203
rect 46296 11160 46348 11169
rect 46480 11067 46532 11076
rect 46480 11033 46489 11067
rect 46489 11033 46523 11067
rect 46523 11033 46532 11067
rect 46480 11024 46532 11033
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 3148 10956 3200 11008
rect 10784 10956 10836 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 46480 10752 46532 10804
rect 29552 10616 29604 10668
rect 36636 10616 36688 10668
rect 47400 10616 47452 10668
rect 46296 10455 46348 10464
rect 46296 10421 46305 10455
rect 46305 10421 46339 10455
rect 46339 10421 46348 10455
rect 46296 10412 46348 10421
rect 46480 10412 46532 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 46480 10115 46532 10124
rect 46480 10081 46489 10115
rect 46489 10081 46523 10115
rect 46523 10081 46532 10115
rect 46480 10072 46532 10081
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 47860 9571 47912 9580
rect 47860 9537 47869 9571
rect 47869 9537 47903 9571
rect 47903 9537 47912 9571
rect 47860 9528 47912 9537
rect 46112 9392 46164 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 47768 8891 47820 8900
rect 47768 8857 47777 8891
rect 47777 8857 47811 8891
rect 47811 8857 47820 8891
rect 47768 8848 47820 8857
rect 29828 8780 29880 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 45284 8440 45336 8492
rect 1860 8372 1912 8424
rect 18604 8236 18656 8288
rect 36176 8236 36228 8288
rect 45744 8236 45796 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 36176 8032 36228 8084
rect 46848 8032 46900 8084
rect 45100 7964 45152 8016
rect 47492 7896 47544 7948
rect 47308 7871 47360 7880
rect 47308 7837 47317 7871
rect 47317 7837 47351 7871
rect 47351 7837 47360 7871
rect 47308 7828 47360 7837
rect 45284 7803 45336 7812
rect 45284 7769 45293 7803
rect 45293 7769 45327 7803
rect 45327 7769 45336 7803
rect 45284 7760 45336 7769
rect 45376 7803 45428 7812
rect 45376 7769 45385 7803
rect 45385 7769 45419 7803
rect 45419 7769 45428 7803
rect 45376 7760 45428 7769
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 45100 7488 45152 7540
rect 45744 7463 45796 7472
rect 45744 7429 45753 7463
rect 45753 7429 45787 7463
rect 45787 7429 45796 7463
rect 45744 7420 45796 7429
rect 48228 7352 48280 7404
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3424 6808 3476 6860
rect 23940 6808 23992 6860
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 42340 6400 42392 6452
rect 47952 6307 48004 6316
rect 47952 6273 47961 6307
rect 47961 6273 47995 6307
rect 47995 6273 48004 6307
rect 47952 6264 48004 6273
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 40132 5695 40184 5704
rect 40132 5661 40141 5695
rect 40141 5661 40175 5695
rect 40175 5661 40184 5695
rect 40132 5652 40184 5661
rect 40224 5559 40276 5568
rect 40224 5525 40233 5559
rect 40233 5525 40267 5559
rect 40267 5525 40276 5559
rect 40224 5516 40276 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3976 5244 4028 5296
rect 37464 5287 37516 5296
rect 37464 5253 37473 5287
rect 37473 5253 37507 5287
rect 37507 5253 37516 5287
rect 37464 5244 37516 5253
rect 40132 5312 40184 5364
rect 40316 5312 40368 5364
rect 40592 5312 40644 5364
rect 18328 5219 18380 5228
rect 18328 5185 18337 5219
rect 18337 5185 18371 5219
rect 18371 5185 18380 5219
rect 18328 5176 18380 5185
rect 23848 5176 23900 5228
rect 23204 5108 23256 5160
rect 37372 5151 37424 5160
rect 37372 5117 37381 5151
rect 37381 5117 37415 5151
rect 37415 5117 37424 5151
rect 39212 5176 39264 5228
rect 40592 5176 40644 5228
rect 40868 5219 40920 5228
rect 40868 5185 40877 5219
rect 40877 5185 40911 5219
rect 40911 5185 40920 5219
rect 40868 5176 40920 5185
rect 37372 5108 37424 5117
rect 38476 5108 38528 5160
rect 40316 5108 40368 5160
rect 42524 5244 42576 5296
rect 47952 5176 48004 5228
rect 43628 5108 43680 5160
rect 43812 5108 43864 5160
rect 24952 5040 25004 5092
rect 18052 4972 18104 5024
rect 22468 4972 22520 5024
rect 22928 4972 22980 5024
rect 40408 4972 40460 5024
rect 40868 5015 40920 5024
rect 40868 4981 40877 5015
rect 40877 4981 40911 5015
rect 40911 4981 40920 5015
rect 40868 4972 40920 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 39212 4811 39264 4820
rect 39212 4777 39221 4811
rect 39221 4777 39255 4811
rect 39255 4777 39264 4811
rect 39212 4768 39264 4777
rect 39304 4768 39356 4820
rect 40868 4768 40920 4820
rect 42524 4811 42576 4820
rect 42524 4777 42533 4811
rect 42533 4777 42567 4811
rect 42567 4777 42576 4811
rect 42524 4768 42576 4777
rect 23664 4700 23716 4752
rect 24400 4632 24452 4684
rect 38476 4675 38528 4684
rect 38476 4641 38485 4675
rect 38485 4641 38519 4675
rect 38519 4641 38528 4675
rect 38476 4632 38528 4641
rect 40224 4675 40276 4684
rect 40224 4641 40233 4675
rect 40233 4641 40267 4675
rect 40267 4641 40276 4675
rect 40224 4632 40276 4641
rect 40408 4675 40460 4684
rect 40408 4641 40417 4675
rect 40417 4641 40451 4675
rect 40451 4641 40460 4675
rect 40408 4632 40460 4641
rect 45376 4632 45428 4684
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 18236 4564 18288 4616
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 21916 4564 21968 4616
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22100 4564 22152 4573
rect 22468 4564 22520 4616
rect 23480 4564 23532 4616
rect 25504 4564 25556 4616
rect 40132 4564 40184 4616
rect 42892 4564 42944 4616
rect 45008 4564 45060 4616
rect 46848 4564 46900 4616
rect 20996 4496 21048 4548
rect 23020 4496 23072 4548
rect 37280 4496 37332 4548
rect 37556 4539 37608 4548
rect 37556 4505 37565 4539
rect 37565 4505 37599 4539
rect 37599 4505 37608 4539
rect 37556 4496 37608 4505
rect 42156 4496 42208 4548
rect 42616 4496 42668 4548
rect 18144 4471 18196 4480
rect 18144 4437 18153 4471
rect 18153 4437 18187 4471
rect 18187 4437 18196 4471
rect 18144 4428 18196 4437
rect 19340 4471 19392 4480
rect 19340 4437 19349 4471
rect 19349 4437 19383 4471
rect 19383 4437 19392 4471
rect 19340 4428 19392 4437
rect 21456 4428 21508 4480
rect 24308 4428 24360 4480
rect 46480 4428 46532 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 17224 4224 17276 4276
rect 20996 4267 21048 4276
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 5264 4088 5316 4140
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 13728 4131 13780 4140
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 18144 4156 18196 4208
rect 17960 4131 18012 4140
rect 17960 4097 17969 4131
rect 17969 4097 18003 4131
rect 18003 4097 18012 4131
rect 17960 4088 18012 4097
rect 3424 3952 3476 4004
rect 17224 3952 17276 4004
rect 18328 4020 18380 4072
rect 20996 4233 21005 4267
rect 21005 4233 21039 4267
rect 21039 4233 21048 4267
rect 20996 4224 21048 4233
rect 21916 4267 21968 4276
rect 21916 4233 21925 4267
rect 21925 4233 21959 4267
rect 21959 4233 21968 4267
rect 21916 4224 21968 4233
rect 37464 4224 37516 4276
rect 40592 4224 40644 4276
rect 18972 4131 19024 4140
rect 18972 4097 18981 4131
rect 18981 4097 19015 4131
rect 19015 4097 19024 4131
rect 18972 4088 19024 4097
rect 19064 4088 19116 4140
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 21364 4088 21416 4140
rect 21456 4088 21508 4140
rect 23112 4131 23164 4140
rect 18512 3952 18564 4004
rect 18604 3952 18656 4004
rect 1400 3884 1452 3936
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 2964 3927 3016 3936
rect 2964 3893 2973 3927
rect 2973 3893 3007 3927
rect 3007 3893 3016 3927
rect 2964 3884 3016 3893
rect 5908 3884 5960 3936
rect 6920 3884 6972 3936
rect 8116 3884 8168 3936
rect 9404 3884 9456 3936
rect 11520 3884 11572 3936
rect 14004 3884 14056 3936
rect 17500 3884 17552 3936
rect 18788 3884 18840 3936
rect 20812 3952 20864 4004
rect 23112 4097 23121 4131
rect 23121 4097 23155 4131
rect 23155 4097 23164 4131
rect 23112 4088 23164 4097
rect 23204 4131 23256 4140
rect 23204 4097 23213 4131
rect 23213 4097 23247 4131
rect 23247 4097 23256 4131
rect 23204 4088 23256 4097
rect 24492 4088 24544 4140
rect 24860 4088 24912 4140
rect 40040 4199 40092 4208
rect 40040 4165 40049 4199
rect 40049 4165 40083 4199
rect 40083 4165 40092 4199
rect 40040 4156 40092 4165
rect 40500 4199 40552 4208
rect 40500 4165 40509 4199
rect 40509 4165 40543 4199
rect 40543 4165 40552 4199
rect 40500 4156 40552 4165
rect 42800 4156 42852 4208
rect 43812 4199 43864 4208
rect 43812 4165 43821 4199
rect 43821 4165 43855 4199
rect 43855 4165 43864 4199
rect 43812 4156 43864 4165
rect 47768 4199 47820 4208
rect 47768 4165 47777 4199
rect 47777 4165 47811 4199
rect 47811 4165 47820 4199
rect 47768 4156 47820 4165
rect 23848 4063 23900 4072
rect 23848 4029 23857 4063
rect 23857 4029 23891 4063
rect 23891 4029 23900 4063
rect 23848 4020 23900 4029
rect 24952 4020 25004 4072
rect 37740 4088 37792 4140
rect 40224 4088 40276 4140
rect 46756 4131 46808 4140
rect 46756 4097 46765 4131
rect 46765 4097 46799 4131
rect 46799 4097 46808 4131
rect 46756 4088 46808 4097
rect 26240 4020 26292 4072
rect 26884 4020 26936 4072
rect 30012 4020 30064 4072
rect 37280 4020 37332 4072
rect 39948 4020 40000 4072
rect 45284 4020 45336 4072
rect 20076 3884 20128 3936
rect 20904 3884 20956 3936
rect 22468 3884 22520 3936
rect 29552 3952 29604 4004
rect 23572 3884 23624 3936
rect 30932 3884 30984 3936
rect 32680 3884 32732 3936
rect 46296 3927 46348 3936
rect 46296 3893 46305 3927
rect 46305 3893 46339 3927
rect 46339 3893 46348 3927
rect 46296 3884 46348 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 18236 3680 18288 3732
rect 18696 3680 18748 3732
rect 20168 3680 20220 3732
rect 20260 3680 20312 3732
rect 21364 3680 21416 3732
rect 23112 3680 23164 3732
rect 24492 3723 24544 3732
rect 24492 3689 24501 3723
rect 24501 3689 24535 3723
rect 24535 3689 24544 3723
rect 24492 3680 24544 3689
rect 24584 3680 24636 3732
rect 30932 3680 30984 3732
rect 31116 3680 31168 3732
rect 664 3612 716 3664
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 2228 3544 2280 3596
rect 5264 3612 5316 3664
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 9496 3544 9548 3596
rect 9588 3544 9640 3596
rect 2044 3408 2096 3460
rect 5264 3519 5316 3528
rect 5264 3485 5273 3519
rect 5273 3485 5307 3519
rect 5307 3485 5316 3519
rect 5264 3476 5316 3485
rect 7932 3476 7984 3528
rect 9404 3451 9456 3460
rect 9404 3417 9413 3451
rect 9413 3417 9447 3451
rect 9447 3417 9456 3451
rect 9404 3408 9456 3417
rect 18144 3612 18196 3664
rect 18328 3612 18380 3664
rect 26700 3612 26752 3664
rect 32864 3680 32916 3732
rect 39304 3680 39356 3732
rect 40132 3723 40184 3732
rect 40132 3689 40141 3723
rect 40141 3689 40175 3723
rect 40175 3689 40184 3723
rect 40132 3680 40184 3689
rect 13820 3476 13872 3528
rect 33784 3612 33836 3664
rect 34060 3612 34112 3664
rect 42524 3612 42576 3664
rect 46572 3612 46624 3664
rect 46296 3587 46348 3596
rect 17500 3476 17552 3528
rect 17776 3476 17828 3528
rect 19340 3476 19392 3528
rect 16120 3408 16172 3460
rect 18236 3408 18288 3460
rect 18972 3408 19024 3460
rect 11704 3340 11756 3392
rect 17408 3340 17460 3392
rect 18144 3340 18196 3392
rect 20352 3519 20404 3528
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 20352 3476 20404 3485
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 20904 3476 20956 3528
rect 22284 3476 22336 3528
rect 23020 3519 23072 3528
rect 23020 3485 23029 3519
rect 23029 3485 23063 3519
rect 23063 3485 23072 3519
rect 23020 3476 23072 3485
rect 23664 3519 23716 3528
rect 23664 3485 23673 3519
rect 23673 3485 23707 3519
rect 23707 3485 23716 3519
rect 23664 3476 23716 3485
rect 24400 3519 24452 3528
rect 24400 3485 24409 3519
rect 24409 3485 24443 3519
rect 24443 3485 24452 3519
rect 24400 3476 24452 3485
rect 25504 3519 25556 3528
rect 25504 3485 25513 3519
rect 25513 3485 25547 3519
rect 25547 3485 25556 3519
rect 25504 3476 25556 3485
rect 20720 3408 20772 3460
rect 22100 3408 22152 3460
rect 19984 3340 20036 3392
rect 20628 3340 20680 3392
rect 24584 3340 24636 3392
rect 25780 3408 25832 3460
rect 33876 3519 33928 3528
rect 32864 3340 32916 3392
rect 33140 3383 33192 3392
rect 33140 3349 33149 3383
rect 33149 3349 33183 3383
rect 33183 3349 33192 3383
rect 33140 3340 33192 3349
rect 33876 3485 33885 3519
rect 33885 3485 33919 3519
rect 33919 3485 33928 3519
rect 33876 3476 33928 3485
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 40040 3519 40092 3528
rect 40040 3485 40049 3519
rect 40049 3485 40083 3519
rect 40083 3485 40092 3519
rect 40040 3476 40092 3485
rect 40776 3519 40828 3528
rect 40776 3485 40785 3519
rect 40785 3485 40819 3519
rect 40819 3485 40828 3519
rect 40776 3476 40828 3485
rect 39672 3408 39724 3460
rect 41144 3340 41196 3392
rect 43904 3519 43956 3528
rect 43904 3485 43913 3519
rect 43913 3485 43947 3519
rect 43947 3485 43956 3519
rect 43904 3476 43956 3485
rect 45192 3519 45244 3528
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 42616 3451 42668 3460
rect 42616 3417 42625 3451
rect 42625 3417 42659 3451
rect 42659 3417 42668 3451
rect 42616 3408 42668 3417
rect 47492 3408 47544 3460
rect 48964 3408 49016 3460
rect 43076 3340 43128 3392
rect 45376 3340 45428 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 8852 3136 8904 3188
rect 37464 3136 37516 3188
rect 37740 3179 37792 3188
rect 37740 3145 37749 3179
rect 37749 3145 37783 3179
rect 37783 3145 37792 3179
rect 37740 3136 37792 3145
rect 39672 3179 39724 3188
rect 39672 3145 39681 3179
rect 39681 3145 39715 3179
rect 39715 3145 39724 3179
rect 39672 3136 39724 3145
rect 40776 3136 40828 3188
rect 47676 3136 47728 3188
rect 2964 3068 3016 3120
rect 8116 3111 8168 3120
rect 8116 3077 8125 3111
rect 8125 3077 8159 3111
rect 8159 3077 8168 3111
rect 8116 3068 8168 3077
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 14004 3111 14056 3120
rect 14004 3077 14013 3111
rect 14013 3077 14047 3111
rect 14047 3077 14056 3111
rect 14004 3068 14056 3077
rect 17776 3111 17828 3120
rect 17776 3077 17785 3111
rect 17785 3077 17819 3111
rect 17819 3077 17828 3111
rect 17776 3068 17828 3077
rect 19064 3068 19116 3120
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 7932 3043 7984 3052
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 2964 2975 3016 2984
rect 2964 2941 2973 2975
rect 2973 2941 3007 2975
rect 3007 2941 3016 2975
rect 2964 2932 3016 2941
rect 7748 2932 7800 2984
rect 10968 2932 11020 2984
rect 14188 2932 14240 2984
rect 15200 2932 15252 2984
rect 6736 2839 6788 2848
rect 6736 2805 6745 2839
rect 6745 2805 6779 2839
rect 6779 2805 6788 2839
rect 6736 2796 6788 2805
rect 9036 2796 9088 2848
rect 9588 2796 9640 2848
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 19708 3068 19760 3120
rect 21088 3068 21140 3120
rect 22468 3111 22520 3120
rect 22468 3077 22477 3111
rect 22477 3077 22511 3111
rect 22511 3077 22520 3111
rect 22468 3068 22520 3077
rect 24308 3068 24360 3120
rect 26056 3068 26108 3120
rect 26240 3068 26292 3120
rect 26700 3068 26752 3120
rect 32220 3068 32272 3120
rect 33140 3111 33192 3120
rect 33140 3077 33149 3111
rect 33149 3077 33183 3111
rect 33183 3077 33192 3111
rect 33140 3068 33192 3077
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 27160 3043 27212 3052
rect 20352 2932 20404 2984
rect 19892 2864 19944 2916
rect 19984 2864 20036 2916
rect 22560 2932 22612 2984
rect 20536 2864 20588 2916
rect 24860 2864 24912 2916
rect 25136 2864 25188 2916
rect 25780 2864 25832 2916
rect 27160 3009 27169 3043
rect 27169 3009 27203 3043
rect 27203 3009 27212 3043
rect 27160 3000 27212 3009
rect 37556 3000 37608 3052
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 42616 3068 42668 3120
rect 43076 3111 43128 3120
rect 43076 3077 43085 3111
rect 43085 3077 43119 3111
rect 43119 3077 43128 3111
rect 43076 3068 43128 3077
rect 45376 3111 45428 3120
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 40592 3000 40644 3052
rect 41236 3000 41288 3052
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 48320 3000 48372 3052
rect 26056 2796 26108 2848
rect 33876 2864 33928 2916
rect 39948 2932 40000 2984
rect 40040 2932 40092 2984
rect 40408 2932 40460 2984
rect 40224 2864 40276 2916
rect 43904 2932 43956 2984
rect 43168 2864 43220 2916
rect 47676 2932 47728 2984
rect 37372 2839 37424 2848
rect 37372 2805 37381 2839
rect 37381 2805 37415 2839
rect 37415 2805 37424 2839
rect 37372 2796 37424 2805
rect 37464 2796 37516 2848
rect 45652 2796 45704 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 6920 2524 6972 2576
rect 9312 2592 9364 2644
rect 15200 2592 15252 2644
rect 6736 2499 6788 2508
rect 6736 2465 6745 2499
rect 6745 2465 6779 2499
rect 6779 2465 6788 2499
rect 6736 2456 6788 2465
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 7196 2456 7248 2508
rect 17316 2592 17368 2644
rect 17960 2592 18012 2644
rect 19248 2592 19300 2644
rect 21272 2524 21324 2576
rect 24216 2592 24268 2644
rect 26240 2592 26292 2644
rect 27160 2524 27212 2576
rect 5172 2388 5224 2440
rect 8484 2388 8536 2440
rect 1308 2320 1360 2372
rect 2596 2320 2648 2372
rect 15476 2320 15528 2372
rect 16120 2388 16172 2440
rect 17408 2431 17460 2440
rect 17408 2397 17417 2431
rect 17417 2397 17451 2431
rect 17451 2397 17460 2431
rect 17408 2388 17460 2397
rect 18052 2431 18104 2440
rect 18052 2397 18061 2431
rect 18061 2397 18095 2431
rect 18095 2397 18104 2431
rect 18052 2388 18104 2397
rect 22928 2431 22980 2440
rect 22928 2397 22937 2431
rect 22937 2397 22971 2431
rect 22971 2397 22980 2431
rect 22928 2388 22980 2397
rect 20628 2320 20680 2372
rect 21916 2320 21968 2372
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 2136 2252 2188 2261
rect 4068 2252 4120 2304
rect 7196 2252 7248 2304
rect 15752 2295 15804 2304
rect 15752 2261 15761 2295
rect 15761 2261 15795 2295
rect 15795 2261 15804 2295
rect 15752 2252 15804 2261
rect 17316 2252 17368 2304
rect 22836 2252 22888 2304
rect 24492 2320 24544 2372
rect 27436 2456 27488 2508
rect 28356 2592 28408 2644
rect 29736 2635 29788 2644
rect 29736 2601 29745 2635
rect 29745 2601 29779 2635
rect 29779 2601 29788 2635
rect 29736 2592 29788 2601
rect 32312 2592 32364 2644
rect 35624 2592 35676 2644
rect 36360 2635 36412 2644
rect 36360 2601 36369 2635
rect 36369 2601 36403 2635
rect 36403 2601 36412 2635
rect 36360 2592 36412 2601
rect 40592 2635 40644 2644
rect 30104 2524 30156 2576
rect 24860 2388 24912 2440
rect 26424 2388 26476 2440
rect 27712 2388 27764 2440
rect 29644 2388 29696 2440
rect 35900 2524 35952 2576
rect 35992 2524 36044 2576
rect 40592 2601 40601 2635
rect 40601 2601 40635 2635
rect 40635 2601 40644 2635
rect 40592 2592 40644 2601
rect 42892 2635 42944 2644
rect 33692 2456 33744 2508
rect 40500 2524 40552 2576
rect 42432 2524 42484 2576
rect 42892 2601 42901 2635
rect 42901 2601 42935 2635
rect 42935 2601 42944 2635
rect 42892 2592 42944 2601
rect 35440 2388 35492 2440
rect 27068 2320 27120 2372
rect 28356 2320 28408 2372
rect 29736 2320 29788 2372
rect 35992 2320 36044 2372
rect 36084 2320 36136 2372
rect 24952 2252 25004 2304
rect 26240 2252 26292 2304
rect 35624 2252 35676 2304
rect 40224 2388 40276 2440
rect 40408 2431 40460 2440
rect 40408 2397 40417 2431
rect 40417 2397 40451 2431
rect 40451 2397 40460 2431
rect 40408 2388 40460 2397
rect 40592 2388 40644 2440
rect 42800 2388 42852 2440
rect 47860 2499 47912 2508
rect 47860 2465 47869 2499
rect 47869 2465 47903 2499
rect 47903 2465 47912 2499
rect 47860 2456 47912 2465
rect 43812 2388 43864 2440
rect 38016 2320 38068 2372
rect 39304 2320 39356 2372
rect 47032 2388 47084 2440
rect 48044 2388 48096 2440
rect 37648 2252 37700 2304
rect 46388 2320 46440 2372
rect 41328 2252 41380 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 27436 2048 27488 2100
rect 32036 2048 32088 2100
rect 35900 2048 35952 2100
rect 40684 2048 40736 2100
rect 22376 1980 22428 2032
rect 41328 1980 41380 2032
rect 2136 1912 2188 1964
rect 26976 1912 27028 1964
rect 15752 1844 15804 1896
rect 37372 1844 37424 1896
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4752 49314
rect 4498 49200 4610 49286
rect 32 21962 60 49200
rect 1858 47696 1914 47705
rect 1858 47631 1914 47640
rect 1872 46646 1900 47631
rect 1964 47054 1992 49200
rect 2044 47456 2096 47462
rect 2044 47398 2096 47404
rect 2056 47122 2084 47398
rect 2044 47116 2096 47122
rect 2044 47058 2096 47064
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2608 46918 2636 49200
rect 3252 47054 3280 49200
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3422 47016 3478 47025
rect 3056 46980 3108 46986
rect 3422 46951 3478 46960
rect 3056 46922 3108 46928
rect 2596 46912 2648 46918
rect 2596 46854 2648 46860
rect 1860 46640 1912 46646
rect 1860 46582 1912 46588
rect 2320 46368 2372 46374
rect 2872 46368 2924 46374
rect 2320 46310 2372 46316
rect 2778 46336 2834 46345
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1492 43240 1544 43246
rect 1492 43182 1544 43188
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1400 40520 1452 40526
rect 1400 40462 1452 40468
rect 1412 40225 1440 40462
rect 1398 40216 1454 40225
rect 1398 40151 1454 40160
rect 1400 35488 1452 35494
rect 1400 35430 1452 35436
rect 1412 33522 1440 35430
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1398 33416 1454 33425
rect 1398 33351 1454 33360
rect 1412 32978 1440 33351
rect 1400 32972 1452 32978
rect 1400 32914 1452 32920
rect 1504 26234 1532 43182
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1584 41540 1636 41546
rect 1858 41511 1914 41520
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 2136 41132 2188 41138
rect 2136 41074 2188 41080
rect 1676 40384 1728 40390
rect 1676 40326 1728 40332
rect 1688 35894 1716 40326
rect 1952 37256 2004 37262
rect 1952 37198 2004 37204
rect 1964 36786 1992 37198
rect 1952 36780 2004 36786
rect 1952 36722 2004 36728
rect 1688 35866 1808 35894
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1596 35465 1624 35634
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1676 33108 1728 33114
rect 1676 33050 1728 33056
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 1596 31822 1624 32671
rect 1688 32026 1716 33050
rect 1676 32020 1728 32026
rect 1676 31962 1728 31968
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1780 28218 1808 35866
rect 2044 32224 2096 32230
rect 2044 32166 2096 32172
rect 2056 31346 2084 32166
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 1768 28212 1820 28218
rect 1768 28154 1820 28160
rect 1504 26206 1716 26234
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1412 23225 1440 23666
rect 1582 23624 1638 23633
rect 1582 23559 1584 23568
rect 1636 23559 1638 23568
rect 1584 23530 1636 23536
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 20 21956 72 21962
rect 20 21898 72 21904
rect 1688 19514 1716 26206
rect 1860 25288 1912 25294
rect 1858 25256 1860 25265
rect 1912 25256 1914 25265
rect 1858 25191 1914 25200
rect 1860 25152 1912 25158
rect 1860 25094 1912 25100
rect 1676 19508 1728 19514
rect 1676 19450 1728 19456
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17785 1440 18226
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1780 17202 1808 17614
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1872 8430 1900 25094
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 2056 18970 2084 19246
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2148 17678 2176 41074
rect 2332 25362 2360 46310
rect 2872 46310 2924 46316
rect 2778 46271 2834 46280
rect 2792 45354 2820 46271
rect 2884 45422 2912 46310
rect 2964 45824 3016 45830
rect 2964 45766 3016 45772
rect 2976 45558 3004 45766
rect 2964 45552 3016 45558
rect 2964 45494 3016 45500
rect 2872 45416 2924 45422
rect 2872 45358 2924 45364
rect 2780 45348 2832 45354
rect 2780 45290 2832 45296
rect 2962 36816 3018 36825
rect 2962 36751 3018 36760
rect 2976 36718 3004 36751
rect 2872 36712 2924 36718
rect 2872 36654 2924 36660
rect 2964 36712 3016 36718
rect 2964 36654 3016 36660
rect 2884 36378 2912 36654
rect 2872 36372 2924 36378
rect 2872 36314 2924 36320
rect 2780 32904 2832 32910
rect 2780 32846 2832 32852
rect 2792 32502 2820 32846
rect 2780 32496 2832 32502
rect 2780 32438 2832 32444
rect 2596 32360 2648 32366
rect 2596 32302 2648 32308
rect 2320 25356 2372 25362
rect 2320 25298 2372 25304
rect 2608 21078 2636 32302
rect 2778 32056 2834 32065
rect 2778 31991 2834 32000
rect 2792 31278 2820 31991
rect 2964 31680 3016 31686
rect 2964 31622 3016 31628
rect 2976 31414 3004 31622
rect 2964 31408 3016 31414
rect 2964 31350 3016 31356
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 3068 21690 3096 46922
rect 3148 45960 3200 45966
rect 3148 45902 3200 45908
rect 3160 32570 3188 45902
rect 3330 44976 3386 44985
rect 3330 44911 3386 44920
rect 3344 38894 3372 44911
rect 3332 38888 3384 38894
rect 3332 38830 3384 38836
rect 3148 32564 3200 32570
rect 3148 32506 3200 32512
rect 3160 31822 3188 32506
rect 3148 31816 3200 31822
rect 3148 31758 3200 31764
rect 3056 21684 3108 21690
rect 3056 21626 3108 21632
rect 3436 21146 3464 46951
rect 3896 46594 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4724 47054 4752 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49314 7186 50000
rect 7074 49286 7328 49314
rect 7074 49200 7186 49286
rect 5828 47054 5856 49200
rect 6644 47524 6696 47530
rect 6644 47466 6696 47472
rect 6656 47122 6684 47466
rect 6644 47116 6696 47122
rect 6644 47058 6696 47064
rect 7300 47054 7328 49286
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49200 13626 50000
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49314 16202 50000
rect 16090 49286 16528 49314
rect 16090 49200 16202 49286
rect 4712 47048 4764 47054
rect 4712 46990 4764 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7288 47048 7340 47054
rect 7288 46990 7340 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 3896 46566 4016 46594
rect 3988 46510 4016 46566
rect 3884 46504 3936 46510
rect 3884 46446 3936 46452
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 3896 46170 3924 46446
rect 3884 46164 3936 46170
rect 3884 46106 3936 46112
rect 3606 43616 3662 43625
rect 3606 43551 3662 43560
rect 3514 39536 3570 39545
rect 3514 39471 3570 39480
rect 3528 39030 3556 39471
rect 3516 39024 3568 39030
rect 3516 38966 3568 38972
rect 3516 38888 3568 38894
rect 3516 38830 3568 38836
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 2596 21072 2648 21078
rect 2596 21014 2648 21020
rect 3056 20596 3108 20602
rect 3056 20538 3108 20544
rect 3068 19825 3096 20538
rect 3528 20058 3556 38830
rect 3620 24614 3648 43551
rect 3700 33448 3752 33454
rect 3700 33390 3752 33396
rect 3712 33114 3740 33390
rect 3700 33108 3752 33114
rect 3700 33050 3752 33056
rect 3882 31376 3938 31385
rect 3882 31311 3938 31320
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3896 23322 3924 31311
rect 3974 28656 4030 28665
rect 3974 28591 4030 28600
rect 3988 27674 4016 28591
rect 3976 27668 4028 27674
rect 3976 27610 4028 27616
rect 3884 23316 3936 23322
rect 3884 23258 3936 23264
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3054 19816 3110 19825
rect 3054 19751 3110 19760
rect 3056 19440 3108 19446
rect 3056 19382 3108 19388
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2792 19145 2820 19246
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 3068 18970 3096 19382
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2976 18426 3004 18702
rect 3330 18456 3386 18465
rect 2964 18420 3016 18426
rect 3330 18391 3386 18400
rect 2964 18362 3016 18368
rect 3344 18154 3372 18391
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17270 1992 17478
rect 2148 17338 2176 17614
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 1952 17264 2004 17270
rect 1952 17206 2004 17212
rect 2780 17128 2832 17134
rect 3528 17105 3556 17546
rect 2780 17070 2832 17076
rect 3514 17096 3570 17105
rect 2792 16425 2820 17070
rect 3514 17031 3570 17040
rect 2778 16416 2834 16425
rect 2778 16351 2834 16360
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 2148 4146 2176 14350
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10305 3188 10950
rect 3146 10296 3202 10305
rect 3146 10231 3202 10240
rect 3344 7585 3372 14214
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3436 13705 3464 13738
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 3330 7576 3386 7585
rect 3330 7511 3386 7520
rect 4080 6914 4108 46922
rect 7472 46912 7524 46918
rect 7472 46854 7524 46860
rect 4620 46436 4672 46442
rect 4620 46378 4672 46384
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4632 46170 4660 46378
rect 4620 46164 4672 46170
rect 4620 46106 4672 46112
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 6644 36168 6696 36174
rect 6644 36110 6696 36116
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4620 33448 4672 33454
rect 4620 33390 4672 33396
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4632 32366 4660 33390
rect 4620 32360 4672 32366
rect 4620 32302 4672 32308
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4632 18358 4660 32302
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3422 6896 3478 6905
rect 3422 6831 3424 6840
rect 3476 6831 3478 6840
rect 3988 6886 4108 6914
rect 3424 6802 3476 6808
rect 3988 5302 4016 6886
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 3424 4004 3476 4010
rect 3424 3946 3476 3952
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 664 3664 716 3670
rect 664 3606 716 3612
rect 676 800 704 3606
rect 1412 3602 1440 3878
rect 2240 3602 2268 3878
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2044 3460 2096 3466
rect 2044 3402 2096 3408
rect 2056 3058 2084 3402
rect 2976 3126 3004 3878
rect 3436 3505 3464 3946
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 5276 3670 5304 4082
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5264 3664 5316 3670
rect 3882 3632 3938 3641
rect 5264 3606 5316 3612
rect 3882 3567 3938 3576
rect 3422 3496 3478 3505
rect 3422 3431 3478 3440
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 1320 800 1348 2314
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2148 1970 2176 2246
rect 2136 1964 2188 1970
rect 2136 1906 2188 1912
rect 2608 800 2636 2314
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 2976 785 3004 2926
rect 3896 800 3924 3567
rect 5276 3534 5304 3606
rect 5920 3602 5948 3878
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4080 1465 4108 2246
rect 4066 1456 4122 1465
rect 4066 1391 4122 1400
rect 5184 800 5212 2382
rect 6472 800 6500 3538
rect 6656 3058 6684 36110
rect 7484 27062 7512 46854
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 10508 46368 10560 46374
rect 10508 46310 10560 46316
rect 10520 46034 10548 46310
rect 10980 46034 11008 49200
rect 11624 47054 11652 49200
rect 12268 47054 12296 49200
rect 12912 47054 12940 49200
rect 13360 47592 13412 47598
rect 13360 47534 13412 47540
rect 13372 47258 13400 47534
rect 13360 47252 13412 47258
rect 13360 47194 13412 47200
rect 11612 47048 11664 47054
rect 11612 46990 11664 46996
rect 12256 47048 12308 47054
rect 12256 46990 12308 46996
rect 12900 47048 12952 47054
rect 12900 46990 12952 46996
rect 11704 46980 11756 46986
rect 11704 46922 11756 46928
rect 12440 46980 12492 46986
rect 12440 46922 12492 46928
rect 10508 46028 10560 46034
rect 10508 45970 10560 45976
rect 10968 46028 11020 46034
rect 10968 45970 11020 45976
rect 10692 45892 10744 45898
rect 10692 45834 10744 45840
rect 10600 45824 10652 45830
rect 10600 45766 10652 45772
rect 8312 45526 8432 45554
rect 7564 39024 7616 39030
rect 7564 38966 7616 38972
rect 7576 27946 7604 38966
rect 8312 32502 8340 45526
rect 10612 45490 10640 45766
rect 10704 45626 10732 45834
rect 10692 45620 10744 45626
rect 10692 45562 10744 45568
rect 10600 45484 10652 45490
rect 10600 45426 10652 45432
rect 9588 32904 9640 32910
rect 9588 32846 9640 32852
rect 8300 32496 8352 32502
rect 8300 32438 8352 32444
rect 9600 31822 9628 32846
rect 9772 32360 9824 32366
rect 9772 32302 9824 32308
rect 10784 32360 10836 32366
rect 10784 32302 10836 32308
rect 9784 32026 9812 32302
rect 10796 32026 10824 32302
rect 9772 32020 9824 32026
rect 9772 31962 9824 31968
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 11716 31958 11744 46922
rect 12452 37262 12480 46922
rect 13556 46918 13584 49200
rect 14200 47954 14228 49200
rect 14200 47926 14320 47954
rect 13544 46912 13596 46918
rect 13544 46854 13596 46860
rect 14292 46510 14320 47926
rect 14740 46980 14792 46986
rect 14740 46922 14792 46928
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 14200 46170 14228 46446
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 12440 37256 12492 37262
rect 12440 37198 12492 37204
rect 13360 33448 13412 33454
rect 13360 33390 13412 33396
rect 14188 33448 14240 33454
rect 14188 33390 14240 33396
rect 13268 32972 13320 32978
rect 13268 32914 13320 32920
rect 12532 32496 12584 32502
rect 12532 32438 12584 32444
rect 11796 32360 11848 32366
rect 11796 32302 11848 32308
rect 11808 32026 11836 32302
rect 12544 32026 12572 32438
rect 13280 32366 13308 32914
rect 13268 32360 13320 32366
rect 13268 32302 13320 32308
rect 12992 32224 13044 32230
rect 12992 32166 13044 32172
rect 11796 32020 11848 32026
rect 11796 31962 11848 31968
rect 12532 32020 12584 32026
rect 12532 31962 12584 31968
rect 11704 31952 11756 31958
rect 11704 31894 11756 31900
rect 9588 31816 9640 31822
rect 9588 31758 9640 31764
rect 10692 31816 10744 31822
rect 10692 31758 10744 31764
rect 12440 31816 12492 31822
rect 12440 31758 12492 31764
rect 9312 29844 9364 29850
rect 9312 29786 9364 29792
rect 9036 29504 9088 29510
rect 9036 29446 9088 29452
rect 7564 27940 7616 27946
rect 7564 27882 7616 27888
rect 7472 27056 7524 27062
rect 7472 26998 7524 27004
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8404 24274 8432 24686
rect 8392 24268 8444 24274
rect 8392 24210 8444 24216
rect 8772 23866 8800 24686
rect 8760 23860 8812 23866
rect 8760 23802 8812 23808
rect 8944 23724 8996 23730
rect 8944 23666 8996 23672
rect 8956 22642 8984 23666
rect 8944 22636 8996 22642
rect 8944 22578 8996 22584
rect 8956 22030 8984 22578
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8852 21956 8904 21962
rect 8852 21898 8904 21904
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8772 21622 8800 21830
rect 8760 21616 8812 21622
rect 8760 21558 8812 21564
rect 8864 21486 8892 21898
rect 8956 21622 8984 21966
rect 8944 21616 8996 21622
rect 8944 21558 8996 21564
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 9048 17610 9076 29446
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 9140 20874 9168 22374
rect 9128 20868 9180 20874
rect 9128 20810 9180 20816
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6748 2514 6776 2790
rect 6932 2582 6960 3878
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7944 3058 7972 3470
rect 8128 3126 8156 3878
rect 8864 3194 8892 4082
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7116 800 7144 2450
rect 7208 2310 7236 2450
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7760 800 7788 2926
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8496 1306 8524 2382
rect 8404 1278 8524 1306
rect 8404 800 8432 1278
rect 9048 800 9076 2790
rect 9324 2650 9352 29786
rect 9600 29170 9628 31758
rect 10704 31346 10732 31758
rect 12256 31748 12308 31754
rect 12256 31690 12308 31696
rect 12268 31346 12296 31690
rect 12452 31686 12480 31758
rect 12440 31680 12492 31686
rect 12440 31622 12492 31628
rect 10692 31340 10744 31346
rect 10692 31282 10744 31288
rect 10876 31340 10928 31346
rect 10876 31282 10928 31288
rect 12256 31340 12308 31346
rect 12256 31282 12308 31288
rect 10784 31136 10836 31142
rect 10784 31078 10836 31084
rect 10796 30802 10824 31078
rect 10784 30796 10836 30802
rect 10784 30738 10836 30744
rect 10600 30252 10652 30258
rect 10600 30194 10652 30200
rect 10692 30252 10744 30258
rect 10692 30194 10744 30200
rect 9680 29572 9732 29578
rect 9680 29514 9732 29520
rect 9692 29306 9720 29514
rect 9680 29300 9732 29306
rect 9680 29242 9732 29248
rect 9588 29164 9640 29170
rect 9588 29106 9640 29112
rect 9600 27470 9628 29106
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 10152 28558 10180 28902
rect 10612 28694 10640 30194
rect 10704 28966 10732 30194
rect 10692 28960 10744 28966
rect 10692 28902 10744 28908
rect 10888 28778 10916 31282
rect 12348 31136 12400 31142
rect 12348 31078 12400 31084
rect 12360 30666 12388 31078
rect 11060 30660 11112 30666
rect 11060 30602 11112 30608
rect 12348 30660 12400 30666
rect 12348 30602 12400 30608
rect 11072 30394 11100 30602
rect 11060 30388 11112 30394
rect 11060 30330 11112 30336
rect 12452 30258 12480 31622
rect 13004 30870 13032 32166
rect 13372 31822 13400 33390
rect 14004 32904 14056 32910
rect 14004 32846 14056 32852
rect 14016 32434 14044 32846
rect 14200 32502 14228 33390
rect 14188 32496 14240 32502
rect 14188 32438 14240 32444
rect 14004 32428 14056 32434
rect 14004 32370 14056 32376
rect 13544 32360 13596 32366
rect 13544 32302 13596 32308
rect 13176 31816 13228 31822
rect 13176 31758 13228 31764
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 12992 30864 13044 30870
rect 12992 30806 13044 30812
rect 12624 30592 12676 30598
rect 12624 30534 12676 30540
rect 12636 30394 12664 30534
rect 12624 30388 12676 30394
rect 12624 30330 12676 30336
rect 12716 30320 12768 30326
rect 12716 30262 12768 30268
rect 10968 30252 11020 30258
rect 10968 30194 11020 30200
rect 12440 30252 12492 30258
rect 12440 30194 12492 30200
rect 10980 29714 11008 30194
rect 12452 30054 12480 30194
rect 12440 30048 12492 30054
rect 12440 29990 12492 29996
rect 10968 29708 11020 29714
rect 10968 29650 11020 29656
rect 12728 28966 12756 30262
rect 13188 30258 13216 31758
rect 13372 30666 13400 31758
rect 13556 31686 13584 32302
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14568 31890 14596 32166
rect 14556 31884 14608 31890
rect 14556 31826 14608 31832
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14464 31816 14516 31822
rect 14464 31758 14516 31764
rect 13544 31680 13596 31686
rect 13544 31622 13596 31628
rect 14096 31680 14148 31686
rect 14096 31622 14148 31628
rect 13556 30734 13584 31622
rect 14108 31414 14136 31622
rect 14096 31408 14148 31414
rect 14096 31350 14148 31356
rect 14292 30802 14320 31758
rect 14280 30796 14332 30802
rect 14280 30738 14332 30744
rect 13544 30728 13596 30734
rect 13544 30670 13596 30676
rect 13360 30660 13412 30666
rect 13360 30602 13412 30608
rect 13372 30326 13400 30602
rect 14188 30592 14240 30598
rect 14188 30534 14240 30540
rect 13360 30320 13412 30326
rect 13360 30262 13412 30268
rect 14200 30258 14228 30534
rect 14292 30394 14320 30738
rect 14372 30728 14424 30734
rect 14372 30670 14424 30676
rect 14280 30388 14332 30394
rect 14280 30330 14332 30336
rect 13176 30252 13228 30258
rect 13176 30194 13228 30200
rect 14188 30252 14240 30258
rect 14188 30194 14240 30200
rect 13188 29238 13216 30194
rect 13176 29232 13228 29238
rect 13176 29174 13228 29180
rect 13544 29164 13596 29170
rect 13544 29106 13596 29112
rect 12716 28960 12768 28966
rect 12716 28902 12768 28908
rect 10796 28750 10916 28778
rect 10600 28688 10652 28694
rect 10600 28630 10652 28636
rect 10140 28552 10192 28558
rect 10140 28494 10192 28500
rect 10796 28014 10824 28750
rect 10876 28688 10928 28694
rect 10876 28630 10928 28636
rect 9680 28008 9732 28014
rect 9680 27950 9732 27956
rect 10784 28008 10836 28014
rect 10784 27950 10836 27956
rect 9692 27606 9720 27950
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9600 26858 9628 27406
rect 10796 26994 10824 27950
rect 10888 27452 10916 28630
rect 12728 28626 12756 28902
rect 12716 28620 12768 28626
rect 12716 28562 12768 28568
rect 10968 28552 11020 28558
rect 10968 28494 11020 28500
rect 10980 28150 11008 28494
rect 11980 28484 12032 28490
rect 11980 28426 12032 28432
rect 10968 28144 11020 28150
rect 10968 28086 11020 28092
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 10968 27464 11020 27470
rect 10888 27424 10968 27452
rect 10968 27406 11020 27412
rect 10876 27328 10928 27334
rect 10876 27270 10928 27276
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 9588 26852 9640 26858
rect 9588 26794 9640 26800
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10612 26450 10640 26726
rect 10888 26450 10916 27270
rect 10980 27130 11008 27406
rect 10968 27124 11020 27130
rect 10968 27066 11020 27072
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10600 26444 10652 26450
rect 10600 26386 10652 26392
rect 10876 26444 10928 26450
rect 10876 26386 10928 26392
rect 10980 25906 11008 26930
rect 11348 26586 11376 28018
rect 11992 27606 12020 28426
rect 13556 27878 13584 29106
rect 13636 29028 13688 29034
rect 13636 28970 13688 28976
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 11980 27600 12032 27606
rect 11980 27542 12032 27548
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 13360 27464 13412 27470
rect 13360 27406 13412 27412
rect 11520 27396 11572 27402
rect 11520 27338 11572 27344
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 11348 25906 11376 26522
rect 11428 25968 11480 25974
rect 11428 25910 11480 25916
rect 10968 25900 11020 25906
rect 10968 25842 11020 25848
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9692 25362 9720 25638
rect 10980 25430 11008 25842
rect 11440 25702 11468 25910
rect 11532 25770 11560 27338
rect 12636 26994 12664 27406
rect 12624 26988 12676 26994
rect 12624 26930 12676 26936
rect 11612 26784 11664 26790
rect 11612 26726 11664 26732
rect 11624 26314 11652 26726
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 12360 25974 12388 26522
rect 12348 25968 12400 25974
rect 12348 25910 12400 25916
rect 11888 25900 11940 25906
rect 11888 25842 11940 25848
rect 11520 25764 11572 25770
rect 11520 25706 11572 25712
rect 11428 25696 11480 25702
rect 11428 25638 11480 25644
rect 10968 25424 11020 25430
rect 10968 25366 11020 25372
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9956 25220 10008 25226
rect 9956 25162 10008 25168
rect 9968 24410 9996 25162
rect 10876 25152 10928 25158
rect 10876 25094 10928 25100
rect 10888 24886 10916 25094
rect 10876 24880 10928 24886
rect 10876 24822 10928 24828
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 10888 24274 10916 24822
rect 11440 24682 11468 25638
rect 11796 24744 11848 24750
rect 11796 24686 11848 24692
rect 11428 24676 11480 24682
rect 11428 24618 11480 24624
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 11440 24206 11468 24618
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 11624 24206 11652 24550
rect 11808 24410 11836 24686
rect 11900 24562 11928 25842
rect 12348 25356 12400 25362
rect 12348 25298 12400 25304
rect 11980 24608 12032 24614
rect 11900 24556 11980 24562
rect 11900 24550 12032 24556
rect 11900 24534 12020 24550
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 11808 24070 11836 24346
rect 11900 24206 11928 24534
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11072 23866 11100 24006
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9784 21894 9812 22578
rect 11072 22574 11100 23802
rect 11440 23594 11468 24006
rect 11428 23588 11480 23594
rect 11428 23530 11480 23536
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11716 23186 11744 23462
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11060 22568 11112 22574
rect 11060 22510 11112 22516
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10152 22234 10180 22374
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 10704 22098 10732 22374
rect 10692 22092 10744 22098
rect 10692 22034 10744 22040
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 11072 21894 11100 22034
rect 11348 21894 11376 22578
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 9784 20806 9812 21830
rect 11348 21554 11376 21830
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 10796 11014 10824 20810
rect 10980 20602 11008 21354
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 10980 19922 11008 20538
rect 11348 20466 11376 21490
rect 11440 21418 11468 23054
rect 11612 22432 11664 22438
rect 11612 22374 11664 22380
rect 11624 21962 11652 22374
rect 11808 22098 11836 24006
rect 11900 23866 11928 24142
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 12084 23186 12112 23258
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11612 21956 11664 21962
rect 11612 21898 11664 21904
rect 11428 21412 11480 21418
rect 11428 21354 11480 21360
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 11348 19378 11376 20402
rect 11796 20392 11848 20398
rect 11796 20334 11848 20340
rect 11808 19990 11836 20334
rect 11796 19984 11848 19990
rect 11796 19926 11848 19932
rect 11900 19854 11928 22510
rect 12360 22030 12388 25298
rect 12636 25294 12664 26930
rect 13372 26246 13400 27406
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 13372 25378 13400 26182
rect 13372 25350 13492 25378
rect 13464 25294 13492 25350
rect 13556 25294 13584 27814
rect 13648 27334 13676 28970
rect 14096 28688 14148 28694
rect 14096 28630 14148 28636
rect 14108 28218 14136 28630
rect 14200 28626 14228 30194
rect 14188 28620 14240 28626
rect 14188 28562 14240 28568
rect 14200 28218 14228 28562
rect 14384 28422 14412 30670
rect 14476 30190 14504 31758
rect 14568 31498 14596 31826
rect 14568 31482 14688 31498
rect 14568 31476 14700 31482
rect 14568 31470 14648 31476
rect 14648 31418 14700 31424
rect 14464 30184 14516 30190
rect 14464 30126 14516 30132
rect 14464 29232 14516 29238
rect 14464 29174 14516 29180
rect 14476 28762 14504 29174
rect 14752 28966 14780 46922
rect 15488 45554 15516 49200
rect 16500 47054 16528 49286
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49314 27150 50000
rect 26620 49286 27150 49314
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 16948 47048 17000 47054
rect 16948 46990 17000 46996
rect 15936 45620 15988 45626
rect 15936 45562 15988 45568
rect 15488 45526 15884 45554
rect 15856 33590 15884 45526
rect 15844 33584 15896 33590
rect 15844 33526 15896 33532
rect 15948 32978 15976 45562
rect 16960 33318 16988 46990
rect 17420 45626 17448 49200
rect 18708 47122 18736 49200
rect 19996 47122 20024 49200
rect 20536 47592 20588 47598
rect 20536 47534 20588 47540
rect 18696 47116 18748 47122
rect 18696 47058 18748 47064
rect 19984 47116 20036 47122
rect 19984 47058 20036 47064
rect 20352 47048 20404 47054
rect 20352 46990 20404 46996
rect 18696 46980 18748 46986
rect 18696 46922 18748 46928
rect 17408 45620 17460 45626
rect 17408 45562 17460 45568
rect 16948 33312 17000 33318
rect 16948 33254 17000 33260
rect 15936 32972 15988 32978
rect 15936 32914 15988 32920
rect 15108 32020 15160 32026
rect 15108 31962 15160 31968
rect 15120 31346 15148 31962
rect 16856 31748 16908 31754
rect 16856 31690 16908 31696
rect 16868 31346 16896 31690
rect 15108 31340 15160 31346
rect 15108 31282 15160 31288
rect 15292 31340 15344 31346
rect 15292 31282 15344 31288
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 15304 30258 15332 31282
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 15660 30728 15712 30734
rect 15660 30670 15712 30676
rect 15672 30394 15700 30670
rect 16684 30666 16712 31078
rect 16672 30660 16724 30666
rect 16672 30602 16724 30608
rect 15660 30388 15712 30394
rect 15660 30330 15712 30336
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15304 29646 15332 30194
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 15200 29164 15252 29170
rect 15200 29106 15252 29112
rect 14740 28960 14792 28966
rect 14740 28902 14792 28908
rect 14464 28756 14516 28762
rect 14464 28698 14516 28704
rect 15212 28558 15240 29106
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 14556 28484 14608 28490
rect 14556 28426 14608 28432
rect 14372 28416 14424 28422
rect 14372 28358 14424 28364
rect 14096 28212 14148 28218
rect 14096 28154 14148 28160
rect 14188 28212 14240 28218
rect 14188 28154 14240 28160
rect 14384 27946 14412 28358
rect 14568 28082 14596 28426
rect 14752 28082 14780 28494
rect 15304 28404 15332 29582
rect 15752 29572 15804 29578
rect 15752 29514 15804 29520
rect 15660 29164 15712 29170
rect 15660 29106 15712 29112
rect 15476 29096 15528 29102
rect 15476 29038 15528 29044
rect 15212 28376 15332 28404
rect 14556 28076 14608 28082
rect 14556 28018 14608 28024
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14372 27940 14424 27946
rect 14372 27882 14424 27888
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 13636 27328 13688 27334
rect 13636 27270 13688 27276
rect 13648 27130 13676 27270
rect 13636 27124 13688 27130
rect 13636 27066 13688 27072
rect 14108 26994 14136 27406
rect 13912 26988 13964 26994
rect 13912 26930 13964 26936
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 13268 25288 13320 25294
rect 13452 25288 13504 25294
rect 13320 25236 13400 25242
rect 13268 25230 13400 25236
rect 13452 25230 13504 25236
rect 13544 25288 13596 25294
rect 13544 25230 13596 25236
rect 13280 25214 13400 25230
rect 12624 24676 12676 24682
rect 12624 24618 12676 24624
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12452 23798 12480 24210
rect 12636 24138 12664 24618
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12440 23792 12492 23798
rect 12440 23734 12492 23740
rect 13096 23322 13124 24142
rect 13372 24070 13400 25214
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 12440 23044 12492 23050
rect 12440 22986 12492 22992
rect 12452 22778 12480 22986
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 13096 22094 13124 23258
rect 13372 22642 13400 24006
rect 13464 23118 13492 25230
rect 13556 24206 13584 25230
rect 13636 25152 13688 25158
rect 13636 25094 13688 25100
rect 13648 24886 13676 25094
rect 13636 24880 13688 24886
rect 13636 24822 13688 24828
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13176 22094 13228 22098
rect 13096 22092 13228 22094
rect 13096 22066 13176 22092
rect 13176 22034 13228 22040
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13372 21622 13400 21966
rect 13360 21616 13412 21622
rect 13360 21558 13412 21564
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 12820 19990 12848 20470
rect 13556 20398 13584 24142
rect 13648 23730 13676 24142
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 13832 23322 13860 23598
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 13924 22642 13952 26930
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 14200 26042 14228 26318
rect 14188 26036 14240 26042
rect 14188 25978 14240 25984
rect 14280 25968 14332 25974
rect 14280 25910 14332 25916
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 14200 25770 14228 25842
rect 14188 25764 14240 25770
rect 14188 25706 14240 25712
rect 14200 25226 14228 25706
rect 14292 25498 14320 25910
rect 14280 25492 14332 25498
rect 14280 25434 14332 25440
rect 14188 25220 14240 25226
rect 14188 25162 14240 25168
rect 14096 23656 14148 23662
rect 14096 23598 14148 23604
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 14016 22030 14044 22374
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 13636 21956 13688 21962
rect 13636 21898 13688 21904
rect 13648 21622 13676 21898
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 12808 19984 12860 19990
rect 12808 19926 12860 19932
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 12360 19378 12388 19858
rect 13096 19854 13124 20198
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11808 18834 11836 19110
rect 12084 18834 12112 19110
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 13004 18222 13032 18362
rect 13096 18290 13124 19790
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13740 19174 13768 19722
rect 13832 19446 13860 20538
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 14016 19718 14044 20402
rect 14108 20330 14136 23598
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14200 20602 14228 21422
rect 14292 20602 14320 25434
rect 14384 24750 14412 27882
rect 14568 26858 14596 28018
rect 14556 26852 14608 26858
rect 14556 26794 14608 26800
rect 14568 25702 14596 26794
rect 14752 26586 14780 28018
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 14936 26586 14964 26930
rect 15212 26926 15240 28376
rect 15488 28150 15516 29038
rect 15568 28484 15620 28490
rect 15568 28426 15620 28432
rect 15476 28144 15528 28150
rect 15476 28086 15528 28092
rect 15580 28082 15608 28426
rect 15568 28076 15620 28082
rect 15672 28064 15700 29106
rect 15764 29102 15792 29514
rect 16868 29170 16896 31282
rect 17132 30116 17184 30122
rect 17132 30058 17184 30064
rect 17144 29850 17172 30058
rect 17132 29844 17184 29850
rect 17132 29786 17184 29792
rect 16948 29572 17000 29578
rect 16948 29514 17000 29520
rect 16960 29306 16988 29514
rect 17868 29504 17920 29510
rect 17868 29446 17920 29452
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 15752 29096 15804 29102
rect 15752 29038 15804 29044
rect 16672 28620 16724 28626
rect 16672 28562 16724 28568
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 15948 28150 15976 28494
rect 16304 28484 16356 28490
rect 16304 28426 16356 28432
rect 16316 28218 16344 28426
rect 16304 28212 16356 28218
rect 16304 28154 16356 28160
rect 15936 28144 15988 28150
rect 15936 28086 15988 28092
rect 15752 28076 15804 28082
rect 15672 28036 15752 28064
rect 15568 28018 15620 28024
rect 15752 28018 15804 28024
rect 15764 27606 15792 28018
rect 15752 27600 15804 27606
rect 15752 27542 15804 27548
rect 15384 27328 15436 27334
rect 15384 27270 15436 27276
rect 15292 27124 15344 27130
rect 15292 27066 15344 27072
rect 15200 26920 15252 26926
rect 15200 26862 15252 26868
rect 14740 26580 14792 26586
rect 14740 26522 14792 26528
rect 14924 26580 14976 26586
rect 14924 26522 14976 26528
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14752 25906 14780 26318
rect 14936 25974 14964 26522
rect 14924 25968 14976 25974
rect 14924 25910 14976 25916
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 14556 25696 14608 25702
rect 14608 25656 14688 25684
rect 14556 25638 14608 25644
rect 14464 25152 14516 25158
rect 14464 25094 14516 25100
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14476 24682 14504 25094
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 14384 21622 14412 21830
rect 14372 21616 14424 21622
rect 14372 21558 14424 21564
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14096 20324 14148 20330
rect 14096 20266 14148 20272
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 14016 19446 14044 19654
rect 13820 19440 13872 19446
rect 13820 19382 13872 19388
rect 14004 19440 14056 19446
rect 14004 19382 14056 19388
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13832 18970 13860 19382
rect 14108 18970 14136 19722
rect 14476 19446 14504 20402
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18426 13216 18702
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13740 18222 13768 18838
rect 14292 18766 14320 19246
rect 14476 19174 14504 19382
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9416 3466 9444 3878
rect 9508 3602 9536 4558
rect 13740 4146 13768 18158
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 16658 14412 16934
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14568 13802 14596 24686
rect 14660 17746 14688 25656
rect 14752 25226 14780 25842
rect 15212 25498 15240 26862
rect 15304 26042 15332 27066
rect 15396 26994 15424 27270
rect 15948 27130 15976 28086
rect 16488 28076 16540 28082
rect 16488 28018 16540 28024
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 16408 26994 16436 27406
rect 16500 27334 16528 28018
rect 16684 27538 16712 28562
rect 17776 28552 17828 28558
rect 17776 28494 17828 28500
rect 17316 28484 17368 28490
rect 17316 28426 17368 28432
rect 16672 27532 16724 27538
rect 16672 27474 16724 27480
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 17328 27130 17356 28426
rect 17788 27470 17816 28494
rect 17880 27606 17908 29446
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 18064 28082 18092 28358
rect 18248 28150 18276 28358
rect 18236 28144 18288 28150
rect 18236 28086 18288 28092
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 17868 27600 17920 27606
rect 17868 27542 17920 27548
rect 17776 27464 17828 27470
rect 17776 27406 17828 27412
rect 17316 27124 17368 27130
rect 17316 27066 17368 27072
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16672 26988 16724 26994
rect 16672 26930 16724 26936
rect 15660 26784 15712 26790
rect 15660 26726 15712 26732
rect 15844 26784 15896 26790
rect 15844 26726 15896 26732
rect 15384 26308 15436 26314
rect 15384 26250 15436 26256
rect 15292 26036 15344 26042
rect 15292 25978 15344 25984
rect 15396 25498 15424 26250
rect 15200 25492 15252 25498
rect 15200 25434 15252 25440
rect 15384 25492 15436 25498
rect 15384 25434 15436 25440
rect 15672 25294 15700 26726
rect 15856 26450 15884 26726
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 16028 26308 16080 26314
rect 16028 26250 16080 26256
rect 16040 26042 16068 26250
rect 16028 26036 16080 26042
rect 16028 25978 16080 25984
rect 16684 25906 16712 26930
rect 17788 26246 17816 27406
rect 17880 26994 17908 27542
rect 18052 27328 18104 27334
rect 18052 27270 18104 27276
rect 18064 27062 18092 27270
rect 18052 27056 18104 27062
rect 18052 26998 18104 27004
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17776 26240 17828 26246
rect 17776 26182 17828 26188
rect 17788 26042 17816 26182
rect 17776 26036 17828 26042
rect 17776 25978 17828 25984
rect 16672 25900 16724 25906
rect 16672 25842 16724 25848
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 14740 25220 14792 25226
rect 14740 25162 14792 25168
rect 14752 18578 14780 25162
rect 15856 24342 15884 25230
rect 16684 25158 16712 25842
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 15844 24336 15896 24342
rect 15844 24278 15896 24284
rect 15384 24268 15436 24274
rect 15384 24210 15436 24216
rect 15200 24064 15252 24070
rect 15200 24006 15252 24012
rect 15108 23112 15160 23118
rect 15212 23066 15240 24006
rect 15160 23060 15240 23066
rect 15108 23054 15240 23060
rect 15120 23038 15240 23054
rect 15396 23050 15424 24210
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16592 23322 16620 24074
rect 16684 23730 16712 25094
rect 17040 24744 17092 24750
rect 17040 24686 17092 24692
rect 17052 24410 17080 24686
rect 17040 24404 17092 24410
rect 17040 24346 17092 24352
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16684 23118 16712 23666
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16776 23050 16804 23462
rect 15384 23044 15436 23050
rect 15384 22986 15436 22992
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16212 21956 16264 21962
rect 16212 21898 16264 21904
rect 16026 21584 16082 21593
rect 16026 21519 16028 21528
rect 16080 21519 16082 21528
rect 16028 21490 16080 21496
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14844 19446 14872 19654
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 14844 18766 14872 19382
rect 15028 18766 15056 19382
rect 15672 19378 15700 20198
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15764 19446 15792 19722
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 14752 18550 14872 18578
rect 14844 17814 14872 18550
rect 14832 17808 14884 17814
rect 14832 17750 14884 17756
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14844 17678 14872 17750
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 15028 17542 15056 18702
rect 15120 18630 15148 19110
rect 15108 18624 15160 18630
rect 15108 18566 15160 18572
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14660 16046 14688 16458
rect 14936 16114 14964 17070
rect 15028 16182 15056 17478
rect 15120 16250 15148 18566
rect 15672 17202 15700 19314
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15396 16522 15424 16934
rect 15672 16658 15700 17138
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 14648 16040 14700 16046
rect 16040 15994 16068 16050
rect 14648 15982 14700 15988
rect 15948 15966 16068 15994
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 14936 15570 14964 15846
rect 15212 15570 15240 15846
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15948 15366 15976 15966
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15948 14482 15976 15302
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16132 14482 16160 14758
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 14556 13796 14608 13802
rect 14556 13738 14608 13744
rect 14832 13456 14884 13462
rect 14832 13398 14884 13404
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 9600 2854 9628 3538
rect 11532 3058 11560 3878
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11716 3126 11744 3334
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 13832 3058 13860 3470
rect 14016 3126 14044 3878
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 10980 800 11008 2926
rect 14200 800 14228 2926
rect 14844 800 14872 13398
rect 16224 6914 16252 21898
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16316 18290 16344 19654
rect 16592 19378 16620 22578
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16684 21418 16712 22510
rect 16868 21894 16896 24142
rect 17236 22710 17264 25842
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 17972 24886 18000 25094
rect 17960 24880 18012 24886
rect 17960 24822 18012 24828
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 17684 24064 17736 24070
rect 17684 24006 17736 24012
rect 17696 23730 17724 24006
rect 18064 23866 18092 24686
rect 18144 24336 18196 24342
rect 18144 24278 18196 24284
rect 18052 23860 18104 23866
rect 18052 23802 18104 23808
rect 18156 23730 18184 24278
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 17500 22976 17552 22982
rect 17500 22918 17552 22924
rect 17512 22710 17540 22918
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 17224 22704 17276 22710
rect 17224 22646 17276 22652
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 16948 22568 17000 22574
rect 16948 22510 17000 22516
rect 16960 22234 16988 22510
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 17972 22030 18000 22714
rect 18156 22658 18184 23666
rect 18236 22704 18288 22710
rect 18156 22652 18236 22658
rect 18156 22646 18288 22652
rect 18156 22630 18276 22646
rect 18156 22098 18184 22630
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 18524 22030 18552 22374
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 16868 21554 16896 21830
rect 18156 21622 18184 21830
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16672 21412 16724 21418
rect 16672 21354 16724 21360
rect 16868 20942 16896 21490
rect 17224 21480 17276 21486
rect 17224 21422 17276 21428
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 17052 21146 17080 21286
rect 17236 21146 17264 21422
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 16856 20936 16908 20942
rect 16856 20878 16908 20884
rect 16868 20466 16896 20878
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 16868 19922 16896 20198
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 18156 19786 18184 20198
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18144 19780 18196 19786
rect 18144 19722 18196 19728
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16592 18766 16620 19314
rect 18340 19310 18368 19858
rect 18616 19718 18644 20198
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17144 17882 17172 18158
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17328 17678 17356 18566
rect 18524 17678 18552 19382
rect 18616 19378 18644 19654
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16592 16250 16620 16458
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16592 12850 16620 16186
rect 16960 15502 16988 16390
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 17328 15026 17356 17614
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17604 15366 17632 16594
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17880 15994 17908 16118
rect 17972 16114 18000 16934
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 18156 15994 18184 16526
rect 18248 16182 18276 16594
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 17788 15706 17816 15982
rect 17880 15966 18184 15994
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17972 15434 18000 15846
rect 18156 15638 18184 15966
rect 18144 15632 18196 15638
rect 18144 15574 18196 15580
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17972 15026 18000 15370
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 16776 13938 16804 14962
rect 17972 14822 18000 14962
rect 18156 14958 18184 15302
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 16776 13394 16804 13670
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16960 12918 16988 13670
rect 17972 13258 18000 14758
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16132 6886 16252 6914
rect 16132 3466 16160 6886
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17236 4010 17264 4218
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17512 3534 17540 3878
rect 17500 3528 17552 3534
rect 17776 3528 17828 3534
rect 17500 3470 17552 3476
rect 17590 3496 17646 3505
rect 16120 3460 16172 3466
rect 17776 3470 17828 3476
rect 17590 3431 17646 3440
rect 16120 3402 16172 3408
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15212 2650 15240 2926
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15488 800 15516 2314
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15764 1902 15792 2246
rect 15752 1896 15804 1902
rect 15752 1838 15804 1844
rect 16132 800 16160 2382
rect 17328 2310 17356 2586
rect 17420 2446 17448 3334
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17604 1034 17632 3431
rect 17788 3126 17816 3470
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17972 2650 18000 4082
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18064 2446 18092 4966
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18156 4214 18184 4422
rect 18144 4208 18196 4214
rect 18144 4150 18196 4156
rect 18248 3738 18276 4558
rect 18340 4078 18368 5170
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18524 4010 18552 17614
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18616 15502 18644 15846
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18616 13938 18644 15438
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18616 8294 18644 12718
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 18156 3398 18184 3606
rect 18236 3460 18288 3466
rect 18340 3448 18368 3606
rect 18616 3482 18644 3946
rect 18708 3738 18736 46922
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19432 46504 19484 46510
rect 19432 46446 19484 46452
rect 20260 46504 20312 46510
rect 20260 46446 20312 46452
rect 19444 46170 19472 46446
rect 19432 46164 19484 46170
rect 19432 46106 19484 46112
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 20272 45626 20300 46446
rect 20260 45620 20312 45626
rect 20260 45562 20312 45568
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 20260 35080 20312 35086
rect 20260 35022 20312 35028
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 20076 34060 20128 34066
rect 20076 34002 20128 34008
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 20088 33590 20116 34002
rect 20076 33584 20128 33590
rect 20076 33526 20128 33532
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 18880 31272 18932 31278
rect 18880 31214 18932 31220
rect 18892 30802 18920 31214
rect 20088 30802 20116 33526
rect 20168 31816 20220 31822
rect 20168 31758 20220 31764
rect 20180 31414 20208 31758
rect 20168 31408 20220 31414
rect 20168 31350 20220 31356
rect 18880 30796 18932 30802
rect 18880 30738 18932 30744
rect 20076 30796 20128 30802
rect 20076 30738 20128 30744
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19432 28484 19484 28490
rect 19432 28426 19484 28432
rect 19248 27124 19300 27130
rect 19248 27066 19300 27072
rect 19260 25770 19288 27066
rect 19444 26450 19472 28426
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 20272 28082 20300 35022
rect 20364 32502 20392 46990
rect 20548 35630 20576 47534
rect 20640 46510 20668 49200
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 20812 46368 20864 46374
rect 20812 46310 20864 46316
rect 20824 46034 20852 46310
rect 21284 46034 21312 49200
rect 24860 47048 24912 47054
rect 24860 46990 24912 46996
rect 24872 46646 24900 46990
rect 24860 46640 24912 46646
rect 24860 46582 24912 46588
rect 25148 46510 25176 49200
rect 25504 47048 25556 47054
rect 25504 46990 25556 46996
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 25136 46504 25188 46510
rect 25136 46446 25188 46452
rect 24780 46170 24808 46446
rect 24768 46164 24820 46170
rect 24768 46106 24820 46112
rect 25516 46034 25544 46990
rect 20812 46028 20864 46034
rect 20812 45970 20864 45976
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 25504 46028 25556 46034
rect 25504 45970 25556 45976
rect 24860 45960 24912 45966
rect 24860 45902 24912 45908
rect 20996 45892 21048 45898
rect 20996 45834 21048 45840
rect 21008 45626 21036 45834
rect 20996 45620 21048 45626
rect 20996 45562 21048 45568
rect 24872 45490 24900 45902
rect 25412 45892 25464 45898
rect 25412 45834 25464 45840
rect 25424 45626 25452 45834
rect 25792 45830 25820 49200
rect 25780 45824 25832 45830
rect 25780 45766 25832 45772
rect 25412 45620 25464 45626
rect 25412 45562 25464 45568
rect 26620 45554 26648 49286
rect 27038 49200 27150 49286
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49200 31014 50000
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49200 40030 50000
rect 40562 49200 40674 50000
rect 41206 49314 41318 50000
rect 40788 49286 41318 49314
rect 28368 47054 28396 49200
rect 29000 47184 29052 47190
rect 29000 47126 29052 47132
rect 28908 47116 28960 47122
rect 28908 47058 28960 47064
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 28722 47016 28778 47025
rect 28722 46951 28724 46960
rect 28776 46951 28778 46960
rect 28724 46922 28776 46928
rect 27344 45824 27396 45830
rect 27344 45766 27396 45772
rect 26344 45526 26648 45554
rect 20812 45484 20864 45490
rect 20812 45426 20864 45432
rect 24860 45484 24912 45490
rect 24860 45426 24912 45432
rect 25320 45484 25372 45490
rect 25320 45426 25372 45432
rect 20824 41414 20852 45426
rect 20732 41386 20852 41414
rect 20732 37806 20760 41386
rect 20720 37800 20772 37806
rect 20720 37742 20772 37748
rect 20536 35624 20588 35630
rect 20536 35566 20588 35572
rect 20548 35086 20576 35566
rect 20536 35080 20588 35086
rect 20536 35022 20588 35028
rect 20536 33856 20588 33862
rect 20536 33798 20588 33804
rect 20548 33590 20576 33798
rect 20536 33584 20588 33590
rect 20536 33526 20588 33532
rect 20352 32496 20404 32502
rect 20352 32438 20404 32444
rect 20628 31272 20680 31278
rect 20628 31214 20680 31220
rect 20640 30326 20668 31214
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20536 30184 20588 30190
rect 20536 30126 20588 30132
rect 20548 29850 20576 30126
rect 20536 29844 20588 29850
rect 20536 29786 20588 29792
rect 20536 28484 20588 28490
rect 20536 28426 20588 28432
rect 20548 28218 20576 28426
rect 20536 28212 20588 28218
rect 20536 28154 20588 28160
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 20640 27062 20668 28018
rect 20628 27056 20680 27062
rect 20628 26998 20680 27004
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 20626 26888 20682 26897
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19248 25764 19300 25770
rect 19248 25706 19300 25712
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 19616 24744 19668 24750
rect 19616 24686 19668 24692
rect 18788 24268 18840 24274
rect 18788 24210 18840 24216
rect 18800 23798 18828 24210
rect 18984 24138 19012 24686
rect 19628 24410 19656 24686
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 18972 24132 19024 24138
rect 18972 24074 19024 24080
rect 18984 23866 19012 24074
rect 19076 23866 19104 24346
rect 19892 24200 19944 24206
rect 19944 24160 20024 24188
rect 19892 24142 19944 24148
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 18972 23860 19024 23866
rect 18972 23802 19024 23808
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 18788 23792 18840 23798
rect 18788 23734 18840 23740
rect 18800 22642 18828 23734
rect 19996 23730 20024 24160
rect 18880 23724 18932 23730
rect 18880 23666 18932 23672
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 18892 22778 18920 23666
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19444 23118 19472 23462
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 19156 22772 19208 22778
rect 19156 22714 19208 22720
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18800 21486 18828 22578
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 19076 19446 19104 22510
rect 19064 19440 19116 19446
rect 19064 19382 19116 19388
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18800 16522 18828 18158
rect 19168 17678 19196 22714
rect 19352 22030 19380 22918
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19996 22574 20024 23666
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19260 21146 19288 21490
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19260 20466 19288 20878
rect 19352 20602 19380 21966
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19260 19718 19288 20402
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19352 19242 19380 20538
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19444 19378 19472 19858
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19996 19446 20024 19790
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 18788 16516 18840 16522
rect 18788 16458 18840 16464
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19352 16114 19380 16390
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19812 15502 19840 16050
rect 19996 15502 20024 16594
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 15042 19472 15302
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19444 15014 19564 15042
rect 19536 14958 19564 15014
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18616 3454 18736 3482
rect 18288 3420 18368 3448
rect 18236 3402 18288 3408
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 17420 1006 17632 1034
rect 17420 800 17448 1006
rect 18708 800 18736 3454
rect 18800 3058 18828 3878
rect 18984 3466 19012 4082
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 19076 3126 19104 4082
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 19260 2650 19288 4558
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19352 3534 19380 4422
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 20088 3942 20116 26862
rect 20626 26823 20682 26832
rect 20640 26790 20668 26823
rect 20628 26784 20680 26790
rect 20628 26726 20680 26732
rect 20536 25696 20588 25702
rect 20536 25638 20588 25644
rect 20548 25362 20576 25638
rect 20536 25356 20588 25362
rect 20536 25298 20588 25304
rect 20168 24132 20220 24138
rect 20168 24074 20220 24080
rect 20180 23866 20208 24074
rect 20548 24070 20576 25298
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 20548 23118 20576 24006
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20272 19310 20300 20198
rect 20732 19938 20760 37742
rect 25332 36854 25360 45426
rect 26344 41414 26372 45526
rect 26344 41386 26464 41414
rect 25780 37120 25832 37126
rect 25780 37062 25832 37068
rect 25320 36848 25372 36854
rect 25320 36790 25372 36796
rect 25688 36780 25740 36786
rect 25688 36722 25740 36728
rect 22376 36576 22428 36582
rect 22376 36518 22428 36524
rect 22388 36106 22416 36518
rect 24400 36168 24452 36174
rect 24400 36110 24452 36116
rect 22376 36100 22428 36106
rect 22376 36042 22428 36048
rect 22836 36100 22888 36106
rect 22836 36042 22888 36048
rect 22848 35834 22876 36042
rect 22836 35828 22888 35834
rect 22836 35770 22888 35776
rect 22376 35760 22428 35766
rect 22376 35702 22428 35708
rect 22008 35692 22060 35698
rect 22008 35634 22060 35640
rect 20812 34944 20864 34950
rect 20812 34886 20864 34892
rect 20824 34610 20852 34886
rect 22020 34610 22048 35634
rect 20812 34604 20864 34610
rect 20812 34546 20864 34552
rect 22008 34604 22060 34610
rect 22008 34546 22060 34552
rect 20824 33998 20852 34546
rect 22192 34536 22244 34542
rect 22192 34478 22244 34484
rect 20812 33992 20864 33998
rect 20812 33934 20864 33940
rect 20824 31890 20852 33934
rect 22204 33930 22232 34478
rect 21640 33924 21692 33930
rect 21640 33866 21692 33872
rect 22192 33924 22244 33930
rect 22192 33866 22244 33872
rect 21652 33658 21680 33866
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 22192 33584 22244 33590
rect 22192 33526 22244 33532
rect 21916 33516 21968 33522
rect 21836 33476 21916 33504
rect 20996 33448 21048 33454
rect 20996 33390 21048 33396
rect 21008 33114 21036 33390
rect 21088 33312 21140 33318
rect 21088 33254 21140 33260
rect 20996 33108 21048 33114
rect 20996 33050 21048 33056
rect 21100 32910 21128 33254
rect 21548 32972 21600 32978
rect 21548 32914 21600 32920
rect 21088 32904 21140 32910
rect 21088 32846 21140 32852
rect 21272 32904 21324 32910
rect 21272 32846 21324 32852
rect 21100 32026 21128 32846
rect 21284 32502 21312 32846
rect 21272 32496 21324 32502
rect 21272 32438 21324 32444
rect 21456 32496 21508 32502
rect 21456 32438 21508 32444
rect 21088 32020 21140 32026
rect 21088 31962 21140 31968
rect 21468 31890 21496 32438
rect 20812 31884 20864 31890
rect 20812 31826 20864 31832
rect 21456 31884 21508 31890
rect 21456 31826 21508 31832
rect 20824 31346 20852 31826
rect 21364 31816 21416 31822
rect 21364 31758 21416 31764
rect 20904 31476 20956 31482
rect 20904 31418 20956 31424
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 20916 30258 20944 31418
rect 21272 31340 21324 31346
rect 21272 31282 21324 31288
rect 21180 31136 21232 31142
rect 21180 31078 21232 31084
rect 21192 30734 21220 31078
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 21088 28960 21140 28966
rect 21088 28902 21140 28908
rect 20996 28552 21048 28558
rect 20996 28494 21048 28500
rect 21008 27962 21036 28494
rect 21100 28082 21128 28902
rect 21180 28484 21232 28490
rect 21180 28426 21232 28432
rect 21192 28218 21220 28426
rect 21180 28212 21232 28218
rect 21180 28154 21232 28160
rect 21088 28076 21140 28082
rect 21088 28018 21140 28024
rect 21008 27934 21128 27962
rect 20996 27532 21048 27538
rect 20996 27474 21048 27480
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20916 26994 20944 27270
rect 20904 26988 20956 26994
rect 20904 26930 20956 26936
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20824 26314 20852 26726
rect 20812 26308 20864 26314
rect 20812 26250 20864 26256
rect 21008 25906 21036 27474
rect 21100 27470 21128 27934
rect 21192 27674 21220 28154
rect 21180 27668 21232 27674
rect 21180 27610 21232 27616
rect 21284 27470 21312 31282
rect 21376 30938 21404 31758
rect 21468 31482 21496 31826
rect 21456 31476 21508 31482
rect 21456 31418 21508 31424
rect 21364 30932 21416 30938
rect 21364 30874 21416 30880
rect 21376 30818 21404 30874
rect 21560 30870 21588 32914
rect 21732 32428 21784 32434
rect 21732 32370 21784 32376
rect 21640 31680 21692 31686
rect 21640 31622 21692 31628
rect 21548 30864 21600 30870
rect 21376 30790 21496 30818
rect 21548 30806 21600 30812
rect 21364 30660 21416 30666
rect 21364 30602 21416 30608
rect 21376 30122 21404 30602
rect 21468 30394 21496 30790
rect 21456 30388 21508 30394
rect 21456 30330 21508 30336
rect 21364 30116 21416 30122
rect 21364 30058 21416 30064
rect 21560 29850 21588 30806
rect 21548 29844 21600 29850
rect 21548 29786 21600 29792
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 21364 28416 21416 28422
rect 21364 28358 21416 28364
rect 21376 28218 21404 28358
rect 21364 28212 21416 28218
rect 21364 28154 21416 28160
rect 21376 28082 21404 28154
rect 21364 28076 21416 28082
rect 21364 28018 21416 28024
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21100 26314 21128 27406
rect 21088 26308 21140 26314
rect 21088 26250 21140 26256
rect 21284 25906 21312 27406
rect 21364 27396 21416 27402
rect 21364 27338 21416 27344
rect 21376 26314 21404 27338
rect 21364 26308 21416 26314
rect 21364 26250 21416 26256
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 21272 25900 21324 25906
rect 21272 25842 21324 25848
rect 21376 25838 21404 26250
rect 21364 25832 21416 25838
rect 21364 25774 21416 25780
rect 21272 24880 21324 24886
rect 21270 24848 21272 24857
rect 21324 24848 21326 24857
rect 21270 24783 21326 24792
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20916 22710 20944 23054
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 21192 22778 21220 22986
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 20904 22704 20956 22710
rect 20904 22646 20956 22652
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 21008 22098 21036 22374
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 20824 20466 20852 21966
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20916 21554 20944 21830
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20916 20942 20944 21286
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20916 20074 20944 20878
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 20916 20046 21036 20074
rect 20732 19910 20944 19938
rect 21008 19922 21036 20046
rect 20536 19780 20588 19786
rect 20536 19722 20588 19728
rect 20548 19310 20576 19722
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20272 18834 20300 19246
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18902 20760 19110
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20824 18426 20852 18702
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20444 17060 20496 17066
rect 20444 17002 20496 17008
rect 20456 16114 20484 17002
rect 20916 16574 20944 19910
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 21008 18290 21036 19858
rect 21192 19378 21220 20402
rect 21284 19378 21312 20538
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21008 17678 21036 18226
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17270 21036 17614
rect 21088 17604 21140 17610
rect 21088 17546 21140 17552
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 20732 16546 20944 16574
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 20180 15094 20208 15302
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20272 3738 20300 4082
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20180 3618 20208 3674
rect 20180 3590 20576 3618
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19708 3120 19760 3126
rect 19536 3080 19708 3108
rect 19536 2972 19564 3080
rect 19996 3074 20024 3334
rect 19708 3062 19760 3068
rect 19352 2944 19564 2972
rect 19904 3046 20024 3074
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19352 800 19380 2944
rect 19904 2922 19932 3046
rect 20364 2990 20392 3470
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20548 2922 20576 3590
rect 20640 3398 20668 13806
rect 20732 3466 20760 16546
rect 21008 16250 21036 17070
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20916 15570 20944 15846
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 21008 4282 21036 4490
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20824 3534 20852 3946
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20916 3534 20944 3878
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 21100 3126 21128 17546
rect 21468 6914 21496 29446
rect 21652 29238 21680 31622
rect 21744 31482 21772 32370
rect 21732 31476 21784 31482
rect 21732 31418 21784 31424
rect 21732 31136 21784 31142
rect 21732 31078 21784 31084
rect 21744 30258 21772 31078
rect 21836 30326 21864 33476
rect 21916 33458 21968 33464
rect 22204 33318 22232 33526
rect 22388 33522 22416 35702
rect 23480 34536 23532 34542
rect 23480 34478 23532 34484
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 23492 34406 23520 34478
rect 23480 34400 23532 34406
rect 23480 34342 23532 34348
rect 23492 34066 23520 34342
rect 23480 34060 23532 34066
rect 23480 34002 23532 34008
rect 22376 33516 22428 33522
rect 22376 33458 22428 33464
rect 22836 33516 22888 33522
rect 22836 33458 22888 33464
rect 22376 33380 22428 33386
rect 22376 33322 22428 33328
rect 22192 33312 22244 33318
rect 22192 33254 22244 33260
rect 22008 32972 22060 32978
rect 22008 32914 22060 32920
rect 22020 32484 22048 32914
rect 22388 32910 22416 33322
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 22560 32904 22612 32910
rect 22560 32846 22612 32852
rect 22100 32496 22152 32502
rect 22020 32456 22100 32484
rect 22100 32438 22152 32444
rect 21916 32428 21968 32434
rect 21916 32370 21968 32376
rect 21928 32314 21956 32370
rect 21928 32286 22140 32314
rect 22112 31890 22140 32286
rect 22284 32292 22336 32298
rect 22284 32234 22336 32240
rect 22100 31884 22152 31890
rect 22100 31826 22152 31832
rect 22296 31346 22324 32234
rect 22572 32230 22600 32846
rect 22744 32768 22796 32774
rect 22744 32710 22796 32716
rect 22560 32224 22612 32230
rect 22560 32166 22612 32172
rect 22572 32026 22600 32166
rect 22756 32026 22784 32710
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22744 32020 22796 32026
rect 22744 31962 22796 31968
rect 22560 31884 22612 31890
rect 22560 31826 22612 31832
rect 22572 31754 22600 31826
rect 22744 31816 22796 31822
rect 22744 31758 22796 31764
rect 22480 31726 22600 31754
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22480 31278 22508 31726
rect 22468 31272 22520 31278
rect 22468 31214 22520 31220
rect 22284 31204 22336 31210
rect 22284 31146 22336 31152
rect 22296 30734 22324 31146
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22376 30728 22428 30734
rect 22376 30670 22428 30676
rect 21916 30592 21968 30598
rect 21916 30534 21968 30540
rect 21824 30320 21876 30326
rect 21824 30262 21876 30268
rect 21928 30258 21956 30534
rect 22388 30394 22416 30670
rect 22376 30388 22428 30394
rect 22376 30330 22428 30336
rect 22388 30258 22416 30330
rect 21732 30252 21784 30258
rect 21732 30194 21784 30200
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 22376 30252 22428 30258
rect 22376 30194 22428 30200
rect 22284 30184 22336 30190
rect 22204 30144 22284 30172
rect 22100 29640 22152 29646
rect 22100 29582 22152 29588
rect 21640 29232 21692 29238
rect 21640 29174 21692 29180
rect 21652 28778 21680 29174
rect 21824 29028 21876 29034
rect 21824 28970 21876 28976
rect 21560 28750 21680 28778
rect 21560 27674 21588 28750
rect 21730 28656 21786 28665
rect 21640 28620 21692 28626
rect 21730 28591 21786 28600
rect 21640 28562 21692 28568
rect 21652 28150 21680 28562
rect 21744 28490 21772 28591
rect 21836 28558 21864 28970
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21732 28484 21784 28490
rect 21732 28426 21784 28432
rect 21640 28144 21692 28150
rect 21640 28086 21692 28092
rect 21548 27668 21600 27674
rect 21548 27610 21600 27616
rect 21560 25770 21588 27610
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21652 26450 21680 27270
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21548 25764 21600 25770
rect 21548 25706 21600 25712
rect 21744 25158 21772 28426
rect 22008 28416 22060 28422
rect 22008 28358 22060 28364
rect 22020 28082 22048 28358
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 22112 27418 22140 29582
rect 22020 27390 22140 27418
rect 21824 27328 21876 27334
rect 21824 27270 21876 27276
rect 21836 27130 21864 27270
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 22020 26994 22048 27390
rect 22100 27328 22152 27334
rect 22100 27270 22152 27276
rect 22112 26994 22140 27270
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 22112 26602 22140 26930
rect 22020 26574 22140 26602
rect 21916 26444 21968 26450
rect 21916 26386 21968 26392
rect 21928 26314 21956 26386
rect 22020 26382 22048 26574
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 21916 26308 21968 26314
rect 21916 26250 21968 26256
rect 21732 25152 21784 25158
rect 21732 25094 21784 25100
rect 21822 24168 21878 24177
rect 21822 24103 21824 24112
rect 21876 24103 21878 24112
rect 21824 24074 21876 24080
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22204 22930 22232 30144
rect 22284 30126 22336 30132
rect 22480 29170 22508 31214
rect 22756 31210 22784 31758
rect 22744 31204 22796 31210
rect 22744 31146 22796 31152
rect 22560 30660 22612 30666
rect 22560 30602 22612 30608
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22572 28966 22600 30602
rect 22652 30252 22704 30258
rect 22848 30240 22876 33458
rect 22928 33312 22980 33318
rect 22928 33254 22980 33260
rect 22940 32026 22968 33254
rect 23388 32224 23440 32230
rect 23388 32166 23440 32172
rect 22928 32020 22980 32026
rect 22928 31962 22980 31968
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 22704 30212 22876 30240
rect 22652 30194 22704 30200
rect 22560 28960 22612 28966
rect 22560 28902 22612 28908
rect 22572 28490 22600 28902
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22296 28082 22324 28358
rect 22376 28212 22428 28218
rect 22376 28154 22428 28160
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22388 27470 22416 28154
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 22664 26994 22692 30194
rect 22940 28694 22968 31282
rect 23400 30734 23428 32166
rect 23492 31414 23520 34002
rect 23572 33856 23624 33862
rect 23572 33798 23624 33804
rect 23584 33590 23612 33798
rect 23768 33658 23796 34478
rect 24412 34406 24440 36110
rect 24952 36100 25004 36106
rect 24952 36042 25004 36048
rect 25136 36100 25188 36106
rect 25136 36042 25188 36048
rect 24964 35834 24992 36042
rect 24952 35828 25004 35834
rect 24952 35770 25004 35776
rect 24584 35488 24636 35494
rect 24584 35430 24636 35436
rect 24596 35086 24624 35430
rect 25148 35290 25176 36042
rect 25700 36038 25728 36722
rect 25688 36032 25740 36038
rect 25688 35974 25740 35980
rect 25596 35556 25648 35562
rect 25596 35498 25648 35504
rect 25136 35284 25188 35290
rect 25136 35226 25188 35232
rect 24584 35080 24636 35086
rect 24584 35022 24636 35028
rect 25320 35080 25372 35086
rect 25320 35022 25372 35028
rect 25412 35080 25464 35086
rect 25412 35022 25464 35028
rect 24400 34400 24452 34406
rect 24400 34342 24452 34348
rect 24596 33998 24624 35022
rect 25136 35012 25188 35018
rect 25136 34954 25188 34960
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 24872 34202 24900 34546
rect 24860 34196 24912 34202
rect 24860 34138 24912 34144
rect 24584 33992 24636 33998
rect 24584 33934 24636 33940
rect 24768 33924 24820 33930
rect 24768 33866 24820 33872
rect 24676 33856 24728 33862
rect 24676 33798 24728 33804
rect 23756 33652 23808 33658
rect 23756 33594 23808 33600
rect 23572 33584 23624 33590
rect 23572 33526 23624 33532
rect 24124 33448 24176 33454
rect 24124 33390 24176 33396
rect 24688 33402 24716 33798
rect 24780 33522 24808 33866
rect 24768 33516 24820 33522
rect 24768 33458 24820 33464
rect 23480 31408 23532 31414
rect 23480 31350 23532 31356
rect 23388 30728 23440 30734
rect 23388 30670 23440 30676
rect 23020 30320 23072 30326
rect 23020 30262 23072 30268
rect 23032 29782 23060 30262
rect 24136 30122 24164 33390
rect 24688 33374 24808 33402
rect 24584 32972 24636 32978
rect 24584 32914 24636 32920
rect 24596 32026 24624 32914
rect 24780 32910 24808 33374
rect 25044 33312 25096 33318
rect 25044 33254 25096 33260
rect 25056 33114 25084 33254
rect 25044 33108 25096 33114
rect 25044 33050 25096 33056
rect 24768 32904 24820 32910
rect 24768 32846 24820 32852
rect 24780 32434 24808 32846
rect 25056 32502 25084 33050
rect 25044 32496 25096 32502
rect 25044 32438 25096 32444
rect 24768 32428 24820 32434
rect 24768 32370 24820 32376
rect 24584 32020 24636 32026
rect 24584 31962 24636 31968
rect 24492 31680 24544 31686
rect 24492 31622 24544 31628
rect 24504 31278 24532 31622
rect 24492 31272 24544 31278
rect 24492 31214 24544 31220
rect 24216 30252 24268 30258
rect 24216 30194 24268 30200
rect 24124 30116 24176 30122
rect 24124 30058 24176 30064
rect 23020 29776 23072 29782
rect 23020 29718 23072 29724
rect 24228 29578 24256 30194
rect 24216 29572 24268 29578
rect 24216 29514 24268 29520
rect 24492 29572 24544 29578
rect 24492 29514 24544 29520
rect 23296 29164 23348 29170
rect 23296 29106 23348 29112
rect 22744 28688 22796 28694
rect 22744 28630 22796 28636
rect 22928 28688 22980 28694
rect 22928 28630 22980 28636
rect 22756 28558 22784 28630
rect 22744 28552 22796 28558
rect 22744 28494 22796 28500
rect 23112 27872 23164 27878
rect 23112 27814 23164 27820
rect 23124 27062 23152 27814
rect 23308 27538 23336 29106
rect 24216 27600 24268 27606
rect 24216 27542 24268 27548
rect 23296 27532 23348 27538
rect 23296 27474 23348 27480
rect 23112 27056 23164 27062
rect 23112 26998 23164 27004
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22572 26586 22600 26726
rect 22560 26580 22612 26586
rect 22560 26522 22612 26528
rect 22284 26512 22336 26518
rect 22284 26454 22336 26460
rect 22296 25226 22324 26454
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22388 25362 22416 25638
rect 23124 25514 23152 26998
rect 24228 26858 24256 27542
rect 24504 27130 24532 29514
rect 24596 28558 24624 31962
rect 25044 31952 25096 31958
rect 25044 31894 25096 31900
rect 25056 31822 25084 31894
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 25148 31754 25176 34954
rect 25228 34536 25280 34542
rect 25228 34478 25280 34484
rect 25240 33454 25268 34478
rect 25332 33998 25360 35022
rect 25424 34542 25452 35022
rect 25412 34536 25464 34542
rect 25412 34478 25464 34484
rect 25608 34134 25636 35498
rect 25700 34746 25728 35974
rect 25792 35630 25820 37062
rect 26332 36712 26384 36718
rect 26332 36654 26384 36660
rect 26148 36032 26200 36038
rect 26148 35974 26200 35980
rect 26160 35766 26188 35974
rect 26148 35760 26200 35766
rect 26148 35702 26200 35708
rect 25780 35624 25832 35630
rect 25780 35566 25832 35572
rect 25792 35086 25820 35566
rect 25872 35488 25924 35494
rect 26056 35488 26108 35494
rect 25924 35436 26056 35442
rect 25872 35430 26108 35436
rect 25884 35414 26096 35430
rect 26160 35154 26188 35702
rect 26240 35624 26292 35630
rect 26240 35566 26292 35572
rect 26252 35290 26280 35566
rect 26344 35290 26372 36654
rect 26240 35284 26292 35290
rect 26240 35226 26292 35232
rect 26332 35284 26384 35290
rect 26332 35226 26384 35232
rect 25964 35148 26016 35154
rect 25964 35090 26016 35096
rect 26148 35148 26200 35154
rect 26148 35090 26200 35096
rect 25780 35080 25832 35086
rect 25780 35022 25832 35028
rect 25688 34740 25740 34746
rect 25688 34682 25740 34688
rect 25780 34536 25832 34542
rect 25780 34478 25832 34484
rect 25596 34128 25648 34134
rect 25596 34070 25648 34076
rect 25792 34066 25820 34478
rect 25976 34406 26004 35090
rect 25964 34400 26016 34406
rect 25964 34342 26016 34348
rect 26148 34400 26200 34406
rect 26148 34342 26200 34348
rect 26056 34196 26108 34202
rect 26056 34138 26108 34144
rect 25780 34060 25832 34066
rect 25780 34002 25832 34008
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25688 33516 25740 33522
rect 25688 33458 25740 33464
rect 25228 33448 25280 33454
rect 25228 33390 25280 33396
rect 25240 32910 25268 33390
rect 25412 33380 25464 33386
rect 25412 33322 25464 33328
rect 25228 32904 25280 32910
rect 25228 32846 25280 32852
rect 25424 31822 25452 33322
rect 25596 32972 25648 32978
rect 25596 32914 25648 32920
rect 25504 32496 25556 32502
rect 25504 32438 25556 32444
rect 25412 31816 25464 31822
rect 25412 31758 25464 31764
rect 25148 31726 25268 31754
rect 24676 31408 24728 31414
rect 24676 31350 24728 31356
rect 24688 30598 24716 31350
rect 24952 31136 25004 31142
rect 24952 31078 25004 31084
rect 24860 30660 24912 30666
rect 24860 30602 24912 30608
rect 24676 30592 24728 30598
rect 24676 30534 24728 30540
rect 24688 29714 24716 30534
rect 24768 30184 24820 30190
rect 24768 30126 24820 30132
rect 24780 29850 24808 30126
rect 24872 30054 24900 30602
rect 24860 30048 24912 30054
rect 24860 29990 24912 29996
rect 24768 29844 24820 29850
rect 24768 29786 24820 29792
rect 24676 29708 24728 29714
rect 24676 29650 24728 29656
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24780 28490 24808 29446
rect 24768 28484 24820 28490
rect 24768 28426 24820 28432
rect 24872 27470 24900 29990
rect 24964 29850 24992 31078
rect 25044 30184 25096 30190
rect 25044 30126 25096 30132
rect 24952 29844 25004 29850
rect 24952 29786 25004 29792
rect 24964 29186 24992 29786
rect 25056 29646 25084 30126
rect 25044 29640 25096 29646
rect 25044 29582 25096 29588
rect 24964 29158 25084 29186
rect 24952 29096 25004 29102
rect 24952 29038 25004 29044
rect 24860 27464 24912 27470
rect 24860 27406 24912 27412
rect 24964 27402 24992 29038
rect 25056 27441 25084 29158
rect 25042 27432 25098 27441
rect 24952 27396 25004 27402
rect 25042 27367 25098 27376
rect 25136 27396 25188 27402
rect 24952 27338 25004 27344
rect 25136 27338 25188 27344
rect 24492 27124 24544 27130
rect 24492 27066 24544 27072
rect 24308 26988 24360 26994
rect 24308 26930 24360 26936
rect 24216 26852 24268 26858
rect 24216 26794 24268 26800
rect 23848 26784 23900 26790
rect 23848 26726 23900 26732
rect 23664 26308 23716 26314
rect 23664 26250 23716 26256
rect 23032 25486 23152 25514
rect 22376 25356 22428 25362
rect 22376 25298 22428 25304
rect 22284 25220 22336 25226
rect 22284 25162 22336 25168
rect 22296 23866 22324 25162
rect 23032 24818 23060 25486
rect 23676 25430 23704 26250
rect 23860 26042 23888 26726
rect 24320 26314 24348 26930
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24676 26852 24728 26858
rect 24676 26794 24728 26800
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24596 26518 24624 26726
rect 24584 26512 24636 26518
rect 24584 26454 24636 26460
rect 24308 26308 24360 26314
rect 24308 26250 24360 26256
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 24596 25906 24624 26454
rect 24688 26382 24716 26794
rect 24872 26382 24900 26862
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24688 25906 24716 26318
rect 24216 25900 24268 25906
rect 24216 25842 24268 25848
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 23664 25424 23716 25430
rect 23664 25366 23716 25372
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23492 24818 23520 25230
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23032 24698 23060 24754
rect 23032 24670 23152 24698
rect 23020 24608 23072 24614
rect 23020 24550 23072 24556
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 23032 23798 23060 24550
rect 23124 24206 23152 24670
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 23020 23792 23072 23798
rect 23020 23734 23072 23740
rect 23124 23662 23152 24142
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23492 23798 23520 24006
rect 23480 23792 23532 23798
rect 23480 23734 23532 23740
rect 23112 23656 23164 23662
rect 23112 23598 23164 23604
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22296 23118 22324 23462
rect 23480 23180 23532 23186
rect 23480 23122 23532 23128
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 22020 21622 22048 22374
rect 22112 21894 22140 22918
rect 22204 22902 22324 22930
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22204 22030 22232 22578
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 21744 20330 21772 21490
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 21732 20324 21784 20330
rect 21732 20266 21784 20272
rect 21824 20324 21876 20330
rect 21824 20266 21876 20272
rect 21744 19990 21772 20266
rect 21732 19984 21784 19990
rect 21732 19926 21784 19932
rect 21744 19446 21772 19926
rect 21836 19718 21864 20266
rect 21916 19780 21968 19786
rect 21916 19722 21968 19728
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21836 19378 21864 19654
rect 21928 19446 21956 19722
rect 21916 19440 21968 19446
rect 21916 19382 21968 19388
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 22112 19310 22140 20470
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22204 17270 22232 18226
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22296 17218 22324 22902
rect 23492 22574 23520 23122
rect 23112 22568 23164 22574
rect 23112 22510 23164 22516
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23124 22234 23152 22510
rect 23848 22500 23900 22506
rect 23848 22442 23900 22448
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 22652 20868 22704 20874
rect 22652 20810 22704 20816
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 22664 20398 22692 20810
rect 23400 20602 23428 20810
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23492 20466 23520 22374
rect 23860 21146 23888 22442
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 23860 20534 23888 21082
rect 23848 20528 23900 20534
rect 23848 20470 23900 20476
rect 23480 20460 23532 20466
rect 23532 20420 23612 20448
rect 23480 20402 23532 20408
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22388 18698 22416 19110
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 22572 18630 22600 19246
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 22744 17808 22796 17814
rect 22744 17750 22796 17756
rect 22756 17270 22784 17750
rect 22744 17264 22796 17270
rect 22296 17190 22416 17218
rect 22744 17206 22796 17212
rect 21824 17060 21876 17066
rect 21824 17002 21876 17008
rect 21836 13938 21864 17002
rect 22100 16516 22152 16522
rect 22100 16458 22152 16464
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21928 15434 21956 16390
rect 22112 16114 22140 16458
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 22112 15366 22140 16050
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 22112 14958 22140 15302
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22296 14550 22324 14894
rect 22284 14544 22336 14550
rect 22284 14486 22336 14492
rect 22192 14340 22244 14346
rect 22192 14282 22244 14288
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 22020 14006 22048 14214
rect 22008 14000 22060 14006
rect 22008 13942 22060 13948
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 22204 13530 22232 14282
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 21284 6886 21496 6914
rect 21088 3120 21140 3126
rect 21088 3062 21140 3068
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2858
rect 21284 2582 21312 6886
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 21468 4146 21496 4422
rect 21928 4282 21956 4558
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21376 3738 21404 4082
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 22112 3466 22140 4558
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 22296 3058 22324 3470
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 21272 2576 21324 2582
rect 21272 2518 21324 2524
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 20640 800 20668 2314
rect 21928 800 21956 2314
rect 22388 2038 22416 17190
rect 22468 17196 22520 17202
rect 22468 17138 22520 17144
rect 22480 17066 22508 17138
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22480 16726 22508 17002
rect 23124 16794 23152 18566
rect 23308 18290 23336 19654
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 23296 17604 23348 17610
rect 23296 17546 23348 17552
rect 23308 17066 23336 17546
rect 23400 17270 23428 17682
rect 23492 17678 23520 18158
rect 23584 17882 23612 20420
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23768 18902 23796 19314
rect 23756 18896 23808 18902
rect 23756 18838 23808 18844
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 23492 17202 23520 17614
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 22468 16720 22520 16726
rect 22468 16662 22520 16668
rect 22572 16114 22600 16730
rect 23492 16114 23520 16934
rect 23676 16522 23704 17478
rect 23664 16516 23716 16522
rect 23664 16458 23716 16464
rect 23768 16114 23796 17818
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23860 16658 23888 17478
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23860 16182 23888 16594
rect 23848 16176 23900 16182
rect 23848 16118 23900 16124
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23756 16108 23808 16114
rect 23756 16050 23808 16056
rect 22572 15502 22600 16050
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 23124 15570 23152 15846
rect 23492 15706 23520 16050
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23860 15586 23888 16118
rect 23768 15570 23888 15586
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 23756 15564 23888 15570
rect 23808 15558 23888 15564
rect 23756 15506 23808 15512
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22480 13326 22508 14418
rect 22572 14278 22600 15438
rect 23940 14952 23992 14958
rect 23940 14894 23992 14900
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22480 4622 22508 4966
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22480 3126 22508 3878
rect 22468 3120 22520 3126
rect 22468 3062 22520 3068
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22376 2032 22428 2038
rect 22376 1974 22428 1980
rect 22572 800 22600 2926
rect 22848 2310 22876 13806
rect 23204 5160 23256 5166
rect 23204 5102 23256 5108
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 22940 2446 22968 4966
rect 23020 4548 23072 4554
rect 23020 4490 23072 4496
rect 23032 3534 23060 4490
rect 23216 4146 23244 5102
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23124 3738 23152 4082
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23492 2802 23520 4558
rect 23584 3942 23612 14418
rect 23952 6866 23980 14894
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23664 4752 23716 4758
rect 23664 4694 23716 4700
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23676 3534 23704 4694
rect 23860 4078 23888 5170
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23216 2774 23520 2802
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 23216 800 23244 2774
rect 24228 2650 24256 25842
rect 24872 25838 24900 26318
rect 25044 26240 25096 26246
rect 25044 26182 25096 26188
rect 24860 25832 24912 25838
rect 24860 25774 24912 25780
rect 24768 25696 24820 25702
rect 24768 25638 24820 25644
rect 24676 25424 24728 25430
rect 24676 25366 24728 25372
rect 24688 24818 24716 25366
rect 24780 25362 24808 25638
rect 24768 25356 24820 25362
rect 24768 25298 24820 25304
rect 24676 24812 24728 24818
rect 24676 24754 24728 24760
rect 24872 23662 24900 25774
rect 25056 25294 25084 26182
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24400 23588 24452 23594
rect 24400 23530 24452 23536
rect 24412 19242 24440 23530
rect 24492 20460 24544 20466
rect 24492 20402 24544 20408
rect 24504 19854 24532 20402
rect 24584 20324 24636 20330
rect 24584 20266 24636 20272
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24596 19378 24624 20266
rect 24766 19408 24822 19417
rect 24584 19372 24636 19378
rect 24766 19343 24822 19352
rect 24584 19314 24636 19320
rect 24400 19236 24452 19242
rect 24400 19178 24452 19184
rect 24412 18766 24440 19178
rect 24400 18760 24452 18766
rect 24400 18702 24452 18708
rect 24412 17678 24440 18702
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 24504 18086 24532 18362
rect 24492 18080 24544 18086
rect 24492 18022 24544 18028
rect 24596 17814 24624 19314
rect 24780 18766 24808 19343
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24872 18834 24900 19110
rect 24860 18828 24912 18834
rect 24860 18770 24912 18776
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24688 18222 24716 18253
rect 24676 18216 24728 18222
rect 24780 18170 24808 18702
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24728 18164 24808 18170
rect 24676 18158 24808 18164
rect 24688 18142 24808 18158
rect 24584 17808 24636 17814
rect 24584 17750 24636 17756
rect 24688 17746 24716 18142
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 24504 16250 24532 17070
rect 24688 16726 24716 17478
rect 24780 17270 24808 18022
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24872 16454 24900 18226
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24492 16244 24544 16250
rect 24492 16186 24544 16192
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24412 15502 24440 15846
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24964 5098 24992 24754
rect 25148 23866 25176 27338
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25148 23118 25176 23802
rect 25240 23594 25268 31726
rect 25424 30410 25452 31758
rect 25516 31754 25544 32438
rect 25608 32434 25636 32914
rect 25700 32842 25728 33458
rect 25792 32842 25820 34002
rect 25872 33992 25924 33998
rect 25872 33934 25924 33940
rect 25884 33130 25912 33934
rect 25884 33102 26004 33130
rect 25976 33046 26004 33102
rect 25964 33040 26016 33046
rect 25964 32982 26016 32988
rect 25688 32836 25740 32842
rect 25688 32778 25740 32784
rect 25780 32836 25832 32842
rect 25780 32778 25832 32784
rect 25976 32502 26004 32982
rect 25964 32496 26016 32502
rect 25964 32438 26016 32444
rect 25596 32428 25648 32434
rect 25596 32370 25648 32376
rect 25964 32292 26016 32298
rect 25964 32234 26016 32240
rect 25976 32026 26004 32234
rect 25964 32020 26016 32026
rect 25964 31962 26016 31968
rect 25872 31952 25924 31958
rect 25872 31894 25924 31900
rect 25688 31816 25740 31822
rect 25688 31758 25740 31764
rect 25780 31816 25832 31822
rect 25780 31758 25832 31764
rect 25516 31726 25636 31754
rect 25608 30546 25636 31726
rect 25700 30938 25728 31758
rect 25688 30932 25740 30938
rect 25688 30874 25740 30880
rect 25608 30518 25728 30546
rect 25424 30382 25544 30410
rect 25412 30252 25464 30258
rect 25412 30194 25464 30200
rect 25424 29306 25452 30194
rect 25412 29300 25464 29306
rect 25412 29242 25464 29248
rect 25320 28960 25372 28966
rect 25320 28902 25372 28908
rect 25332 28490 25360 28902
rect 25320 28484 25372 28490
rect 25320 28426 25372 28432
rect 25412 28484 25464 28490
rect 25412 28426 25464 28432
rect 25424 28218 25452 28426
rect 25412 28212 25464 28218
rect 25412 28154 25464 28160
rect 25516 26314 25544 30382
rect 25700 30326 25728 30518
rect 25688 30320 25740 30326
rect 25688 30262 25740 30268
rect 25596 29232 25648 29238
rect 25596 29174 25648 29180
rect 25608 28218 25636 29174
rect 25596 28212 25648 28218
rect 25596 28154 25648 28160
rect 25688 27872 25740 27878
rect 25688 27814 25740 27820
rect 25700 26994 25728 27814
rect 25688 26988 25740 26994
rect 25688 26930 25740 26936
rect 25504 26308 25556 26314
rect 25504 26250 25556 26256
rect 25516 26042 25544 26250
rect 25504 26036 25556 26042
rect 25504 25978 25556 25984
rect 25412 25152 25464 25158
rect 25412 25094 25464 25100
rect 25228 23588 25280 23594
rect 25228 23530 25280 23536
rect 25136 23112 25188 23118
rect 25136 23054 25188 23060
rect 25148 22030 25176 23054
rect 25424 22234 25452 25094
rect 25516 24274 25544 25978
rect 25700 25770 25728 26930
rect 25688 25764 25740 25770
rect 25688 25706 25740 25712
rect 25688 25492 25740 25498
rect 25688 25434 25740 25440
rect 25700 25294 25728 25434
rect 25792 25362 25820 31758
rect 25780 25356 25832 25362
rect 25780 25298 25832 25304
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25792 24886 25820 25298
rect 25884 25158 25912 31894
rect 26068 31822 26096 34138
rect 26160 33590 26188 34342
rect 26148 33584 26200 33590
rect 26148 33526 26200 33532
rect 26240 33108 26292 33114
rect 26160 33068 26240 33096
rect 26160 32026 26188 33068
rect 26240 33050 26292 33056
rect 26148 32020 26200 32026
rect 26148 31962 26200 31968
rect 26056 31816 26108 31822
rect 26056 31758 26108 31764
rect 26056 31680 26108 31686
rect 26056 31622 26108 31628
rect 26068 31142 26096 31622
rect 26056 31136 26108 31142
rect 26056 31078 26108 31084
rect 26068 30734 26096 31078
rect 26160 30802 26188 31962
rect 26436 31754 26464 41386
rect 27356 36922 27384 45766
rect 28080 44872 28132 44878
rect 28080 44814 28132 44820
rect 27528 37188 27580 37194
rect 27528 37130 27580 37136
rect 27344 36916 27396 36922
rect 27344 36858 27396 36864
rect 27540 36718 27568 37130
rect 27528 36712 27580 36718
rect 27528 36654 27580 36660
rect 27160 35624 27212 35630
rect 27160 35566 27212 35572
rect 27172 34474 27200 35566
rect 27252 35284 27304 35290
rect 27252 35226 27304 35232
rect 27264 34932 27292 35226
rect 27540 35170 27568 36654
rect 28092 35290 28120 44814
rect 28172 36168 28224 36174
rect 28172 36110 28224 36116
rect 28184 35494 28212 36110
rect 28540 36032 28592 36038
rect 28540 35974 28592 35980
rect 28552 35698 28580 35974
rect 28540 35692 28592 35698
rect 28540 35634 28592 35640
rect 28448 35624 28500 35630
rect 28448 35566 28500 35572
rect 28172 35488 28224 35494
rect 28172 35430 28224 35436
rect 28080 35284 28132 35290
rect 28080 35226 28132 35232
rect 27448 35142 27568 35170
rect 28184 35170 28212 35430
rect 28184 35142 28304 35170
rect 27344 34944 27396 34950
rect 27264 34904 27344 34932
rect 27160 34468 27212 34474
rect 27160 34410 27212 34416
rect 27264 34406 27292 34904
rect 27344 34886 27396 34892
rect 27252 34400 27304 34406
rect 27252 34342 27304 34348
rect 27160 32496 27212 32502
rect 27160 32438 27212 32444
rect 26792 32224 26844 32230
rect 26792 32166 26844 32172
rect 26804 31822 26832 32166
rect 27172 32026 27200 32438
rect 27160 32020 27212 32026
rect 27160 31962 27212 31968
rect 26792 31816 26844 31822
rect 26792 31758 26844 31764
rect 26436 31726 26556 31754
rect 26332 31340 26384 31346
rect 26332 31282 26384 31288
rect 26344 30938 26372 31282
rect 26332 30932 26384 30938
rect 26332 30874 26384 30880
rect 26148 30796 26200 30802
rect 26148 30738 26200 30744
rect 26056 30728 26108 30734
rect 26056 30670 26108 30676
rect 25964 30320 26016 30326
rect 25964 30262 26016 30268
rect 25976 29646 26004 30262
rect 26068 30258 26096 30670
rect 26056 30252 26108 30258
rect 26056 30194 26108 30200
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 25976 29016 26004 29582
rect 26068 29578 26096 30194
rect 26160 29646 26188 30738
rect 26240 30728 26292 30734
rect 26240 30670 26292 30676
rect 26148 29640 26200 29646
rect 26148 29582 26200 29588
rect 26056 29572 26108 29578
rect 26056 29514 26108 29520
rect 26056 29028 26108 29034
rect 25976 28988 26056 29016
rect 26056 28970 26108 28976
rect 26068 28626 26096 28970
rect 26056 28620 26108 28626
rect 26056 28562 26108 28568
rect 26160 27470 26188 29582
rect 26252 28762 26280 30670
rect 26240 28756 26292 28762
rect 26240 28698 26292 28704
rect 26252 28098 26280 28698
rect 26332 28552 26384 28558
rect 26332 28494 26384 28500
rect 26344 28218 26372 28494
rect 26332 28212 26384 28218
rect 26332 28154 26384 28160
rect 26252 28070 26372 28098
rect 26344 28014 26372 28070
rect 26424 28076 26476 28082
rect 26424 28018 26476 28024
rect 26332 28008 26384 28014
rect 26332 27950 26384 27956
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26240 27328 26292 27334
rect 26240 27270 26292 27276
rect 26148 27124 26200 27130
rect 26148 27066 26200 27072
rect 25872 25152 25924 25158
rect 25872 25094 25924 25100
rect 25884 24954 25912 25094
rect 25872 24948 25924 24954
rect 25872 24890 25924 24896
rect 25780 24880 25832 24886
rect 25780 24822 25832 24828
rect 25688 24812 25740 24818
rect 25688 24754 25740 24760
rect 25504 24268 25556 24274
rect 25504 24210 25556 24216
rect 25700 24138 25728 24754
rect 25884 24682 25912 24890
rect 26160 24886 26188 27066
rect 26252 26858 26280 27270
rect 26240 26852 26292 26858
rect 26240 26794 26292 26800
rect 26344 26314 26372 27950
rect 26436 27674 26464 28018
rect 26424 27668 26476 27674
rect 26424 27610 26476 27616
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26148 24880 26200 24886
rect 26148 24822 26200 24828
rect 26424 24812 26476 24818
rect 26424 24754 26476 24760
rect 25872 24676 25924 24682
rect 25872 24618 25924 24624
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25976 24206 26004 24550
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 25688 24132 25740 24138
rect 25688 24074 25740 24080
rect 25504 24064 25556 24070
rect 25504 24006 25556 24012
rect 25516 23186 25544 24006
rect 25504 23180 25556 23186
rect 25504 23122 25556 23128
rect 25412 22228 25464 22234
rect 25412 22170 25464 22176
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25148 21554 25176 21966
rect 25688 21956 25740 21962
rect 25688 21898 25740 21904
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25700 21078 25728 21898
rect 25688 21072 25740 21078
rect 25688 21014 25740 21020
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25240 19922 25268 20198
rect 25516 19922 25544 20198
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25412 19780 25464 19786
rect 25412 19722 25464 19728
rect 25044 19304 25096 19310
rect 25044 19246 25096 19252
rect 25056 19174 25084 19246
rect 25044 19168 25096 19174
rect 25044 19110 25096 19116
rect 25424 18766 25452 19722
rect 25792 19514 25820 20402
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26252 19786 26280 20198
rect 26240 19780 26292 19786
rect 26240 19722 26292 19728
rect 25780 19508 25832 19514
rect 25780 19450 25832 19456
rect 25594 19408 25650 19417
rect 25594 19343 25596 19352
rect 25648 19343 25650 19352
rect 25596 19314 25648 19320
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25148 17134 25176 17614
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 25504 17264 25556 17270
rect 25504 17206 25556 17212
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25240 15026 25268 16594
rect 25516 16590 25544 17206
rect 25608 16658 25636 17478
rect 25780 17060 25832 17066
rect 25780 17002 25832 17008
rect 25792 16794 25820 17002
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 25332 15162 25360 15370
rect 25320 15156 25372 15162
rect 25320 15098 25372 15104
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 26436 12646 26464 24754
rect 26528 23594 26556 31726
rect 26804 30938 26832 31758
rect 27160 31476 27212 31482
rect 27160 31418 27212 31424
rect 26792 30932 26844 30938
rect 26792 30874 26844 30880
rect 26608 30048 26660 30054
rect 26608 29990 26660 29996
rect 26620 29510 26648 29990
rect 26608 29504 26660 29510
rect 26608 29446 26660 29452
rect 26620 25702 26648 29446
rect 26976 28484 27028 28490
rect 26976 28426 27028 28432
rect 26988 27713 27016 28426
rect 27172 28218 27200 31418
rect 27160 28212 27212 28218
rect 27160 28154 27212 28160
rect 27172 28098 27200 28154
rect 27080 28070 27200 28098
rect 27080 27878 27108 28070
rect 27160 28008 27212 28014
rect 27160 27950 27212 27956
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 26974 27704 27030 27713
rect 26804 27662 26974 27690
rect 26700 27396 26752 27402
rect 26700 27338 26752 27344
rect 26712 26382 26740 27338
rect 26700 26376 26752 26382
rect 26700 26318 26752 26324
rect 26804 26194 26832 27662
rect 26974 27639 27030 27648
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 27080 26586 27108 27406
rect 27068 26580 27120 26586
rect 27068 26522 27120 26528
rect 27172 26518 27200 27950
rect 27264 27606 27292 34342
rect 27342 28656 27398 28665
rect 27342 28591 27398 28600
rect 27252 27600 27304 27606
rect 27252 27542 27304 27548
rect 27264 27130 27292 27542
rect 27356 27282 27384 28591
rect 27448 28218 27476 35142
rect 28276 35086 28304 35142
rect 28172 35080 28224 35086
rect 28172 35022 28224 35028
rect 28264 35080 28316 35086
rect 28264 35022 28316 35028
rect 27620 35012 27672 35018
rect 27620 34954 27672 34960
rect 27632 34542 27660 34954
rect 27620 34536 27672 34542
rect 27620 34478 27672 34484
rect 28080 34536 28132 34542
rect 28080 34478 28132 34484
rect 27712 33516 27764 33522
rect 27712 33458 27764 33464
rect 27724 33114 27752 33458
rect 27988 33448 28040 33454
rect 27988 33390 28040 33396
rect 27712 33108 27764 33114
rect 27712 33050 27764 33056
rect 28000 33046 28028 33390
rect 27988 33040 28040 33046
rect 27988 32982 28040 32988
rect 27988 32428 28040 32434
rect 27988 32370 28040 32376
rect 27896 32360 27948 32366
rect 27896 32302 27948 32308
rect 27908 31890 27936 32302
rect 27896 31884 27948 31890
rect 27896 31826 27948 31832
rect 27804 31816 27856 31822
rect 27804 31758 27856 31764
rect 27528 31748 27580 31754
rect 27528 31690 27580 31696
rect 27540 31482 27568 31690
rect 27528 31476 27580 31482
rect 27528 31418 27580 31424
rect 27816 31396 27844 31758
rect 28000 31754 28028 32370
rect 28092 32366 28120 34478
rect 28184 33998 28212 35022
rect 28172 33992 28224 33998
rect 28172 33934 28224 33940
rect 28080 32360 28132 32366
rect 28080 32302 28132 32308
rect 27908 31726 28028 31754
rect 27908 31498 27936 31726
rect 27908 31470 28120 31498
rect 27816 31368 28028 31396
rect 27712 30320 27764 30326
rect 27712 30262 27764 30268
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 27540 29034 27568 30194
rect 27620 30048 27672 30054
rect 27620 29990 27672 29996
rect 27528 29028 27580 29034
rect 27528 28970 27580 28976
rect 27540 28558 27568 28970
rect 27528 28552 27580 28558
rect 27528 28494 27580 28500
rect 27436 28212 27488 28218
rect 27436 28154 27488 28160
rect 27448 28082 27476 28154
rect 27632 28150 27660 29990
rect 27724 28694 27752 30262
rect 27804 29572 27856 29578
rect 27804 29514 27856 29520
rect 27816 28762 27844 29514
rect 27896 29164 27948 29170
rect 27896 29106 27948 29112
rect 27804 28756 27856 28762
rect 27804 28698 27856 28704
rect 27712 28688 27764 28694
rect 27710 28656 27712 28665
rect 27764 28656 27766 28665
rect 27710 28591 27766 28600
rect 27804 28552 27856 28558
rect 27724 28512 27804 28540
rect 27620 28144 27672 28150
rect 27620 28086 27672 28092
rect 27436 28076 27488 28082
rect 27436 28018 27488 28024
rect 27620 27532 27672 27538
rect 27620 27474 27672 27480
rect 27356 27254 27476 27282
rect 27252 27124 27304 27130
rect 27252 27066 27304 27072
rect 27252 26920 27304 26926
rect 27252 26862 27304 26868
rect 27264 26586 27292 26862
rect 27344 26784 27396 26790
rect 27344 26726 27396 26732
rect 27252 26580 27304 26586
rect 27252 26522 27304 26528
rect 27160 26512 27212 26518
rect 27160 26454 27212 26460
rect 27172 26382 27200 26454
rect 27160 26376 27212 26382
rect 27160 26318 27212 26324
rect 26712 26166 26832 26194
rect 26608 25696 26660 25702
rect 26608 25638 26660 25644
rect 26516 23588 26568 23594
rect 26516 23530 26568 23536
rect 26712 20942 26740 26166
rect 27264 25906 27292 26522
rect 27356 26518 27384 26726
rect 27344 26512 27396 26518
rect 27344 26454 27396 26460
rect 27252 25900 27304 25906
rect 27252 25842 27304 25848
rect 27160 25696 27212 25702
rect 27160 25638 27212 25644
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 26988 24138 27016 24346
rect 26976 24132 27028 24138
rect 26976 24074 27028 24080
rect 26988 23322 27016 24074
rect 27172 23526 27200 25638
rect 27448 25498 27476 27254
rect 27632 27062 27660 27474
rect 27620 27056 27672 27062
rect 27620 26998 27672 27004
rect 27436 25492 27488 25498
rect 27436 25434 27488 25440
rect 27160 23520 27212 23526
rect 27160 23462 27212 23468
rect 26976 23316 27028 23322
rect 26976 23258 27028 23264
rect 27172 23118 27200 23462
rect 27160 23112 27212 23118
rect 27160 23054 27212 23060
rect 27068 23044 27120 23050
rect 27068 22986 27120 22992
rect 27080 22778 27108 22986
rect 27068 22772 27120 22778
rect 27068 22714 27120 22720
rect 26884 22704 26936 22710
rect 26884 22646 26936 22652
rect 26896 22234 26924 22646
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 26884 22228 26936 22234
rect 26884 22170 26936 22176
rect 26792 22092 26844 22098
rect 26792 22034 26844 22040
rect 26804 21894 26832 22034
rect 27356 22030 27384 22578
rect 27344 22024 27396 22030
rect 27344 21966 27396 21972
rect 26792 21888 26844 21894
rect 26792 21830 26844 21836
rect 27356 21146 27384 21966
rect 27344 21140 27396 21146
rect 27344 21082 27396 21088
rect 27356 20942 27384 21082
rect 26700 20936 26752 20942
rect 26700 20878 26752 20884
rect 27344 20936 27396 20942
rect 27344 20878 27396 20884
rect 26712 17678 26740 20878
rect 27356 20466 27384 20878
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27160 20324 27212 20330
rect 27160 20266 27212 20272
rect 27068 20256 27120 20262
rect 27068 20198 27120 20204
rect 27080 18698 27108 20198
rect 27172 19854 27200 20266
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27172 18902 27200 19790
rect 27632 19258 27660 20402
rect 27540 19230 27660 19258
rect 27160 18896 27212 18902
rect 27160 18838 27212 18844
rect 27068 18692 27120 18698
rect 27068 18634 27120 18640
rect 27540 18290 27568 19230
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 26700 17672 26752 17678
rect 26700 17614 26752 17620
rect 26884 17196 26936 17202
rect 26884 17138 26936 17144
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 26896 16658 26924 17138
rect 27172 16658 27200 17138
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 24952 5092 25004 5098
rect 24952 5034 25004 5040
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 24308 4480 24360 4486
rect 24308 4422 24360 4428
rect 24320 3126 24348 4422
rect 24412 3534 24440 4626
rect 25504 4616 25556 4622
rect 25504 4558 25556 4564
rect 24492 4140 24544 4146
rect 24492 4082 24544 4088
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24504 3738 24532 4082
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 24596 3398 24624 3674
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24308 3120 24360 3126
rect 24308 3062 24360 3068
rect 24872 2922 24900 4082
rect 24952 4072 25004 4078
rect 24952 4014 25004 4020
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24872 2446 24900 2858
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24492 2372 24544 2378
rect 24492 2314 24544 2320
rect 24504 800 24532 2314
rect 24964 2310 24992 4014
rect 25516 3534 25544 4558
rect 26896 4078 26924 16594
rect 27172 6914 27200 16594
rect 27540 14618 27568 18226
rect 27528 14612 27580 14618
rect 27528 14554 27580 14560
rect 26988 6886 27200 6914
rect 26240 4072 26292 4078
rect 26240 4014 26292 4020
rect 26884 4072 26936 4078
rect 26884 4014 26936 4020
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 25780 3460 25832 3466
rect 25780 3402 25832 3408
rect 25792 2922 25820 3402
rect 26252 3126 26280 4014
rect 26700 3664 26752 3670
rect 26700 3606 26752 3612
rect 26712 3126 26740 3606
rect 26056 3120 26108 3126
rect 26056 3062 26108 3068
rect 26240 3120 26292 3126
rect 26240 3062 26292 3068
rect 26700 3120 26752 3126
rect 26700 3062 26752 3068
rect 25136 2916 25188 2922
rect 25136 2858 25188 2864
rect 25780 2916 25832 2922
rect 25780 2858 25832 2864
rect 24952 2304 25004 2310
rect 24952 2246 25004 2252
rect 25148 800 25176 2858
rect 26068 2854 26096 3062
rect 26056 2848 26108 2854
rect 26056 2790 26108 2796
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 26252 2310 26280 2586
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26240 2304 26292 2310
rect 26240 2246 26292 2252
rect 26436 800 26464 2382
rect 26988 1970 27016 6886
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 27172 2582 27200 2994
rect 27160 2576 27212 2582
rect 27160 2518 27212 2524
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 26976 1964 27028 1970
rect 26976 1906 27028 1912
rect 27080 800 27108 2314
rect 27448 2106 27476 2450
rect 27724 2446 27752 28512
rect 27804 28494 27856 28500
rect 27804 28144 27856 28150
rect 27804 28086 27856 28092
rect 27816 26790 27844 28086
rect 27804 26784 27856 26790
rect 27804 26726 27856 26732
rect 27908 24682 27936 29106
rect 28000 28626 28028 31368
rect 27988 28620 28040 28626
rect 27988 28562 28040 28568
rect 28000 27402 28028 28562
rect 28092 28082 28120 31470
rect 28184 30326 28212 33934
rect 28460 33658 28488 35566
rect 28540 35488 28592 35494
rect 28540 35430 28592 35436
rect 28448 33652 28500 33658
rect 28448 33594 28500 33600
rect 28264 33516 28316 33522
rect 28264 33458 28316 33464
rect 28276 33046 28304 33458
rect 28356 33448 28408 33454
rect 28356 33390 28408 33396
rect 28264 33040 28316 33046
rect 28264 32982 28316 32988
rect 28276 32026 28304 32982
rect 28264 32020 28316 32026
rect 28264 31962 28316 31968
rect 28264 31884 28316 31890
rect 28264 31826 28316 31832
rect 28172 30320 28224 30326
rect 28172 30262 28224 30268
rect 28172 30184 28224 30190
rect 28172 30126 28224 30132
rect 28184 28694 28212 30126
rect 28172 28688 28224 28694
rect 28172 28630 28224 28636
rect 28172 28552 28224 28558
rect 28172 28494 28224 28500
rect 28080 28076 28132 28082
rect 28080 28018 28132 28024
rect 28184 27878 28212 28494
rect 28172 27872 28224 27878
rect 28172 27814 28224 27820
rect 28276 27470 28304 31826
rect 28264 27464 28316 27470
rect 28264 27406 28316 27412
rect 27988 27396 28040 27402
rect 27988 27338 28040 27344
rect 28172 27396 28224 27402
rect 28172 27338 28224 27344
rect 28000 27062 28028 27338
rect 27988 27056 28040 27062
rect 27988 26998 28040 27004
rect 27988 26920 28040 26926
rect 28184 26897 28212 27338
rect 27988 26862 28040 26868
rect 28170 26888 28226 26897
rect 28000 26790 28028 26862
rect 28170 26823 28226 26832
rect 27988 26784 28040 26790
rect 27988 26726 28040 26732
rect 27988 26580 28040 26586
rect 27988 26522 28040 26528
rect 28000 24818 28028 26522
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 27896 24676 27948 24682
rect 27896 24618 27948 24624
rect 28080 24608 28132 24614
rect 28080 24550 28132 24556
rect 28092 24274 28120 24550
rect 28080 24268 28132 24274
rect 28080 24210 28132 24216
rect 28092 23662 28120 24210
rect 28184 24206 28212 25298
rect 28264 24744 28316 24750
rect 28264 24686 28316 24692
rect 28276 24410 28304 24686
rect 28264 24404 28316 24410
rect 28264 24346 28316 24352
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28184 23866 28212 24142
rect 28172 23860 28224 23866
rect 28172 23802 28224 23808
rect 28080 23656 28132 23662
rect 28080 23598 28132 23604
rect 28092 22982 28120 23598
rect 28080 22976 28132 22982
rect 28080 22918 28132 22924
rect 28184 22642 28212 23802
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28276 22778 28304 23054
rect 28264 22772 28316 22778
rect 28264 22714 28316 22720
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 28080 22094 28132 22098
rect 28184 22094 28212 22578
rect 28080 22092 28212 22094
rect 28132 22066 28212 22092
rect 28080 22034 28132 22040
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 28000 21622 28028 21830
rect 27988 21616 28040 21622
rect 27988 21558 28040 21564
rect 28172 21616 28224 21622
rect 28172 21558 28224 21564
rect 28184 21146 28212 21558
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28264 19508 28316 19514
rect 28264 19450 28316 19456
rect 28276 19378 28304 19450
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 27804 18828 27856 18834
rect 27804 18770 27856 18776
rect 27816 17678 27844 18770
rect 28172 18624 28224 18630
rect 28172 18566 28224 18572
rect 28184 18290 28212 18566
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27816 17270 27844 17614
rect 27804 17264 27856 17270
rect 27804 17206 27856 17212
rect 28368 2650 28396 33390
rect 28448 33380 28500 33386
rect 28448 33322 28500 33328
rect 28460 32178 28488 33322
rect 28552 32910 28580 35430
rect 28632 34128 28684 34134
rect 28632 34070 28684 34076
rect 28540 32904 28592 32910
rect 28540 32846 28592 32852
rect 28644 32434 28672 34070
rect 28816 33992 28868 33998
rect 28816 33934 28868 33940
rect 28724 33584 28776 33590
rect 28724 33526 28776 33532
rect 28736 32910 28764 33526
rect 28828 33114 28856 33934
rect 28816 33108 28868 33114
rect 28816 33050 28868 33056
rect 28724 32904 28776 32910
rect 28724 32846 28776 32852
rect 28632 32428 28684 32434
rect 28632 32370 28684 32376
rect 28828 32366 28856 33050
rect 28816 32360 28868 32366
rect 28920 32337 28948 47058
rect 29012 34746 29040 47126
rect 29656 47054 29684 49200
rect 29828 47184 29880 47190
rect 29828 47126 29880 47132
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 29840 41414 29868 47126
rect 30944 47054 30972 49200
rect 30932 47048 30984 47054
rect 30932 46990 30984 46996
rect 31392 46980 31444 46986
rect 31392 46922 31444 46928
rect 31404 41414 31432 46922
rect 32232 46442 32260 49200
rect 38028 47682 38056 49200
rect 37292 47654 38056 47682
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 33692 47184 33744 47190
rect 33692 47126 33744 47132
rect 32404 46504 32456 46510
rect 32404 46446 32456 46452
rect 33324 46504 33376 46510
rect 33324 46446 33376 46452
rect 32220 46436 32272 46442
rect 32220 46378 32272 46384
rect 32416 46170 32444 46446
rect 32404 46164 32456 46170
rect 32404 46106 32456 46112
rect 33336 45558 33364 46446
rect 33324 45552 33376 45558
rect 33324 45494 33376 45500
rect 29840 41386 30328 41414
rect 29920 35828 29972 35834
rect 29920 35770 29972 35776
rect 29276 35760 29328 35766
rect 29276 35702 29328 35708
rect 29288 34746 29316 35702
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 29276 34740 29328 34746
rect 29276 34682 29328 34688
rect 29460 34740 29512 34746
rect 29460 34682 29512 34688
rect 29092 34060 29144 34066
rect 29092 34002 29144 34008
rect 29104 33522 29132 34002
rect 29472 33658 29500 34682
rect 29932 34610 29960 35770
rect 29552 34604 29604 34610
rect 29552 34546 29604 34552
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29564 34202 29592 34546
rect 29552 34196 29604 34202
rect 29552 34138 29604 34144
rect 29460 33652 29512 33658
rect 29460 33594 29512 33600
rect 30104 33584 30156 33590
rect 30104 33526 30156 33532
rect 29092 33516 29144 33522
rect 29092 33458 29144 33464
rect 29104 32910 29132 33458
rect 29552 32972 29604 32978
rect 29552 32914 29604 32920
rect 29092 32904 29144 32910
rect 29092 32846 29144 32852
rect 29104 32434 29132 32846
rect 29564 32774 29592 32914
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 29552 32768 29604 32774
rect 29552 32710 29604 32716
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 28816 32302 28868 32308
rect 28906 32328 28962 32337
rect 28906 32263 28962 32272
rect 28460 32150 28994 32178
rect 28448 31884 28500 31890
rect 28448 31826 28500 31832
rect 28460 27674 28488 31826
rect 28540 30796 28592 30802
rect 28540 30738 28592 30744
rect 28552 30122 28580 30738
rect 28724 30728 28776 30734
rect 28724 30670 28776 30676
rect 28632 30660 28684 30666
rect 28632 30602 28684 30608
rect 28540 30116 28592 30122
rect 28540 30058 28592 30064
rect 28552 28558 28580 30058
rect 28644 28626 28672 30602
rect 28736 29594 28764 30670
rect 28828 29714 28856 32150
rect 28966 32042 28994 32150
rect 28966 32014 29040 32042
rect 29104 32026 29132 32370
rect 28906 31920 28962 31929
rect 29012 31906 29040 32014
rect 29092 32020 29144 32026
rect 29092 31962 29144 31968
rect 29276 31952 29328 31958
rect 29012 31900 29276 31906
rect 29012 31894 29328 31900
rect 29012 31878 29316 31894
rect 28906 31855 28962 31864
rect 28816 29708 28868 29714
rect 28816 29650 28868 29656
rect 28736 29566 28856 29594
rect 28828 28762 28856 29566
rect 28816 28756 28868 28762
rect 28816 28698 28868 28704
rect 28632 28620 28684 28626
rect 28632 28562 28684 28568
rect 28540 28552 28592 28558
rect 28540 28494 28592 28500
rect 28538 27704 28594 27713
rect 28448 27668 28500 27674
rect 28538 27639 28540 27648
rect 28448 27610 28500 27616
rect 28592 27639 28594 27648
rect 28540 27610 28592 27616
rect 28460 27334 28488 27610
rect 28540 27464 28592 27470
rect 28540 27406 28592 27412
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 28552 27130 28580 27406
rect 28540 27124 28592 27130
rect 28540 27066 28592 27072
rect 28644 27010 28672 28562
rect 28724 28552 28776 28558
rect 28724 28494 28776 28500
rect 28736 28218 28764 28494
rect 28724 28212 28776 28218
rect 28724 28154 28776 28160
rect 28722 27432 28778 27441
rect 28722 27367 28724 27376
rect 28776 27367 28778 27376
rect 28724 27338 28776 27344
rect 28736 27130 28764 27338
rect 28724 27124 28776 27130
rect 28724 27066 28776 27072
rect 28552 26982 28672 27010
rect 28552 26450 28580 26982
rect 28632 26920 28684 26926
rect 28632 26862 28684 26868
rect 28540 26444 28592 26450
rect 28460 26404 28540 26432
rect 28460 24410 28488 26404
rect 28540 26386 28592 26392
rect 28644 25906 28672 26862
rect 28736 26382 28764 27066
rect 28724 26376 28776 26382
rect 28724 26318 28776 26324
rect 28632 25900 28684 25906
rect 28632 25842 28684 25848
rect 28644 25378 28672 25842
rect 28552 25350 28672 25378
rect 28552 25294 28580 25350
rect 28540 25288 28592 25294
rect 28540 25230 28592 25236
rect 28828 25226 28856 28698
rect 28816 25220 28868 25226
rect 28816 25162 28868 25168
rect 28920 25106 28948 31855
rect 29000 30932 29052 30938
rect 29000 30874 29052 30880
rect 29012 30258 29040 30874
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 29012 29850 29040 30194
rect 29000 29844 29052 29850
rect 29000 29786 29052 29792
rect 29564 29782 29592 32710
rect 29932 32502 29960 32846
rect 29644 32496 29696 32502
rect 29644 32438 29696 32444
rect 29920 32496 29972 32502
rect 29920 32438 29972 32444
rect 29656 30938 29684 32438
rect 30116 32434 30144 33526
rect 30104 32428 30156 32434
rect 30104 32370 30156 32376
rect 30300 31754 30328 41386
rect 31220 41386 31432 41414
rect 30656 35760 30708 35766
rect 30656 35702 30708 35708
rect 30380 35488 30432 35494
rect 30380 35430 30432 35436
rect 30392 34066 30420 35430
rect 30668 35290 30696 35702
rect 30840 35488 30892 35494
rect 30840 35430 30892 35436
rect 30656 35284 30708 35290
rect 30656 35226 30708 35232
rect 30380 34060 30432 34066
rect 30380 34002 30432 34008
rect 30380 33924 30432 33930
rect 30380 33866 30432 33872
rect 30748 33924 30800 33930
rect 30748 33866 30800 33872
rect 30392 33522 30420 33866
rect 30380 33516 30432 33522
rect 30380 33458 30432 33464
rect 30392 33046 30420 33458
rect 30760 33114 30788 33866
rect 30852 33862 30880 35430
rect 31116 35148 31168 35154
rect 31116 35090 31168 35096
rect 31128 34746 31156 35090
rect 31116 34740 31168 34746
rect 31116 34682 31168 34688
rect 30932 34196 30984 34202
rect 30932 34138 30984 34144
rect 30944 33862 30972 34138
rect 30840 33856 30892 33862
rect 30840 33798 30892 33804
rect 30932 33856 30984 33862
rect 30932 33798 30984 33804
rect 30852 33522 30880 33798
rect 30840 33516 30892 33522
rect 30840 33458 30892 33464
rect 30932 33516 30984 33522
rect 30932 33458 30984 33464
rect 30852 33318 30880 33458
rect 30840 33312 30892 33318
rect 30840 33254 30892 33260
rect 30656 33108 30708 33114
rect 30656 33050 30708 33056
rect 30748 33108 30800 33114
rect 30748 33050 30800 33056
rect 30380 33040 30432 33046
rect 30380 32982 30432 32988
rect 30668 32994 30696 33050
rect 30668 32966 30880 32994
rect 30944 32978 30972 33458
rect 30852 32910 30880 32966
rect 30932 32972 30984 32978
rect 30932 32914 30984 32920
rect 30656 32904 30708 32910
rect 30656 32846 30708 32852
rect 30840 32904 30892 32910
rect 30840 32846 30892 32852
rect 30564 32768 30616 32774
rect 30564 32710 30616 32716
rect 30472 32428 30524 32434
rect 30472 32370 30524 32376
rect 30484 31890 30512 32370
rect 30576 32366 30604 32710
rect 30564 32360 30616 32366
rect 30564 32302 30616 32308
rect 30472 31884 30524 31890
rect 30472 31826 30524 31832
rect 30116 31726 30328 31754
rect 30668 31754 30696 32846
rect 30748 32768 30800 32774
rect 30748 32710 30800 32716
rect 30760 32230 30788 32710
rect 30944 32502 30972 32914
rect 30932 32496 30984 32502
rect 30932 32438 30984 32444
rect 31220 32314 31248 41386
rect 33416 36168 33468 36174
rect 33416 36110 33468 36116
rect 33324 36032 33376 36038
rect 33324 35974 33376 35980
rect 31760 34944 31812 34950
rect 31760 34886 31812 34892
rect 31300 34672 31352 34678
rect 31300 34614 31352 34620
rect 31312 33266 31340 34614
rect 31668 34536 31720 34542
rect 31668 34478 31720 34484
rect 31680 34082 31708 34478
rect 31496 34066 31708 34082
rect 31484 34060 31708 34066
rect 31536 34054 31708 34060
rect 31484 34002 31536 34008
rect 31312 33238 31524 33266
rect 31128 32286 31248 32314
rect 30748 32224 30800 32230
rect 30748 32166 30800 32172
rect 31128 31754 31156 32286
rect 31208 32224 31260 32230
rect 31208 32166 31260 32172
rect 31300 32224 31352 32230
rect 31300 32166 31352 32172
rect 31220 31958 31248 32166
rect 31312 31958 31340 32166
rect 31208 31952 31260 31958
rect 31208 31894 31260 31900
rect 31300 31952 31352 31958
rect 31300 31894 31352 31900
rect 30668 31726 30880 31754
rect 29644 30932 29696 30938
rect 29644 30874 29696 30880
rect 29552 29776 29604 29782
rect 29552 29718 29604 29724
rect 29276 29572 29328 29578
rect 29276 29514 29328 29520
rect 29092 28076 29144 28082
rect 29092 28018 29144 28024
rect 29104 27606 29132 28018
rect 29092 27600 29144 27606
rect 29092 27542 29144 27548
rect 29288 27130 29316 29514
rect 29276 27124 29328 27130
rect 29276 27066 29328 27072
rect 29184 26988 29236 26994
rect 29184 26930 29236 26936
rect 29196 26314 29224 26930
rect 29184 26308 29236 26314
rect 29184 26250 29236 26256
rect 29276 25288 29328 25294
rect 29276 25230 29328 25236
rect 29366 25256 29422 25265
rect 28736 25078 28948 25106
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28448 24404 28500 24410
rect 28448 24346 28500 24352
rect 28552 24206 28580 24754
rect 28632 24404 28684 24410
rect 28632 24346 28684 24352
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28448 24064 28500 24070
rect 28448 24006 28500 24012
rect 28460 23730 28488 24006
rect 28644 23730 28672 24346
rect 28448 23724 28500 23730
rect 28448 23666 28500 23672
rect 28632 23724 28684 23730
rect 28632 23666 28684 23672
rect 28460 22642 28488 23666
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28736 19514 28764 25078
rect 29288 24818 29316 25230
rect 29366 25191 29368 25200
rect 29420 25191 29422 25200
rect 29368 25162 29420 25168
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 29564 24342 29592 29718
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29736 29572 29788 29578
rect 29736 29514 29788 29520
rect 29644 26444 29696 26450
rect 29644 26386 29696 26392
rect 29656 26042 29684 26386
rect 29644 26036 29696 26042
rect 29644 25978 29696 25984
rect 29642 25528 29698 25537
rect 29642 25463 29698 25472
rect 29656 25294 29684 25463
rect 29644 25288 29696 25294
rect 29644 25230 29696 25236
rect 29644 25152 29696 25158
rect 29644 25094 29696 25100
rect 29656 24886 29684 25094
rect 29644 24880 29696 24886
rect 29644 24822 29696 24828
rect 29552 24336 29604 24342
rect 29552 24278 29604 24284
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 29564 23866 29592 24142
rect 29552 23860 29604 23866
rect 29552 23802 29604 23808
rect 29642 23760 29698 23769
rect 29642 23695 29644 23704
rect 29696 23695 29698 23704
rect 29644 23666 29696 23672
rect 28816 23248 28868 23254
rect 28816 23190 28868 23196
rect 28828 22030 28856 23190
rect 28908 22636 28960 22642
rect 28908 22578 28960 22584
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 28920 21486 28948 22578
rect 29460 22432 29512 22438
rect 29460 22374 29512 22380
rect 29472 21962 29500 22374
rect 29460 21956 29512 21962
rect 29460 21898 29512 21904
rect 29276 21888 29328 21894
rect 29276 21830 29328 21836
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 28998 21040 29054 21049
rect 28998 20975 29054 20984
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28736 18766 28764 19450
rect 28908 19372 28960 19378
rect 29012 19360 29040 20975
rect 28960 19332 29040 19360
rect 28908 19314 28960 19320
rect 29012 18766 29040 19332
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 29104 18902 29132 19246
rect 29092 18896 29144 18902
rect 29092 18838 29144 18844
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 28736 17746 28764 18702
rect 28724 17740 28776 17746
rect 28724 17682 28776 17688
rect 28632 17672 28684 17678
rect 28632 17614 28684 17620
rect 28644 16794 28672 17614
rect 29012 17610 29040 18702
rect 29000 17604 29052 17610
rect 29000 17546 29052 17552
rect 28632 16788 28684 16794
rect 28632 16730 28684 16736
rect 29288 16658 29316 21830
rect 29748 18426 29776 29514
rect 29840 28762 29868 29582
rect 29828 28756 29880 28762
rect 29828 28698 29880 28704
rect 29828 27464 29880 27470
rect 29828 27406 29880 27412
rect 29840 22574 29868 27406
rect 29920 26784 29972 26790
rect 29920 26726 29972 26732
rect 29932 26382 29960 26726
rect 29920 26376 29972 26382
rect 29920 26318 29972 26324
rect 29920 25288 29972 25294
rect 29920 25230 29972 25236
rect 29932 24954 29960 25230
rect 29920 24948 29972 24954
rect 29920 24890 29972 24896
rect 30012 24948 30064 24954
rect 30012 24890 30064 24896
rect 29920 24812 29972 24818
rect 29920 24754 29972 24760
rect 29932 24206 29960 24754
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 30024 22930 30052 24890
rect 30116 24290 30144 31726
rect 30472 30728 30524 30734
rect 30472 30670 30524 30676
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 30392 29102 30420 29582
rect 30380 29096 30432 29102
rect 30380 29038 30432 29044
rect 30392 28422 30420 29038
rect 30484 28762 30512 30670
rect 30656 30592 30708 30598
rect 30656 30534 30708 30540
rect 30564 30184 30616 30190
rect 30564 30126 30616 30132
rect 30576 29850 30604 30126
rect 30564 29844 30616 29850
rect 30564 29786 30616 29792
rect 30668 29714 30696 30534
rect 30748 29844 30800 29850
rect 30748 29786 30800 29792
rect 30656 29708 30708 29714
rect 30656 29650 30708 29656
rect 30656 29572 30708 29578
rect 30656 29514 30708 29520
rect 30668 29170 30696 29514
rect 30656 29164 30708 29170
rect 30656 29106 30708 29112
rect 30564 29028 30616 29034
rect 30564 28970 30616 28976
rect 30472 28756 30524 28762
rect 30472 28698 30524 28704
rect 30576 28558 30604 28970
rect 30668 28694 30696 29106
rect 30760 29034 30788 29786
rect 30748 29028 30800 29034
rect 30748 28970 30800 28976
rect 30656 28688 30708 28694
rect 30656 28630 30708 28636
rect 30564 28552 30616 28558
rect 30564 28494 30616 28500
rect 30380 28416 30432 28422
rect 30380 28358 30432 28364
rect 30748 27872 30800 27878
rect 30748 27814 30800 27820
rect 30760 27606 30788 27814
rect 30748 27600 30800 27606
rect 30748 27542 30800 27548
rect 30760 27402 30788 27542
rect 30748 27396 30800 27402
rect 30748 27338 30800 27344
rect 30656 27328 30708 27334
rect 30656 27270 30708 27276
rect 30380 26512 30432 26518
rect 30380 26454 30432 26460
rect 30196 26376 30248 26382
rect 30196 26318 30248 26324
rect 30208 26246 30236 26318
rect 30196 26240 30248 26246
rect 30196 26182 30248 26188
rect 30288 25288 30340 25294
rect 30208 25248 30288 25276
rect 30208 24410 30236 25248
rect 30288 25230 30340 25236
rect 30288 24948 30340 24954
rect 30392 24936 30420 26454
rect 30668 25226 30696 27270
rect 30656 25220 30708 25226
rect 30656 25162 30708 25168
rect 30340 24908 30420 24936
rect 30288 24890 30340 24896
rect 30564 24880 30616 24886
rect 30564 24822 30616 24828
rect 30576 24750 30604 24822
rect 30564 24744 30616 24750
rect 30564 24686 30616 24692
rect 30380 24608 30432 24614
rect 30380 24550 30432 24556
rect 30472 24608 30524 24614
rect 30472 24550 30524 24556
rect 30196 24404 30248 24410
rect 30196 24346 30248 24352
rect 30392 24342 30420 24550
rect 30484 24410 30512 24550
rect 30576 24410 30604 24686
rect 30472 24404 30524 24410
rect 30472 24346 30524 24352
rect 30564 24404 30616 24410
rect 30564 24346 30616 24352
rect 30380 24336 30432 24342
rect 30116 24262 30328 24290
rect 30380 24278 30432 24284
rect 30196 24200 30248 24206
rect 30196 24142 30248 24148
rect 30102 23760 30158 23769
rect 30102 23695 30104 23704
rect 30156 23695 30158 23704
rect 30104 23666 30156 23672
rect 30208 23186 30236 24142
rect 30196 23180 30248 23186
rect 30196 23122 30248 23128
rect 30024 22902 30144 22930
rect 29828 22568 29880 22574
rect 29828 22510 29880 22516
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 29460 17128 29512 17134
rect 29460 17070 29512 17076
rect 29472 16794 29500 17070
rect 29460 16788 29512 16794
rect 29460 16730 29512 16736
rect 29276 16652 29328 16658
rect 29276 16594 29328 16600
rect 29552 16584 29604 16590
rect 29552 16526 29604 16532
rect 29564 10674 29592 16526
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 29564 4010 29592 10610
rect 29840 8838 29868 22510
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 30012 20392 30064 20398
rect 30012 20334 30064 20340
rect 29932 19514 29960 20334
rect 30024 20058 30052 20334
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29932 18834 29960 19450
rect 29920 18828 29972 18834
rect 29920 18770 29972 18776
rect 30012 18692 30064 18698
rect 30012 18634 30064 18640
rect 29828 8832 29880 8838
rect 29828 8774 29880 8780
rect 30024 4078 30052 18634
rect 30012 4072 30064 4078
rect 30012 4014 30064 4020
rect 29552 4004 29604 4010
rect 29552 3946 29604 3952
rect 28356 2644 28408 2650
rect 28356 2586 28408 2592
rect 29736 2644 29788 2650
rect 29736 2586 29788 2592
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 27436 2100 27488 2106
rect 27436 2042 27488 2048
rect 28368 800 28396 2314
rect 29656 800 29684 2382
rect 29748 2378 29776 2586
rect 30116 2582 30144 22902
rect 30208 22642 30236 23122
rect 30196 22636 30248 22642
rect 30196 22578 30248 22584
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30208 20806 30236 20946
rect 30300 20874 30328 24262
rect 30576 24070 30604 24346
rect 30564 24064 30616 24070
rect 30564 24006 30616 24012
rect 30668 23882 30696 25162
rect 30576 23854 30696 23882
rect 30472 23724 30524 23730
rect 30392 23684 30472 23712
rect 30392 23322 30420 23684
rect 30472 23666 30524 23672
rect 30380 23316 30432 23322
rect 30380 23258 30432 23264
rect 30392 23118 30420 23258
rect 30380 23112 30432 23118
rect 30380 23054 30432 23060
rect 30576 23050 30604 23854
rect 30564 23044 30616 23050
rect 30564 22986 30616 22992
rect 30576 22778 30604 22986
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30852 22094 30880 31726
rect 30944 31726 31156 31754
rect 30944 23118 30972 31726
rect 31208 31476 31260 31482
rect 31208 31418 31260 31424
rect 31024 30728 31076 30734
rect 31024 30670 31076 30676
rect 31036 29034 31064 30670
rect 31116 30660 31168 30666
rect 31116 30602 31168 30608
rect 31128 30122 31156 30602
rect 31116 30116 31168 30122
rect 31116 30058 31168 30064
rect 31220 30002 31248 31418
rect 31392 30796 31444 30802
rect 31392 30738 31444 30744
rect 31300 30728 31352 30734
rect 31300 30670 31352 30676
rect 31312 30190 31340 30670
rect 31300 30184 31352 30190
rect 31300 30126 31352 30132
rect 31404 30054 31432 30738
rect 31392 30048 31444 30054
rect 31220 29974 31340 30002
rect 31392 29990 31444 29996
rect 31024 29028 31076 29034
rect 31024 28970 31076 28976
rect 31208 28076 31260 28082
rect 31208 28018 31260 28024
rect 31024 27872 31076 27878
rect 31024 27814 31076 27820
rect 31036 27470 31064 27814
rect 31116 27532 31168 27538
rect 31116 27474 31168 27480
rect 31024 27464 31076 27470
rect 31024 27406 31076 27412
rect 31128 27062 31156 27474
rect 31024 27056 31076 27062
rect 31024 26998 31076 27004
rect 31116 27056 31168 27062
rect 31116 26998 31168 27004
rect 31036 26790 31064 26998
rect 31220 26994 31248 28018
rect 31312 27402 31340 29974
rect 31404 29646 31432 29990
rect 31392 29640 31444 29646
rect 31392 29582 31444 29588
rect 31404 29170 31432 29582
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 31404 28626 31432 29106
rect 31496 28762 31524 33238
rect 31576 32020 31628 32026
rect 31576 31962 31628 31968
rect 31588 31929 31616 31962
rect 31574 31920 31630 31929
rect 31574 31855 31630 31864
rect 31576 31816 31628 31822
rect 31576 31758 31628 31764
rect 31588 31482 31616 31758
rect 31576 31476 31628 31482
rect 31576 31418 31628 31424
rect 31680 31362 31708 34054
rect 31772 33930 31800 34886
rect 33336 34678 33364 35974
rect 33428 35834 33456 36110
rect 33704 35834 33732 47126
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 36268 45280 36320 45286
rect 36268 45222 36320 45228
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 33416 35828 33468 35834
rect 33416 35770 33468 35776
rect 33692 35828 33744 35834
rect 33692 35770 33744 35776
rect 33508 35624 33560 35630
rect 33508 35566 33560 35572
rect 33416 35556 33468 35562
rect 33416 35498 33468 35504
rect 33324 34672 33376 34678
rect 33324 34614 33376 34620
rect 31760 33924 31812 33930
rect 31760 33866 31812 33872
rect 32680 33924 32732 33930
rect 32680 33866 32732 33872
rect 32220 33856 32272 33862
rect 32220 33798 32272 33804
rect 32232 33522 32260 33798
rect 32692 33658 32720 33866
rect 32680 33652 32732 33658
rect 32680 33594 32732 33600
rect 32220 33516 32272 33522
rect 32220 33458 32272 33464
rect 32496 33516 32548 33522
rect 32496 33458 32548 33464
rect 32508 33114 32536 33458
rect 33048 33380 33100 33386
rect 33048 33322 33100 33328
rect 32312 33108 32364 33114
rect 32312 33050 32364 33056
rect 32496 33108 32548 33114
rect 32496 33050 32548 33056
rect 32324 32434 32352 33050
rect 32864 33040 32916 33046
rect 32864 32982 32916 32988
rect 32496 32904 32548 32910
rect 32496 32846 32548 32852
rect 32312 32428 32364 32434
rect 32312 32370 32364 32376
rect 31850 31920 31906 31929
rect 31850 31855 31906 31864
rect 31588 31346 31708 31362
rect 31576 31340 31708 31346
rect 31628 31334 31708 31340
rect 31576 31282 31628 31288
rect 31588 30598 31616 31282
rect 31576 30592 31628 30598
rect 31576 30534 31628 30540
rect 31588 30394 31616 30534
rect 31576 30388 31628 30394
rect 31576 30330 31628 30336
rect 31668 30048 31720 30054
rect 31668 29990 31720 29996
rect 31680 29866 31708 29990
rect 31588 29838 31708 29866
rect 31588 29714 31616 29838
rect 31576 29708 31628 29714
rect 31576 29650 31628 29656
rect 31484 28756 31536 28762
rect 31484 28698 31536 28704
rect 31392 28620 31444 28626
rect 31392 28562 31444 28568
rect 31392 28416 31444 28422
rect 31392 28358 31444 28364
rect 31404 28082 31432 28358
rect 31496 28082 31524 28698
rect 31576 28552 31628 28558
rect 31628 28512 31708 28540
rect 31576 28494 31628 28500
rect 31392 28076 31444 28082
rect 31392 28018 31444 28024
rect 31484 28076 31536 28082
rect 31484 28018 31536 28024
rect 31484 27940 31536 27946
rect 31484 27882 31536 27888
rect 31300 27396 31352 27402
rect 31300 27338 31352 27344
rect 31300 27124 31352 27130
rect 31300 27066 31352 27072
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 31024 26784 31076 26790
rect 31024 26726 31076 26732
rect 31024 26444 31076 26450
rect 31024 26386 31076 26392
rect 31036 25702 31064 26386
rect 31312 26042 31340 27066
rect 31392 26580 31444 26586
rect 31392 26522 31444 26528
rect 31404 26450 31432 26522
rect 31392 26444 31444 26450
rect 31392 26386 31444 26392
rect 31300 26036 31352 26042
rect 31300 25978 31352 25984
rect 31392 25968 31444 25974
rect 31392 25910 31444 25916
rect 31024 25696 31076 25702
rect 31024 25638 31076 25644
rect 31208 25356 31260 25362
rect 31208 25298 31260 25304
rect 31220 24886 31248 25298
rect 31208 24880 31260 24886
rect 31208 24822 31260 24828
rect 31300 24812 31352 24818
rect 31300 24754 31352 24760
rect 31312 23866 31340 24754
rect 31404 24614 31432 25910
rect 31496 25838 31524 27882
rect 31680 27470 31708 28512
rect 31668 27464 31720 27470
rect 31668 27406 31720 27412
rect 31864 27402 31892 31855
rect 32324 31822 32352 32370
rect 32508 32366 32536 32846
rect 32876 32502 32904 32982
rect 33060 32910 33088 33322
rect 33140 33312 33192 33318
rect 33140 33254 33192 33260
rect 33324 33312 33376 33318
rect 33324 33254 33376 33260
rect 33152 32978 33180 33254
rect 33140 32972 33192 32978
rect 33140 32914 33192 32920
rect 33048 32904 33100 32910
rect 33048 32846 33100 32852
rect 33060 32774 33088 32846
rect 32956 32768 33008 32774
rect 32956 32710 33008 32716
rect 33048 32768 33100 32774
rect 33048 32710 33100 32716
rect 32968 32586 32996 32710
rect 32968 32558 33180 32586
rect 32864 32496 32916 32502
rect 32864 32438 32916 32444
rect 32496 32360 32548 32366
rect 32496 32302 32548 32308
rect 32680 31952 32732 31958
rect 32494 31920 32550 31929
rect 32680 31894 32732 31900
rect 32494 31855 32550 31864
rect 32508 31822 32536 31855
rect 32692 31822 32720 31894
rect 32312 31816 32364 31822
rect 32312 31758 32364 31764
rect 32496 31816 32548 31822
rect 32496 31758 32548 31764
rect 32680 31816 32732 31822
rect 32680 31758 32732 31764
rect 32324 31482 32352 31758
rect 32312 31476 32364 31482
rect 32312 31418 32364 31424
rect 32312 30660 32364 30666
rect 32312 30602 32364 30608
rect 32220 30592 32272 30598
rect 32220 30534 32272 30540
rect 32232 30326 32260 30534
rect 32220 30320 32272 30326
rect 32220 30262 32272 30268
rect 32036 29640 32088 29646
rect 32036 29582 32088 29588
rect 32048 28558 32076 29582
rect 32324 29306 32352 30602
rect 32404 29640 32456 29646
rect 32404 29582 32456 29588
rect 32416 29306 32444 29582
rect 32312 29300 32364 29306
rect 32312 29242 32364 29248
rect 32404 29300 32456 29306
rect 32404 29242 32456 29248
rect 32036 28552 32088 28558
rect 32036 28494 32088 28500
rect 32324 28150 32352 29242
rect 32312 28144 32364 28150
rect 32312 28086 32364 28092
rect 31944 27464 31996 27470
rect 31944 27406 31996 27412
rect 31852 27396 31904 27402
rect 31852 27338 31904 27344
rect 31576 26920 31628 26926
rect 31576 26862 31628 26868
rect 31588 26586 31616 26862
rect 31576 26580 31628 26586
rect 31576 26522 31628 26528
rect 31588 25906 31616 26522
rect 31576 25900 31628 25906
rect 31576 25842 31628 25848
rect 31484 25832 31536 25838
rect 31484 25774 31536 25780
rect 31496 25702 31524 25774
rect 31484 25696 31536 25702
rect 31484 25638 31536 25644
rect 31392 24608 31444 24614
rect 31392 24550 31444 24556
rect 31404 24138 31432 24550
rect 31496 24206 31524 25638
rect 31588 25498 31616 25842
rect 31576 25492 31628 25498
rect 31576 25434 31628 25440
rect 31850 25256 31906 25265
rect 31576 25220 31628 25226
rect 31850 25191 31906 25200
rect 31576 25162 31628 25168
rect 31484 24200 31536 24206
rect 31484 24142 31536 24148
rect 31392 24132 31444 24138
rect 31392 24074 31444 24080
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31024 23724 31076 23730
rect 31024 23666 31076 23672
rect 31036 23526 31064 23666
rect 31024 23520 31076 23526
rect 31024 23462 31076 23468
rect 31392 23520 31444 23526
rect 31392 23462 31444 23468
rect 30932 23112 30984 23118
rect 30932 23054 30984 23060
rect 31208 22976 31260 22982
rect 31208 22918 31260 22924
rect 31220 22710 31248 22918
rect 31404 22710 31432 23462
rect 31496 23186 31524 24142
rect 31588 23322 31616 25162
rect 31864 25158 31892 25191
rect 31852 25152 31904 25158
rect 31852 25094 31904 25100
rect 31956 24834 31984 27406
rect 32496 26988 32548 26994
rect 32496 26930 32548 26936
rect 32508 26518 32536 26930
rect 32496 26512 32548 26518
rect 32496 26454 32548 26460
rect 32508 25294 32536 26454
rect 32588 26308 32640 26314
rect 32588 26250 32640 26256
rect 32600 26042 32628 26250
rect 32588 26036 32640 26042
rect 32588 25978 32640 25984
rect 32496 25288 32548 25294
rect 32496 25230 32548 25236
rect 31956 24806 32076 24834
rect 31576 23316 31628 23322
rect 31576 23258 31628 23264
rect 31484 23180 31536 23186
rect 31484 23122 31536 23128
rect 31576 23112 31628 23118
rect 31576 23054 31628 23060
rect 31588 22778 31616 23054
rect 31576 22772 31628 22778
rect 31576 22714 31628 22720
rect 31208 22704 31260 22710
rect 31208 22646 31260 22652
rect 31392 22704 31444 22710
rect 31392 22646 31444 22652
rect 31944 22228 31996 22234
rect 31944 22170 31996 22176
rect 30852 22066 30972 22094
rect 30288 20868 30340 20874
rect 30288 20810 30340 20816
rect 30196 20800 30248 20806
rect 30196 20742 30248 20748
rect 30208 20380 30236 20742
rect 30300 20534 30328 20810
rect 30288 20528 30340 20534
rect 30288 20470 30340 20476
rect 30208 20352 30328 20380
rect 30196 20256 30248 20262
rect 30196 20198 30248 20204
rect 30208 19922 30236 20198
rect 30196 19916 30248 19922
rect 30196 19858 30248 19864
rect 30300 18698 30328 20352
rect 30288 18692 30340 18698
rect 30288 18634 30340 18640
rect 30196 18624 30248 18630
rect 30196 18566 30248 18572
rect 30208 17746 30236 18566
rect 30380 18080 30432 18086
rect 30380 18022 30432 18028
rect 30392 17746 30420 18022
rect 30196 17740 30248 17746
rect 30196 17682 30248 17688
rect 30380 17740 30432 17746
rect 30380 17682 30432 17688
rect 30944 3942 30972 22066
rect 31852 21344 31904 21350
rect 31852 21286 31904 21292
rect 31206 21040 31262 21049
rect 31206 20975 31208 20984
rect 31260 20975 31262 20984
rect 31208 20946 31260 20952
rect 31864 20874 31892 21286
rect 31852 20868 31904 20874
rect 31852 20810 31904 20816
rect 31208 20460 31260 20466
rect 31208 20402 31260 20408
rect 31116 18692 31168 18698
rect 31116 18634 31168 18640
rect 31128 18290 31156 18634
rect 31116 18284 31168 18290
rect 31116 18226 31168 18232
rect 31116 17128 31168 17134
rect 31116 17070 31168 17076
rect 30932 3936 30984 3942
rect 30932 3878 30984 3884
rect 31128 3738 31156 17070
rect 31220 14550 31248 20402
rect 31668 19916 31720 19922
rect 31668 19858 31720 19864
rect 31680 19825 31708 19858
rect 31666 19816 31722 19825
rect 31666 19751 31722 19760
rect 31956 18698 31984 22170
rect 31944 18692 31996 18698
rect 31944 18634 31996 18640
rect 31208 14544 31260 14550
rect 31208 14486 31260 14492
rect 30932 3732 30984 3738
rect 30932 3674 30984 3680
rect 31116 3732 31168 3738
rect 31116 3674 31168 3680
rect 30104 2576 30156 2582
rect 30104 2518 30156 2524
rect 29736 2372 29788 2378
rect 29736 2314 29788 2320
rect 30944 800 30972 3674
rect 32048 2106 32076 24806
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 32126 21040 32182 21049
rect 32126 20975 32128 20984
rect 32180 20975 32182 20984
rect 32128 20946 32180 20952
rect 32324 20602 32352 21490
rect 32312 20596 32364 20602
rect 32312 20538 32364 20544
rect 32312 20256 32364 20262
rect 32312 20198 32364 20204
rect 32128 18692 32180 18698
rect 32128 18634 32180 18640
rect 32140 17746 32168 18634
rect 32128 17740 32180 17746
rect 32128 17682 32180 17688
rect 32220 3120 32272 3126
rect 32220 3062 32272 3068
rect 32036 2100 32088 2106
rect 32036 2042 32088 2048
rect 32232 800 32260 3062
rect 32324 2650 32352 20198
rect 32692 3942 32720 31758
rect 33152 29646 33180 32558
rect 33336 32434 33364 33254
rect 33324 32428 33376 32434
rect 33324 32370 33376 32376
rect 33232 31952 33284 31958
rect 33232 31894 33284 31900
rect 33244 31278 33272 31894
rect 33232 31272 33284 31278
rect 33232 31214 33284 31220
rect 33324 30252 33376 30258
rect 33324 30194 33376 30200
rect 33336 29714 33364 30194
rect 33324 29708 33376 29714
rect 33324 29650 33376 29656
rect 33140 29640 33192 29646
rect 33140 29582 33192 29588
rect 33152 27062 33180 29582
rect 33324 29572 33376 29578
rect 33324 29514 33376 29520
rect 33232 28008 33284 28014
rect 33232 27950 33284 27956
rect 33244 27606 33272 27950
rect 33232 27600 33284 27606
rect 33232 27542 33284 27548
rect 33140 27056 33192 27062
rect 33140 26998 33192 27004
rect 32956 26920 33008 26926
rect 33336 26874 33364 29514
rect 33428 28490 33456 35498
rect 33520 35290 33548 35566
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 33508 35284 33560 35290
rect 33508 35226 33560 35232
rect 34612 35080 34664 35086
rect 34612 35022 34664 35028
rect 34624 34542 34652 35022
rect 34796 34672 34848 34678
rect 34796 34614 34848 34620
rect 34612 34536 34664 34542
rect 34612 34478 34664 34484
rect 33508 32904 33560 32910
rect 33508 32846 33560 32852
rect 33520 31414 33548 32846
rect 33784 32836 33836 32842
rect 33784 32778 33836 32784
rect 33796 31686 33824 32778
rect 34428 32768 34480 32774
rect 34428 32710 34480 32716
rect 34440 32434 34468 32710
rect 34428 32428 34480 32434
rect 34428 32370 34480 32376
rect 34520 32428 34572 32434
rect 34520 32370 34572 32376
rect 34532 32298 34560 32370
rect 34520 32292 34572 32298
rect 34520 32234 34572 32240
rect 33784 31680 33836 31686
rect 33784 31622 33836 31628
rect 33508 31408 33560 31414
rect 33508 31350 33560 31356
rect 33520 30326 33548 31350
rect 33796 30734 33824 31622
rect 34532 30802 34560 32234
rect 34520 30796 34572 30802
rect 34520 30738 34572 30744
rect 33784 30728 33836 30734
rect 33784 30670 33836 30676
rect 34520 30660 34572 30666
rect 34520 30602 34572 30608
rect 34152 30592 34204 30598
rect 34152 30534 34204 30540
rect 33508 30320 33560 30326
rect 33508 30262 33560 30268
rect 34164 30258 34192 30534
rect 34152 30252 34204 30258
rect 34152 30194 34204 30200
rect 34164 30054 34192 30194
rect 34244 30184 34296 30190
rect 34244 30126 34296 30132
rect 34152 30048 34204 30054
rect 34152 29990 34204 29996
rect 34164 29102 34192 29990
rect 34256 29170 34284 30126
rect 34428 30048 34480 30054
rect 34428 29990 34480 29996
rect 34440 29578 34468 29990
rect 34532 29646 34560 30602
rect 34624 29646 34652 34478
rect 34808 34202 34836 34614
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34796 34196 34848 34202
rect 34796 34138 34848 34144
rect 35348 33992 35400 33998
rect 35348 33934 35400 33940
rect 35360 33522 35388 33934
rect 35348 33516 35400 33522
rect 35348 33458 35400 33464
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34980 32972 35032 32978
rect 34980 32914 35032 32920
rect 34992 32434 35020 32914
rect 35072 32836 35124 32842
rect 35072 32778 35124 32784
rect 35084 32502 35112 32778
rect 35072 32496 35124 32502
rect 35072 32438 35124 32444
rect 34980 32428 35032 32434
rect 34980 32370 35032 32376
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 35360 31890 35388 33458
rect 35992 33312 36044 33318
rect 35992 33254 36044 33260
rect 36004 32842 36032 33254
rect 35992 32836 36044 32842
rect 35992 32778 36044 32784
rect 35440 32428 35492 32434
rect 35440 32370 35492 32376
rect 35348 31884 35400 31890
rect 35348 31826 35400 31832
rect 34796 31816 34848 31822
rect 34796 31758 34848 31764
rect 34808 31414 34836 31758
rect 34796 31408 34848 31414
rect 34796 31350 34848 31356
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 35164 30728 35216 30734
rect 35164 30670 35216 30676
rect 35176 30394 35204 30670
rect 35256 30592 35308 30598
rect 35256 30534 35308 30540
rect 35164 30388 35216 30394
rect 35164 30330 35216 30336
rect 35268 30326 35296 30534
rect 35256 30320 35308 30326
rect 35256 30262 35308 30268
rect 34796 30116 34848 30122
rect 34796 30058 34848 30064
rect 34808 29850 34836 30058
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34704 29844 34756 29850
rect 34704 29786 34756 29792
rect 34796 29844 34848 29850
rect 34796 29786 34848 29792
rect 34520 29640 34572 29646
rect 34520 29582 34572 29588
rect 34612 29640 34664 29646
rect 34612 29582 34664 29588
rect 34428 29572 34480 29578
rect 34428 29514 34480 29520
rect 34520 29504 34572 29510
rect 34520 29446 34572 29452
rect 34532 29238 34560 29446
rect 34520 29232 34572 29238
rect 34520 29174 34572 29180
rect 34244 29164 34296 29170
rect 34244 29106 34296 29112
rect 34152 29096 34204 29102
rect 34152 29038 34204 29044
rect 33508 28960 33560 28966
rect 33508 28902 33560 28908
rect 33520 28762 33548 28902
rect 33508 28756 33560 28762
rect 33508 28698 33560 28704
rect 33968 28756 34020 28762
rect 33968 28698 34020 28704
rect 33416 28484 33468 28490
rect 33416 28426 33468 28432
rect 33508 28484 33560 28490
rect 33508 28426 33560 28432
rect 33520 27674 33548 28426
rect 33508 27668 33560 27674
rect 33508 27610 33560 27616
rect 33876 27668 33928 27674
rect 33876 27610 33928 27616
rect 33508 27056 33560 27062
rect 33508 26998 33560 27004
rect 33416 26988 33468 26994
rect 33416 26930 33468 26936
rect 32956 26862 33008 26868
rect 32968 25158 32996 26862
rect 33152 26846 33364 26874
rect 33048 25764 33100 25770
rect 33048 25706 33100 25712
rect 32956 25152 33008 25158
rect 32956 25094 33008 25100
rect 32968 24954 32996 25094
rect 32956 24948 33008 24954
rect 32956 24890 33008 24896
rect 33060 24682 33088 25706
rect 33048 24676 33100 24682
rect 33048 24618 33100 24624
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 32876 23866 32904 24142
rect 32864 23860 32916 23866
rect 32864 23802 32916 23808
rect 33152 23633 33180 26846
rect 33324 26784 33376 26790
rect 33324 26726 33376 26732
rect 33336 26382 33364 26726
rect 33428 26450 33456 26930
rect 33416 26444 33468 26450
rect 33416 26386 33468 26392
rect 33520 26382 33548 26998
rect 33692 26444 33744 26450
rect 33692 26386 33744 26392
rect 33324 26376 33376 26382
rect 33324 26318 33376 26324
rect 33508 26376 33560 26382
rect 33508 26318 33560 26324
rect 33600 26376 33652 26382
rect 33600 26318 33652 26324
rect 33612 26042 33640 26318
rect 33600 26036 33652 26042
rect 33600 25978 33652 25984
rect 33232 23792 33284 23798
rect 33232 23734 33284 23740
rect 33138 23624 33194 23633
rect 33138 23559 33194 23568
rect 33244 22642 33272 23734
rect 33416 23044 33468 23050
rect 33416 22986 33468 22992
rect 33428 22778 33456 22986
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33232 22636 33284 22642
rect 33232 22578 33284 22584
rect 32680 3936 32732 3942
rect 32680 3878 32732 3884
rect 32864 3732 32916 3738
rect 32864 3674 32916 3680
rect 32876 3398 32904 3674
rect 32864 3392 32916 3398
rect 32864 3334 32916 3340
rect 33140 3392 33192 3398
rect 33140 3334 33192 3340
rect 33152 3126 33180 3334
rect 33140 3120 33192 3126
rect 33140 3062 33192 3068
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 32312 2644 32364 2650
rect 32312 2586 32364 2592
rect 33520 800 33548 2926
rect 33704 2514 33732 26386
rect 33888 25922 33916 27610
rect 33980 26994 34008 28698
rect 34612 28552 34664 28558
rect 34716 28506 34744 29786
rect 34888 29708 34940 29714
rect 34888 29650 34940 29656
rect 34900 29306 34928 29650
rect 34888 29300 34940 29306
rect 34888 29242 34940 29248
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 35360 28762 35388 31826
rect 35452 30734 35480 32370
rect 35808 30864 35860 30870
rect 35808 30806 35860 30812
rect 35440 30728 35492 30734
rect 35440 30670 35492 30676
rect 35820 29646 35848 30806
rect 35900 30320 35952 30326
rect 35900 30262 35952 30268
rect 35912 29850 35940 30262
rect 35900 29844 35952 29850
rect 35900 29786 35952 29792
rect 35808 29640 35860 29646
rect 35808 29582 35860 29588
rect 35532 29232 35584 29238
rect 35532 29174 35584 29180
rect 35544 28762 35572 29174
rect 35348 28756 35400 28762
rect 35348 28698 35400 28704
rect 35532 28756 35584 28762
rect 35532 28698 35584 28704
rect 35360 28558 35388 28698
rect 34664 28500 34744 28506
rect 34612 28494 34744 28500
rect 35348 28552 35400 28558
rect 35348 28494 35400 28500
rect 34624 28478 34744 28494
rect 34716 28014 34744 28478
rect 35360 28082 35388 28494
rect 35348 28076 35400 28082
rect 35348 28018 35400 28024
rect 34704 28008 34756 28014
rect 34704 27950 34756 27956
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 33968 26988 34020 26994
rect 33968 26930 34020 26936
rect 33980 26382 34008 26930
rect 34704 26784 34756 26790
rect 34704 26726 34756 26732
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 34060 26240 34112 26246
rect 34060 26182 34112 26188
rect 34072 25974 34100 26182
rect 34060 25968 34112 25974
rect 33784 25900 33836 25906
rect 33888 25894 34008 25922
rect 34060 25910 34112 25916
rect 34612 25968 34664 25974
rect 34612 25910 34664 25916
rect 33784 25842 33836 25848
rect 33796 25294 33824 25842
rect 33876 25832 33928 25838
rect 33876 25774 33928 25780
rect 33888 25362 33916 25774
rect 33876 25356 33928 25362
rect 33876 25298 33928 25304
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 33796 24818 33824 25230
rect 33784 24812 33836 24818
rect 33784 24754 33836 24760
rect 33796 23866 33824 24754
rect 33784 23860 33836 23866
rect 33784 23802 33836 23808
rect 33980 23730 34008 25894
rect 34242 25528 34298 25537
rect 34242 25463 34244 25472
rect 34296 25463 34298 25472
rect 34244 25434 34296 25440
rect 34624 25430 34652 25910
rect 34612 25424 34664 25430
rect 34612 25366 34664 25372
rect 34716 25226 34744 26726
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34704 25220 34756 25226
rect 34704 25162 34756 25168
rect 35992 25220 36044 25226
rect 35992 25162 36044 25168
rect 35716 24880 35768 24886
rect 35716 24822 35768 24828
rect 35728 24682 35756 24822
rect 36004 24818 36032 25162
rect 35992 24812 36044 24818
rect 35992 24754 36044 24760
rect 35716 24676 35768 24682
rect 35716 24618 35768 24624
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 36280 24410 36308 45222
rect 37096 36236 37148 36242
rect 37096 36178 37148 36184
rect 36360 24608 36412 24614
rect 36360 24550 36412 24556
rect 36268 24404 36320 24410
rect 36268 24346 36320 24352
rect 36176 24064 36228 24070
rect 36176 24006 36228 24012
rect 33968 23724 34020 23730
rect 33968 23666 34020 23672
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 36188 23186 36216 24006
rect 36280 23798 36308 24346
rect 36372 24206 36400 24550
rect 37108 24274 37136 36178
rect 37096 24268 37148 24274
rect 37096 24210 37148 24216
rect 36360 24200 36412 24206
rect 37292 24177 37320 47654
rect 37372 47524 37424 47530
rect 37372 47466 37424 47472
rect 36360 24142 36412 24148
rect 37278 24168 37334 24177
rect 36268 23792 36320 23798
rect 36268 23734 36320 23740
rect 36176 23180 36228 23186
rect 36176 23122 36228 23128
rect 35992 23112 36044 23118
rect 35992 23054 36044 23060
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34152 22024 34204 22030
rect 34152 21966 34204 21972
rect 34518 21992 34574 22001
rect 34164 21690 34192 21966
rect 34518 21927 34574 21936
rect 34152 21684 34204 21690
rect 34152 21626 34204 21632
rect 33784 21548 33836 21554
rect 33784 21490 33836 21496
rect 33796 20874 33824 21490
rect 34532 21486 34560 21927
rect 34704 21888 34756 21894
rect 34704 21830 34756 21836
rect 34716 21622 34744 21830
rect 34704 21616 34756 21622
rect 34704 21558 34756 21564
rect 34520 21480 34572 21486
rect 34520 21422 34572 21428
rect 35900 21412 35952 21418
rect 35900 21354 35952 21360
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35912 20942 35940 21354
rect 35900 20936 35952 20942
rect 35900 20878 35952 20884
rect 33784 20868 33836 20874
rect 33784 20810 33836 20816
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 36004 19718 36032 23054
rect 35992 19712 36044 19718
rect 35992 19654 36044 19660
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 36280 18970 36308 23734
rect 36372 23730 36400 24142
rect 37278 24103 37334 24112
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 36372 22642 36400 23666
rect 36360 22636 36412 22642
rect 36360 22578 36412 22584
rect 36636 22568 36688 22574
rect 36636 22510 36688 22516
rect 36360 20868 36412 20874
rect 36360 20810 36412 20816
rect 36268 18964 36320 18970
rect 36268 18906 36320 18912
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 36176 8288 36228 8294
rect 36176 8230 36228 8236
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 36188 8090 36216 8230
rect 36176 8084 36228 8090
rect 36176 8026 36228 8032
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 33784 3664 33836 3670
rect 34060 3664 34112 3670
rect 33836 3612 34060 3618
rect 33784 3606 34112 3612
rect 33796 3590 34100 3606
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 33888 2922 33916 3470
rect 33876 2916 33928 2922
rect 33876 2858 33928 2864
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 36372 2650 36400 20810
rect 36648 10674 36676 22510
rect 36636 10668 36688 10674
rect 36636 10610 36688 10616
rect 37384 5166 37412 47466
rect 38200 47456 38252 47462
rect 38200 47398 38252 47404
rect 38212 47258 38240 47398
rect 38200 47252 38252 47258
rect 38200 47194 38252 47200
rect 38200 47048 38252 47054
rect 38200 46990 38252 46996
rect 38212 46578 38240 46990
rect 38200 46572 38252 46578
rect 38200 46514 38252 46520
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 38384 46504 38436 46510
rect 38384 46446 38436 46452
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 38396 46170 38424 46446
rect 38384 46164 38436 46170
rect 38384 46106 38436 46112
rect 39960 45554 39988 49200
rect 40788 47410 40816 49286
rect 41206 49200 41318 49286
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 43782 49200 43894 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49200 46470 50000
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 39868 45526 39988 45554
rect 40052 47382 40816 47410
rect 39868 45422 39896 45526
rect 38660 45416 38712 45422
rect 38660 45358 38712 45364
rect 38844 45416 38896 45422
rect 38844 45358 38896 45364
rect 39856 45416 39908 45422
rect 39856 45358 39908 45364
rect 38672 44742 38700 45358
rect 38752 45348 38804 45354
rect 38752 45290 38804 45296
rect 38764 44878 38792 45290
rect 38856 45082 38884 45358
rect 38844 45076 38896 45082
rect 38844 45018 38896 45024
rect 38752 44872 38804 44878
rect 38752 44814 38804 44820
rect 38660 44736 38712 44742
rect 38660 44678 38712 44684
rect 38764 24206 38792 44814
rect 40052 24857 40080 47382
rect 40500 47252 40552 47258
rect 40500 47194 40552 47200
rect 40408 46980 40460 46986
rect 40408 46922 40460 46928
rect 40316 45960 40368 45966
rect 40316 45902 40368 45908
rect 40132 39432 40184 39438
rect 40132 39374 40184 39380
rect 40144 38962 40172 39374
rect 40132 38956 40184 38962
rect 40132 38898 40184 38904
rect 40144 38282 40172 38898
rect 40328 38894 40356 45902
rect 40316 38888 40368 38894
rect 40316 38830 40368 38836
rect 40132 38276 40184 38282
rect 40132 38218 40184 38224
rect 40144 37874 40172 38218
rect 40132 37868 40184 37874
rect 40132 37810 40184 37816
rect 40144 37262 40172 37810
rect 40132 37256 40184 37262
rect 40132 37198 40184 37204
rect 40316 37188 40368 37194
rect 40316 37130 40368 37136
rect 40328 36922 40356 37130
rect 40316 36916 40368 36922
rect 40316 36858 40368 36864
rect 40420 26926 40448 46922
rect 40408 26920 40460 26926
rect 40408 26862 40460 26868
rect 40038 24848 40094 24857
rect 40038 24783 40094 24792
rect 40040 24744 40092 24750
rect 40040 24686 40092 24692
rect 40316 24744 40368 24750
rect 40316 24686 40368 24692
rect 40408 24744 40460 24750
rect 40408 24686 40460 24692
rect 40052 24342 40080 24686
rect 40040 24336 40092 24342
rect 40040 24278 40092 24284
rect 40328 24206 40356 24686
rect 38752 24200 38804 24206
rect 38752 24142 38804 24148
rect 40316 24200 40368 24206
rect 40316 24142 40368 24148
rect 37648 23792 37700 23798
rect 37648 23734 37700 23740
rect 37660 17338 37688 23734
rect 40420 23594 40448 24686
rect 40408 23588 40460 23594
rect 40408 23530 40460 23536
rect 40408 23112 40460 23118
rect 40408 23054 40460 23060
rect 40420 22778 40448 23054
rect 40408 22772 40460 22778
rect 40408 22714 40460 22720
rect 40316 22636 40368 22642
rect 40316 22578 40368 22584
rect 40328 22030 40356 22578
rect 40512 22438 40540 47194
rect 41892 46918 41920 49200
rect 41880 46912 41932 46918
rect 41880 46854 41932 46860
rect 41420 46368 41472 46374
rect 41420 46310 41472 46316
rect 41432 46034 41460 46310
rect 42536 46034 42564 49200
rect 42708 47048 42760 47054
rect 42708 46990 42760 46996
rect 42720 46578 42748 46990
rect 42892 46912 42944 46918
rect 42892 46854 42944 46860
rect 42708 46572 42760 46578
rect 42708 46514 42760 46520
rect 41420 46028 41472 46034
rect 41420 45970 41472 45976
rect 42524 46028 42576 46034
rect 42524 45970 42576 45976
rect 41604 45892 41656 45898
rect 41604 45834 41656 45840
rect 41616 45558 41644 45834
rect 41604 45552 41656 45558
rect 41604 45494 41656 45500
rect 40960 45484 41012 45490
rect 40960 45426 41012 45432
rect 40972 39506 41000 45426
rect 41420 45280 41472 45286
rect 41420 45222 41472 45228
rect 41432 44946 41460 45222
rect 42904 44946 42932 46854
rect 43180 46646 43208 49200
rect 43824 47054 43852 49200
rect 44468 47122 44496 49200
rect 44456 47116 44508 47122
rect 44456 47058 44508 47064
rect 43812 47048 43864 47054
rect 43812 46990 43864 46996
rect 44364 46980 44416 46986
rect 44364 46922 44416 46928
rect 43352 46912 43404 46918
rect 43352 46854 43404 46860
rect 43168 46640 43220 46646
rect 43168 46582 43220 46588
rect 41420 44940 41472 44946
rect 41420 44882 41472 44888
rect 42892 44940 42944 44946
rect 42892 44882 42944 44888
rect 41604 44804 41656 44810
rect 41604 44746 41656 44752
rect 41616 44538 41644 44746
rect 41604 44532 41656 44538
rect 41604 44474 41656 44480
rect 40776 39500 40828 39506
rect 40776 39442 40828 39448
rect 40960 39500 41012 39506
rect 40960 39442 41012 39448
rect 40684 36916 40736 36922
rect 40684 36858 40736 36864
rect 40592 23724 40644 23730
rect 40592 23666 40644 23672
rect 40500 22432 40552 22438
rect 40500 22374 40552 22380
rect 40512 22030 40540 22374
rect 40316 22024 40368 22030
rect 40316 21966 40368 21972
rect 40500 22024 40552 22030
rect 40500 21966 40552 21972
rect 40328 21350 40356 21966
rect 40500 21888 40552 21894
rect 40500 21830 40552 21836
rect 40316 21344 40368 21350
rect 40316 21286 40368 21292
rect 40132 18284 40184 18290
rect 40132 18226 40184 18232
rect 40040 18148 40092 18154
rect 40040 18090 40092 18096
rect 40052 17338 40080 18090
rect 37648 17332 37700 17338
rect 37648 17274 37700 17280
rect 40040 17332 40092 17338
rect 40040 17274 40092 17280
rect 40144 17270 40172 18226
rect 40132 17264 40184 17270
rect 40132 17206 40184 17212
rect 40132 5704 40184 5710
rect 40132 5646 40184 5652
rect 40144 5370 40172 5646
rect 40224 5568 40276 5574
rect 40224 5510 40276 5516
rect 40132 5364 40184 5370
rect 40132 5306 40184 5312
rect 37464 5296 37516 5302
rect 37464 5238 37516 5244
rect 37372 5160 37424 5166
rect 37372 5102 37424 5108
rect 37280 4548 37332 4554
rect 37280 4490 37332 4496
rect 37292 4078 37320 4490
rect 37476 4282 37504 5238
rect 39212 5228 39264 5234
rect 39212 5170 39264 5176
rect 38476 5160 38528 5166
rect 38476 5102 38528 5108
rect 38488 4690 38516 5102
rect 39224 4826 39252 5170
rect 39212 4820 39264 4826
rect 39212 4762 39264 4768
rect 39304 4820 39356 4826
rect 39304 4762 39356 4768
rect 38476 4684 38528 4690
rect 38476 4626 38528 4632
rect 37556 4548 37608 4554
rect 37556 4490 37608 4496
rect 37464 4276 37516 4282
rect 37464 4218 37516 4224
rect 37280 4072 37332 4078
rect 37280 4014 37332 4020
rect 37464 3188 37516 3194
rect 37464 3130 37516 3136
rect 37476 2854 37504 3130
rect 37568 3058 37596 4490
rect 37740 4140 37792 4146
rect 37740 4082 37792 4088
rect 37752 3194 37780 4082
rect 39316 3738 39344 4762
rect 40236 4690 40264 5510
rect 40316 5364 40368 5370
rect 40316 5306 40368 5312
rect 40328 5166 40356 5306
rect 40316 5160 40368 5166
rect 40316 5102 40368 5108
rect 40408 5024 40460 5030
rect 40408 4966 40460 4972
rect 40420 4690 40448 4966
rect 40224 4684 40276 4690
rect 40224 4626 40276 4632
rect 40408 4684 40460 4690
rect 40408 4626 40460 4632
rect 40132 4616 40184 4622
rect 40132 4558 40184 4564
rect 40040 4208 40092 4214
rect 40040 4150 40092 4156
rect 39948 4072 40000 4078
rect 39948 4014 40000 4020
rect 39304 3732 39356 3738
rect 39304 3674 39356 3680
rect 39672 3460 39724 3466
rect 39672 3402 39724 3408
rect 39684 3194 39712 3402
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 39672 3188 39724 3194
rect 39672 3130 39724 3136
rect 39960 3074 39988 4014
rect 40052 3534 40080 4150
rect 40144 3738 40172 4558
rect 40512 4214 40540 21830
rect 40604 5370 40632 23666
rect 40696 17066 40724 36858
rect 40788 35894 40816 39442
rect 41328 38412 41380 38418
rect 41328 38354 41380 38360
rect 41340 35894 41368 38354
rect 40788 35866 41092 35894
rect 40868 24336 40920 24342
rect 40868 24278 40920 24284
rect 40880 23186 40908 24278
rect 40960 24268 41012 24274
rect 40960 24210 41012 24216
rect 40972 23866 41000 24210
rect 40960 23860 41012 23866
rect 40960 23802 41012 23808
rect 40868 23180 40920 23186
rect 40868 23122 40920 23128
rect 41064 20398 41092 35866
rect 41156 35866 41368 35894
rect 41156 32570 41184 35866
rect 41144 32564 41196 32570
rect 41144 32506 41196 32512
rect 41052 20392 41104 20398
rect 41052 20334 41104 20340
rect 40776 18284 40828 18290
rect 40776 18226 40828 18232
rect 40684 17060 40736 17066
rect 40684 17002 40736 17008
rect 40788 12434 40816 18226
rect 40960 18080 41012 18086
rect 40960 18022 41012 18028
rect 40972 17746 41000 18022
rect 40960 17740 41012 17746
rect 40960 17682 41012 17688
rect 40868 15496 40920 15502
rect 40868 15438 40920 15444
rect 40696 12406 40816 12434
rect 40592 5364 40644 5370
rect 40592 5306 40644 5312
rect 40592 5228 40644 5234
rect 40592 5170 40644 5176
rect 40604 4282 40632 5170
rect 40592 4276 40644 4282
rect 40592 4218 40644 4224
rect 40500 4208 40552 4214
rect 40500 4150 40552 4156
rect 40224 4140 40276 4146
rect 40224 4082 40276 4088
rect 40132 3732 40184 3738
rect 40132 3674 40184 3680
rect 40040 3528 40092 3534
rect 40040 3470 40092 3476
rect 37556 3052 37608 3058
rect 39960 3046 40080 3074
rect 37556 2994 37608 3000
rect 37372 2848 37424 2854
rect 37372 2790 37424 2796
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 35624 2644 35676 2650
rect 35624 2586 35676 2592
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 33692 2508 33744 2514
rect 33692 2450 33744 2456
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35452 800 35480 2382
rect 35636 2310 35664 2586
rect 35900 2576 35952 2582
rect 35900 2518 35952 2524
rect 35992 2576 36044 2582
rect 35992 2518 36044 2524
rect 35624 2304 35676 2310
rect 35624 2246 35676 2252
rect 35912 2106 35940 2518
rect 36004 2378 36032 2518
rect 35992 2372 36044 2378
rect 35992 2314 36044 2320
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 35900 2100 35952 2106
rect 35900 2042 35952 2048
rect 36096 800 36124 2314
rect 37384 1902 37412 2790
rect 37568 2774 37596 2994
rect 40052 2990 40080 3046
rect 39948 2984 40000 2990
rect 39948 2926 40000 2932
rect 40040 2984 40092 2990
rect 40040 2926 40092 2932
rect 37568 2746 37688 2774
rect 37660 2310 37688 2746
rect 38016 2372 38068 2378
rect 38016 2314 38068 2320
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 37648 2304 37700 2310
rect 37648 2246 37700 2252
rect 37372 1896 37424 1902
rect 37372 1838 37424 1844
rect 38028 800 38056 2314
rect 39316 800 39344 2314
rect 39960 800 39988 2926
rect 40236 2922 40264 4082
rect 40408 2984 40460 2990
rect 40408 2926 40460 2932
rect 40224 2916 40276 2922
rect 40224 2858 40276 2864
rect 40236 2446 40264 2858
rect 40420 2446 40448 2926
rect 40512 2582 40540 4150
rect 40592 3052 40644 3058
rect 40592 2994 40644 3000
rect 40604 2650 40632 2994
rect 40592 2644 40644 2650
rect 40592 2586 40644 2592
rect 40500 2576 40552 2582
rect 40500 2518 40552 2524
rect 40224 2440 40276 2446
rect 40224 2382 40276 2388
rect 40408 2440 40460 2446
rect 40408 2382 40460 2388
rect 40592 2440 40644 2446
rect 40592 2382 40644 2388
rect 40604 800 40632 2382
rect 40696 2106 40724 12406
rect 40880 5234 40908 15438
rect 40868 5228 40920 5234
rect 40868 5170 40920 5176
rect 40868 5024 40920 5030
rect 40868 4966 40920 4972
rect 40880 4826 40908 4966
rect 40868 4820 40920 4826
rect 40868 4762 40920 4768
rect 40776 3528 40828 3534
rect 40776 3470 40828 3476
rect 40788 3194 40816 3470
rect 41156 3398 41184 32506
rect 43364 25498 43392 46854
rect 43812 46504 43864 46510
rect 43812 46446 43864 46452
rect 43824 46170 43852 46446
rect 43812 46164 43864 46170
rect 43812 46106 43864 46112
rect 43812 45484 43864 45490
rect 43812 45426 43864 45432
rect 43444 45280 43496 45286
rect 43444 45222 43496 45228
rect 43352 25492 43404 25498
rect 43352 25434 43404 25440
rect 42892 24812 42944 24818
rect 42892 24754 42944 24760
rect 42524 24064 42576 24070
rect 42524 24006 42576 24012
rect 42536 23866 42564 24006
rect 42524 23860 42576 23866
rect 42524 23802 42576 23808
rect 42904 23662 42932 24754
rect 43456 24206 43484 45222
rect 43628 24812 43680 24818
rect 43628 24754 43680 24760
rect 43168 24200 43220 24206
rect 43168 24142 43220 24148
rect 43444 24200 43496 24206
rect 43444 24142 43496 24148
rect 43536 24200 43588 24206
rect 43536 24142 43588 24148
rect 43180 23866 43208 24142
rect 43168 23860 43220 23866
rect 43168 23802 43220 23808
rect 43352 23724 43404 23730
rect 43352 23666 43404 23672
rect 42892 23656 42944 23662
rect 42892 23598 42944 23604
rect 42904 23322 42932 23598
rect 42892 23316 42944 23322
rect 42892 23258 42944 23264
rect 42064 23180 42116 23186
rect 42064 23122 42116 23128
rect 42076 18698 42104 23122
rect 42800 22568 42852 22574
rect 42800 22510 42852 22516
rect 42812 22098 42840 22510
rect 42892 22500 42944 22506
rect 42892 22442 42944 22448
rect 42904 22166 42932 22442
rect 42892 22160 42944 22166
rect 42892 22102 42944 22108
rect 42800 22092 42852 22098
rect 42800 22034 42852 22040
rect 42616 22024 42668 22030
rect 42616 21966 42668 21972
rect 42984 22024 43036 22030
rect 42984 21966 43036 21972
rect 42628 21554 42656 21966
rect 42996 21622 43024 21966
rect 43364 21894 43392 23666
rect 43456 23118 43484 24142
rect 43444 23112 43496 23118
rect 43444 23054 43496 23060
rect 43548 23032 43576 24142
rect 43640 24070 43668 24754
rect 43824 24274 43852 45426
rect 44180 38888 44232 38894
rect 44180 38830 44232 38836
rect 44192 38350 44220 38830
rect 44180 38344 44232 38350
rect 44180 38286 44232 38292
rect 44376 30802 44404 46922
rect 45112 45626 45140 49200
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45100 45620 45152 45626
rect 45100 45562 45152 45568
rect 44456 45416 44508 45422
rect 44456 45358 44508 45364
rect 44468 45082 44496 45358
rect 44456 45076 44508 45082
rect 44456 45018 44508 45024
rect 45008 44872 45060 44878
rect 45008 44814 45060 44820
rect 45020 38418 45048 44814
rect 45204 43994 45232 46990
rect 45468 46980 45520 46986
rect 45468 46922 45520 46928
rect 45376 46504 45428 46510
rect 45376 46446 45428 46452
rect 45388 45082 45416 46446
rect 45480 45354 45508 46922
rect 45560 46436 45612 46442
rect 45560 46378 45612 46384
rect 45468 45348 45520 45354
rect 45468 45290 45520 45296
rect 45376 45076 45428 45082
rect 45376 45018 45428 45024
rect 45572 44402 45600 46378
rect 45756 45966 45784 49200
rect 46400 47410 46428 49200
rect 46400 47382 46888 47410
rect 45836 46028 45888 46034
rect 45836 45970 45888 45976
rect 46756 46028 46808 46034
rect 46756 45970 46808 45976
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 45848 44878 45876 45970
rect 45836 44872 45888 44878
rect 45836 44814 45888 44820
rect 46296 44872 46348 44878
rect 46296 44814 46348 44820
rect 45560 44396 45612 44402
rect 45560 44338 45612 44344
rect 45848 44198 45876 44814
rect 46308 44402 46336 44814
rect 46296 44396 46348 44402
rect 46296 44338 46348 44344
rect 45836 44192 45888 44198
rect 45836 44134 45888 44140
rect 46572 44192 46624 44198
rect 46572 44134 46624 44140
rect 45192 43988 45244 43994
rect 45192 43930 45244 43936
rect 46296 43784 46348 43790
rect 46296 43726 46348 43732
rect 46308 43314 46336 43726
rect 46296 43308 46348 43314
rect 46296 43250 46348 43256
rect 46296 42696 46348 42702
rect 46296 42638 46348 42644
rect 46308 42226 46336 42638
rect 46296 42220 46348 42226
rect 46296 42162 46348 42168
rect 46296 39840 46348 39846
rect 46296 39782 46348 39788
rect 45926 39536 45982 39545
rect 46308 39506 46336 39782
rect 45926 39471 45982 39480
rect 46296 39500 46348 39506
rect 45468 38888 45520 38894
rect 45468 38830 45520 38836
rect 45008 38412 45060 38418
rect 45008 38354 45060 38360
rect 44364 30796 44416 30802
rect 44364 30738 44416 30744
rect 45282 26344 45338 26353
rect 45282 26279 45338 26288
rect 44548 24812 44600 24818
rect 44548 24754 44600 24760
rect 44272 24744 44324 24750
rect 44272 24686 44324 24692
rect 43904 24608 43956 24614
rect 43904 24550 43956 24556
rect 43812 24268 43864 24274
rect 43812 24210 43864 24216
rect 43628 24064 43680 24070
rect 43628 24006 43680 24012
rect 43824 23474 43852 24210
rect 43916 23730 43944 24550
rect 44284 24410 44312 24686
rect 44272 24404 44324 24410
rect 44272 24346 44324 24352
rect 44560 24138 44588 24754
rect 44548 24132 44600 24138
rect 44548 24074 44600 24080
rect 43904 23724 43956 23730
rect 43904 23666 43956 23672
rect 43824 23446 44312 23474
rect 43628 23044 43680 23050
rect 43548 23004 43628 23032
rect 43628 22986 43680 22992
rect 43536 22500 43588 22506
rect 43536 22442 43588 22448
rect 43548 22030 43576 22442
rect 43536 22024 43588 22030
rect 43536 21966 43588 21972
rect 43352 21888 43404 21894
rect 43352 21830 43404 21836
rect 43548 21690 43576 21966
rect 43536 21684 43588 21690
rect 43536 21626 43588 21632
rect 42984 21616 43036 21622
rect 42984 21558 43036 21564
rect 42616 21548 42668 21554
rect 42616 21490 42668 21496
rect 42340 20936 42392 20942
rect 42340 20878 42392 20884
rect 42352 20466 42380 20878
rect 42340 20460 42392 20466
rect 42340 20402 42392 20408
rect 42064 18692 42116 18698
rect 42064 18634 42116 18640
rect 42076 18154 42104 18634
rect 42156 18216 42208 18222
rect 42156 18158 42208 18164
rect 42064 18148 42116 18154
rect 42064 18090 42116 18096
rect 42076 16574 42104 18090
rect 42168 17814 42196 18158
rect 42156 17808 42208 17814
rect 42156 17750 42208 17756
rect 42168 17678 42196 17750
rect 42156 17672 42208 17678
rect 42156 17614 42208 17620
rect 42076 16546 42196 16574
rect 42168 4554 42196 16546
rect 42352 6458 42380 20402
rect 42432 19848 42484 19854
rect 42432 19790 42484 19796
rect 42444 19378 42472 19790
rect 42432 19372 42484 19378
rect 42432 19314 42484 19320
rect 42444 17814 42472 19314
rect 42524 18284 42576 18290
rect 42524 18226 42576 18232
rect 42536 17882 42564 18226
rect 42524 17876 42576 17882
rect 42524 17818 42576 17824
rect 42432 17808 42484 17814
rect 42432 17750 42484 17756
rect 42524 17536 42576 17542
rect 42524 17478 42576 17484
rect 42536 17134 42564 17478
rect 42524 17128 42576 17134
rect 42524 17070 42576 17076
rect 42628 6914 42656 21490
rect 42708 21412 42760 21418
rect 42708 21354 42760 21360
rect 42720 21010 42748 21354
rect 42708 21004 42760 21010
rect 42708 20946 42760 20952
rect 42720 20466 42748 20946
rect 42708 20460 42760 20466
rect 42708 20402 42760 20408
rect 43352 20460 43404 20466
rect 43352 20402 43404 20408
rect 43364 19922 43392 20402
rect 43536 20392 43588 20398
rect 43536 20334 43588 20340
rect 43352 19916 43404 19922
rect 43352 19858 43404 19864
rect 43548 19514 43576 20334
rect 43536 19508 43588 19514
rect 43536 19450 43588 19456
rect 43260 18760 43312 18766
rect 43260 18702 43312 18708
rect 42708 17876 42760 17882
rect 42708 17818 42760 17824
rect 42720 17610 42748 17818
rect 43272 17678 43300 18702
rect 43260 17672 43312 17678
rect 43260 17614 43312 17620
rect 43444 17672 43496 17678
rect 43444 17614 43496 17620
rect 42708 17604 42760 17610
rect 42708 17546 42760 17552
rect 43168 17604 43220 17610
rect 43168 17546 43220 17552
rect 42720 17202 42748 17546
rect 43180 17270 43208 17546
rect 43456 17542 43484 17614
rect 43444 17536 43496 17542
rect 43444 17478 43496 17484
rect 43456 17338 43484 17478
rect 43444 17332 43496 17338
rect 43444 17274 43496 17280
rect 43168 17264 43220 17270
rect 43168 17206 43220 17212
rect 42708 17196 42760 17202
rect 42708 17138 42760 17144
rect 42444 6886 42656 6914
rect 42340 6452 42392 6458
rect 42340 6394 42392 6400
rect 42156 4548 42208 4554
rect 42156 4490 42208 4496
rect 41144 3392 41196 3398
rect 41144 3334 41196 3340
rect 40776 3188 40828 3194
rect 40776 3130 40828 3136
rect 41236 3052 41288 3058
rect 41236 2994 41288 3000
rect 40684 2100 40736 2106
rect 40684 2042 40736 2048
rect 41248 800 41276 2994
rect 42444 2582 42472 6886
rect 42524 5296 42576 5302
rect 42524 5238 42576 5244
rect 42536 4826 42564 5238
rect 43640 5166 43668 22986
rect 43720 22432 43772 22438
rect 43720 22374 43772 22380
rect 43732 21554 43760 22374
rect 43812 21956 43864 21962
rect 43812 21898 43864 21904
rect 43720 21548 43772 21554
rect 43720 21490 43772 21496
rect 43824 21486 43852 21898
rect 43812 21480 43864 21486
rect 43812 21422 43864 21428
rect 43824 19990 43852 21422
rect 43904 20936 43956 20942
rect 43904 20878 43956 20884
rect 44088 20936 44140 20942
rect 44088 20878 44140 20884
rect 43812 19984 43864 19990
rect 43812 19926 43864 19932
rect 43916 19922 43944 20878
rect 43996 20800 44048 20806
rect 43996 20742 44048 20748
rect 44008 20466 44036 20742
rect 44100 20602 44128 20878
rect 44088 20596 44140 20602
rect 44088 20538 44140 20544
rect 43996 20460 44048 20466
rect 43996 20402 44048 20408
rect 43904 19916 43956 19922
rect 43904 19858 43956 19864
rect 43904 19780 43956 19786
rect 43904 19722 43956 19728
rect 43916 19378 43944 19722
rect 43904 19372 43956 19378
rect 43904 19314 43956 19320
rect 43916 18766 43944 19314
rect 43904 18760 43956 18766
rect 43904 18702 43956 18708
rect 43812 18624 43864 18630
rect 43812 18566 43864 18572
rect 43824 18290 43852 18566
rect 43812 18284 43864 18290
rect 43812 18226 43864 18232
rect 43916 17882 43944 18702
rect 44180 18148 44232 18154
rect 44180 18090 44232 18096
rect 43904 17876 43956 17882
rect 43904 17818 43956 17824
rect 43720 17604 43772 17610
rect 43720 17546 43772 17552
rect 43732 17270 43760 17546
rect 43720 17264 43772 17270
rect 43720 17206 43772 17212
rect 44192 17134 44220 18090
rect 43904 17128 43956 17134
rect 43904 17070 43956 17076
rect 44180 17128 44232 17134
rect 44180 17070 44232 17076
rect 43916 16114 43944 17070
rect 44284 17066 44312 23446
rect 44272 17060 44324 17066
rect 44272 17002 44324 17008
rect 43904 16108 43956 16114
rect 43904 16050 43956 16056
rect 44088 16040 44140 16046
rect 44088 15982 44140 15988
rect 44100 15706 44128 15982
rect 44088 15700 44140 15706
rect 44088 15642 44140 15648
rect 44560 13938 44588 24074
rect 44732 23520 44784 23526
rect 44732 23462 44784 23468
rect 44744 21554 44772 23462
rect 45296 23254 45324 26279
rect 45480 25294 45508 38830
rect 45652 38820 45704 38826
rect 45652 38762 45704 38768
rect 45468 25288 45520 25294
rect 45468 25230 45520 25236
rect 45480 24886 45508 25230
rect 45560 25152 45612 25158
rect 45560 25094 45612 25100
rect 45468 24880 45520 24886
rect 45468 24822 45520 24828
rect 45572 24818 45600 25094
rect 45560 24812 45612 24818
rect 45560 24754 45612 24760
rect 45572 24274 45600 24754
rect 45560 24268 45612 24274
rect 45560 24210 45612 24216
rect 45376 23656 45428 23662
rect 45376 23598 45428 23604
rect 45560 23656 45612 23662
rect 45560 23598 45612 23604
rect 45388 23322 45416 23598
rect 45376 23316 45428 23322
rect 45376 23258 45428 23264
rect 45284 23248 45336 23254
rect 45284 23190 45336 23196
rect 45572 23186 45600 23598
rect 45560 23180 45612 23186
rect 45560 23122 45612 23128
rect 45560 23044 45612 23050
rect 45560 22986 45612 22992
rect 45572 22642 45600 22986
rect 45560 22636 45612 22642
rect 45560 22578 45612 22584
rect 44732 21548 44784 21554
rect 44732 21490 44784 21496
rect 44640 21480 44692 21486
rect 44640 21422 44692 21428
rect 44652 20466 44680 21422
rect 45572 20534 45600 22578
rect 45664 20942 45692 38762
rect 45836 25832 45888 25838
rect 45836 25774 45888 25780
rect 45744 24200 45796 24206
rect 45744 24142 45796 24148
rect 45756 23186 45784 24142
rect 45848 24138 45876 25774
rect 45940 24342 45968 39471
rect 46296 39442 46348 39448
rect 46296 38344 46348 38350
rect 46296 38286 46348 38292
rect 46308 37466 46336 38286
rect 46296 37460 46348 37466
rect 46296 37402 46348 37408
rect 46112 33584 46164 33590
rect 46112 33526 46164 33532
rect 46124 31414 46152 33526
rect 46296 32904 46348 32910
rect 46296 32846 46348 32852
rect 46204 32360 46256 32366
rect 46204 32302 46256 32308
rect 46216 32065 46244 32302
rect 46202 32056 46258 32065
rect 46202 31991 46258 32000
rect 46308 31890 46336 32846
rect 46480 32224 46532 32230
rect 46480 32166 46532 32172
rect 46492 31890 46520 32166
rect 46296 31884 46348 31890
rect 46296 31826 46348 31832
rect 46480 31884 46532 31890
rect 46480 31826 46532 31832
rect 46112 31408 46164 31414
rect 46112 31350 46164 31356
rect 46020 31272 46072 31278
rect 46020 31214 46072 31220
rect 45928 24336 45980 24342
rect 45928 24278 45980 24284
rect 45836 24132 45888 24138
rect 45836 24074 45888 24080
rect 45744 23180 45796 23186
rect 45744 23122 45796 23128
rect 45756 22710 45784 23122
rect 45744 22704 45796 22710
rect 45744 22646 45796 22652
rect 45652 20936 45704 20942
rect 45652 20878 45704 20884
rect 45560 20528 45612 20534
rect 45560 20470 45612 20476
rect 44640 20460 44692 20466
rect 44640 20402 44692 20408
rect 45192 20392 45244 20398
rect 45192 20334 45244 20340
rect 45204 20058 45232 20334
rect 45192 20052 45244 20058
rect 45192 19994 45244 20000
rect 44824 19848 44876 19854
rect 44824 19790 44876 19796
rect 44836 17490 44864 19790
rect 45560 19440 45612 19446
rect 45560 19382 45612 19388
rect 45468 19168 45520 19174
rect 45468 19110 45520 19116
rect 45480 18834 45508 19110
rect 45468 18828 45520 18834
rect 45468 18770 45520 18776
rect 44916 18760 44968 18766
rect 44916 18702 44968 18708
rect 45100 18760 45152 18766
rect 45100 18702 45152 18708
rect 44928 17678 44956 18702
rect 45008 18216 45060 18222
rect 45008 18158 45060 18164
rect 44916 17672 44968 17678
rect 44916 17614 44968 17620
rect 44836 17462 44956 17490
rect 44928 16658 44956 17462
rect 44916 16652 44968 16658
rect 44916 16594 44968 16600
rect 44548 13932 44600 13938
rect 44548 13874 44600 13880
rect 44928 6914 44956 16594
rect 45020 15570 45048 18158
rect 45112 17610 45140 18702
rect 45572 17814 45600 19382
rect 45560 17808 45612 17814
rect 45560 17750 45612 17756
rect 45100 17604 45152 17610
rect 45100 17546 45152 17552
rect 45008 15564 45060 15570
rect 45008 15506 45060 15512
rect 45112 8022 45140 17546
rect 45192 16448 45244 16454
rect 45192 16390 45244 16396
rect 45204 15570 45232 16390
rect 45468 16040 45520 16046
rect 45468 15982 45520 15988
rect 45192 15564 45244 15570
rect 45192 15506 45244 15512
rect 45284 8492 45336 8498
rect 45284 8434 45336 8440
rect 45296 8378 45324 8434
rect 45296 8350 45416 8378
rect 45100 8016 45152 8022
rect 45100 7958 45152 7964
rect 45112 7546 45140 7958
rect 45388 7818 45416 8350
rect 45284 7812 45336 7818
rect 45284 7754 45336 7760
rect 45376 7812 45428 7818
rect 45376 7754 45428 7760
rect 45100 7540 45152 7546
rect 45100 7482 45152 7488
rect 44928 6886 45048 6914
rect 43628 5160 43680 5166
rect 43628 5102 43680 5108
rect 43812 5160 43864 5166
rect 43812 5102 43864 5108
rect 42524 4820 42576 4826
rect 42524 4762 42576 4768
rect 42892 4616 42944 4622
rect 42892 4558 42944 4564
rect 42616 4548 42668 4554
rect 42616 4490 42668 4496
rect 42524 3664 42576 3670
rect 42524 3606 42576 3612
rect 42432 2576 42484 2582
rect 42432 2518 42484 2524
rect 41328 2304 41380 2310
rect 41328 2246 41380 2252
rect 41340 2038 41368 2246
rect 41328 2032 41380 2038
rect 41328 1974 41380 1980
rect 42536 800 42564 3606
rect 42628 3466 42656 4490
rect 42800 4208 42852 4214
rect 42800 4150 42852 4156
rect 42616 3460 42668 3466
rect 42616 3402 42668 3408
rect 42628 3126 42656 3402
rect 42616 3120 42668 3126
rect 42616 3062 42668 3068
rect 42812 2446 42840 4150
rect 42904 2650 42932 4558
rect 43824 4214 43852 5102
rect 45020 4622 45048 6886
rect 45008 4616 45060 4622
rect 45008 4558 45060 4564
rect 43812 4208 43864 4214
rect 43812 4150 43864 4156
rect 45296 4078 45324 7754
rect 45388 4690 45416 7754
rect 45376 4684 45428 4690
rect 45376 4626 45428 4632
rect 45284 4072 45336 4078
rect 45284 4014 45336 4020
rect 45480 3618 45508 15982
rect 45112 3590 45508 3618
rect 43904 3528 43956 3534
rect 43904 3470 43956 3476
rect 43076 3392 43128 3398
rect 43076 3334 43128 3340
rect 43088 3126 43116 3334
rect 43076 3120 43128 3126
rect 43076 3062 43128 3068
rect 43916 2990 43944 3470
rect 43904 2984 43956 2990
rect 43904 2926 43956 2932
rect 43168 2916 43220 2922
rect 43168 2858 43220 2864
rect 42892 2644 42944 2650
rect 42892 2586 42944 2592
rect 42800 2440 42852 2446
rect 42800 2382 42852 2388
rect 43180 800 43208 2858
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 45112 800 45140 3590
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 45204 3058 45232 3470
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45388 3126 45416 3334
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 45664 2854 45692 20878
rect 45848 19854 45876 24074
rect 46032 22658 46060 31214
rect 45940 22630 46060 22658
rect 45940 20806 45968 22630
rect 46018 22536 46074 22545
rect 46018 22471 46074 22480
rect 46032 22030 46060 22471
rect 46020 22024 46072 22030
rect 46020 21966 46072 21972
rect 45928 20800 45980 20806
rect 45928 20742 45980 20748
rect 46020 20392 46072 20398
rect 46020 20334 46072 20340
rect 45836 19848 45888 19854
rect 45836 19790 45888 19796
rect 45928 19712 45980 19718
rect 45928 19654 45980 19660
rect 45940 19378 45968 19654
rect 45928 19372 45980 19378
rect 45928 19314 45980 19320
rect 45836 18760 45888 18766
rect 45836 18702 45888 18708
rect 45848 18465 45876 18702
rect 45834 18456 45890 18465
rect 45834 18391 45890 18400
rect 45744 8288 45796 8294
rect 45744 8230 45796 8236
rect 45756 7478 45784 8230
rect 45744 7472 45796 7478
rect 45744 7414 45796 7420
rect 46032 3641 46060 20334
rect 46124 9450 46152 31350
rect 46386 30016 46442 30025
rect 46386 29951 46442 29960
rect 46400 28014 46428 29951
rect 46388 28008 46440 28014
rect 46388 27950 46440 27956
rect 46296 26784 46348 26790
rect 46296 26726 46348 26732
rect 46308 26450 46336 26726
rect 46296 26444 46348 26450
rect 46296 26386 46348 26392
rect 46388 26240 46440 26246
rect 46388 26182 46440 26188
rect 46400 25838 46428 26182
rect 46388 25832 46440 25838
rect 46388 25774 46440 25780
rect 46296 25764 46348 25770
rect 46296 25706 46348 25712
rect 46204 24200 46256 24206
rect 46204 24142 46256 24148
rect 46216 23798 46244 24142
rect 46204 23792 46256 23798
rect 46204 23734 46256 23740
rect 46308 23186 46336 25706
rect 46480 25696 46532 25702
rect 46480 25638 46532 25644
rect 46492 25362 46520 25638
rect 46480 25356 46532 25362
rect 46480 25298 46532 25304
rect 46480 25220 46532 25226
rect 46480 25162 46532 25168
rect 46388 24608 46440 24614
rect 46388 24550 46440 24556
rect 46400 24274 46428 24550
rect 46388 24268 46440 24274
rect 46388 24210 46440 24216
rect 46296 23180 46348 23186
rect 46296 23122 46348 23128
rect 46204 22024 46256 22030
rect 46204 21966 46256 21972
rect 46216 21078 46244 21966
rect 46388 21888 46440 21894
rect 46388 21830 46440 21836
rect 46204 21072 46256 21078
rect 46204 21014 46256 21020
rect 46400 19922 46428 21830
rect 46492 20602 46520 25162
rect 46584 24614 46612 44134
rect 46768 43246 46796 45970
rect 46860 45558 46888 47382
rect 47044 46646 47072 49200
rect 47688 47054 47716 49200
rect 48134 47696 48190 47705
rect 48134 47631 48190 47640
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47032 46640 47084 46646
rect 47032 46582 47084 46588
rect 47952 46572 48004 46578
rect 47952 46514 48004 46520
rect 47860 46368 47912 46374
rect 47964 46345 47992 46514
rect 47860 46310 47912 46316
rect 47950 46336 48006 46345
rect 46940 45892 46992 45898
rect 46940 45834 46992 45840
rect 46848 45552 46900 45558
rect 46848 45494 46900 45500
rect 46952 44538 46980 45834
rect 47492 45484 47544 45490
rect 47492 45426 47544 45432
rect 46940 44532 46992 44538
rect 46940 44474 46992 44480
rect 47504 44402 47532 45426
rect 46848 44396 46900 44402
rect 46848 44338 46900 44344
rect 47492 44396 47544 44402
rect 47492 44338 47544 44344
rect 46756 43240 46808 43246
rect 46756 43182 46808 43188
rect 46860 41138 46888 44338
rect 47308 44328 47360 44334
rect 47308 44270 47360 44276
rect 47320 42226 47348 44270
rect 47308 42220 47360 42226
rect 47308 42162 47360 42168
rect 46940 41540 46992 41546
rect 46940 41482 46992 41488
rect 46952 41274 46980 41482
rect 46940 41268 46992 41274
rect 46940 41210 46992 41216
rect 46848 41132 46900 41138
rect 46848 41074 46900 41080
rect 46756 38956 46808 38962
rect 46756 38898 46808 38904
rect 46768 26246 46796 38898
rect 46860 38826 46888 41074
rect 46940 39364 46992 39370
rect 46940 39306 46992 39312
rect 46952 39098 46980 39306
rect 46940 39092 46992 39098
rect 46940 39034 46992 39040
rect 46848 38820 46900 38826
rect 46848 38762 46900 38768
rect 47124 34944 47176 34950
rect 47124 34886 47176 34892
rect 47032 33040 47084 33046
rect 47032 32982 47084 32988
rect 47044 31278 47072 32982
rect 47136 32978 47164 34886
rect 47216 33312 47268 33318
rect 47216 33254 47268 33260
rect 47124 32972 47176 32978
rect 47124 32914 47176 32920
rect 47228 32842 47256 33254
rect 47216 32836 47268 32842
rect 47216 32778 47268 32784
rect 47032 31272 47084 31278
rect 47032 31214 47084 31220
rect 46846 28656 46902 28665
rect 46846 28591 46902 28600
rect 46860 26466 46888 28591
rect 46940 28552 46992 28558
rect 46940 28494 46992 28500
rect 46952 27606 46980 28494
rect 46940 27600 46992 27606
rect 46940 27542 46992 27548
rect 46860 26438 46980 26466
rect 46848 26308 46900 26314
rect 46848 26250 46900 26256
rect 46756 26240 46808 26246
rect 46860 26217 46888 26250
rect 46756 26182 46808 26188
rect 46846 26208 46902 26217
rect 46846 26143 46902 26152
rect 46952 26058 46980 26438
rect 46768 26030 46980 26058
rect 46664 25900 46716 25906
rect 46664 25842 46716 25848
rect 46572 24608 46624 24614
rect 46572 24550 46624 24556
rect 46480 20596 46532 20602
rect 46480 20538 46532 20544
rect 46492 19990 46520 20538
rect 46480 19984 46532 19990
rect 46480 19926 46532 19932
rect 46388 19916 46440 19922
rect 46388 19858 46440 19864
rect 46204 19168 46256 19174
rect 46204 19110 46256 19116
rect 46216 18358 46244 19110
rect 46204 18352 46256 18358
rect 46204 18294 46256 18300
rect 46296 17672 46348 17678
rect 46296 17614 46348 17620
rect 46308 17202 46336 17614
rect 46296 17196 46348 17202
rect 46296 17138 46348 17144
rect 46296 16516 46348 16522
rect 46296 16458 46348 16464
rect 46308 15745 46336 16458
rect 46294 15736 46350 15745
rect 46294 15671 46350 15680
rect 46480 13728 46532 13734
rect 46480 13670 46532 13676
rect 46492 13394 46520 13670
rect 46480 13388 46532 13394
rect 46480 13330 46532 13336
rect 46296 13320 46348 13326
rect 46296 13262 46348 13268
rect 46308 12850 46336 13262
rect 46296 12844 46348 12850
rect 46296 12786 46348 12792
rect 46296 11552 46348 11558
rect 46296 11494 46348 11500
rect 46308 11218 46336 11494
rect 46296 11212 46348 11218
rect 46296 11154 46348 11160
rect 46480 11076 46532 11082
rect 46480 11018 46532 11024
rect 46492 10810 46520 11018
rect 46480 10804 46532 10810
rect 46480 10746 46532 10752
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46480 10464 46532 10470
rect 46480 10406 46532 10412
rect 46308 10130 46336 10406
rect 46492 10130 46520 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 46480 10124 46532 10130
rect 46480 10066 46532 10072
rect 46112 9444 46164 9450
rect 46112 9386 46164 9392
rect 46480 4480 46532 4486
rect 46480 4422 46532 4428
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46018 3632 46074 3641
rect 46308 3602 46336 3878
rect 46492 3602 46520 4422
rect 46584 3670 46612 24550
rect 46676 23225 46704 25842
rect 46662 23216 46718 23225
rect 46662 23151 46718 23160
rect 46768 21146 46796 26030
rect 46846 25800 46902 25809
rect 46846 25735 46902 25744
rect 46860 24818 46888 25735
rect 46848 24812 46900 24818
rect 46848 24754 46900 24760
rect 46848 24676 46900 24682
rect 46848 24618 46900 24624
rect 46860 23905 46888 24618
rect 46846 23896 46902 23905
rect 46846 23831 46902 23840
rect 46940 23044 46992 23050
rect 46940 22986 46992 22992
rect 46952 22778 46980 22986
rect 46940 22772 46992 22778
rect 46940 22714 46992 22720
rect 47044 21622 47072 31214
rect 47216 29708 47268 29714
rect 47216 29650 47268 29656
rect 47124 24812 47176 24818
rect 47124 24754 47176 24760
rect 47032 21616 47084 21622
rect 47032 21558 47084 21564
rect 46848 21480 46900 21486
rect 46848 21422 46900 21428
rect 46756 21140 46808 21146
rect 46756 21082 46808 21088
rect 46860 19922 46888 21422
rect 46848 19916 46900 19922
rect 46848 19858 46900 19864
rect 46860 18222 46888 19858
rect 47032 18284 47084 18290
rect 47032 18226 47084 18232
rect 46848 18216 46900 18222
rect 46848 18158 46900 18164
rect 46860 17218 46888 18158
rect 47044 17898 47072 18226
rect 47136 18170 47164 24754
rect 47228 22574 47256 29650
rect 47320 22710 47348 42162
rect 47504 32434 47532 44338
rect 47676 44192 47728 44198
rect 47676 44134 47728 44140
rect 47688 43858 47716 44134
rect 47676 43852 47728 43858
rect 47676 43794 47728 43800
rect 47676 42628 47728 42634
rect 47676 42570 47728 42576
rect 47688 42362 47716 42570
rect 47676 42356 47728 42362
rect 47676 42298 47728 42304
rect 47676 41676 47728 41682
rect 47676 41618 47728 41624
rect 47688 40730 47716 41618
rect 47676 40724 47728 40730
rect 47676 40666 47728 40672
rect 47676 38956 47728 38962
rect 47676 38898 47728 38904
rect 47688 38865 47716 38898
rect 47674 38856 47730 38865
rect 47674 38791 47730 38800
rect 47676 38276 47728 38282
rect 47676 38218 47728 38224
rect 47688 38010 47716 38218
rect 47676 38004 47728 38010
rect 47676 37946 47728 37952
rect 47584 37868 47636 37874
rect 47584 37810 47636 37816
rect 47492 32428 47544 32434
rect 47492 32370 47544 32376
rect 47400 29640 47452 29646
rect 47400 29582 47452 29588
rect 47412 29345 47440 29582
rect 47398 29336 47454 29345
rect 47398 29271 47454 29280
rect 47504 23866 47532 32370
rect 47596 28082 47624 37810
rect 47872 35894 47900 46310
rect 47950 46271 48006 46280
rect 48148 46034 48176 47631
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 48136 46028 48188 46034
rect 48136 45970 48188 45976
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 48240 43858 48268 44911
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 48136 41608 48188 41614
rect 48134 41576 48136 41585
rect 48188 41576 48190 41585
rect 48134 41511 48190 41520
rect 47952 41132 48004 41138
rect 47952 41074 48004 41080
rect 47964 40905 47992 41074
rect 48044 40928 48096 40934
rect 47950 40896 48006 40905
rect 48044 40870 48096 40876
rect 47950 40831 48006 40840
rect 47780 35866 47900 35894
rect 47584 28076 47636 28082
rect 47584 28018 47636 28024
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 47688 27538 47716 27814
rect 47676 27532 47728 27538
rect 47676 27474 47728 27480
rect 47780 26234 47808 35866
rect 47860 34400 47912 34406
rect 47860 34342 47912 34348
rect 47872 33318 47900 34342
rect 47952 33992 48004 33998
rect 47952 33934 48004 33940
rect 48056 33946 48084 40870
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48148 39506 48176 40151
rect 48136 39500 48188 39506
rect 48136 39442 48188 39448
rect 48136 38276 48188 38282
rect 48136 38218 48188 38224
rect 48148 38185 48176 38218
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48136 35080 48188 35086
rect 48136 35022 48188 35028
rect 48148 34785 48176 35022
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48136 34604 48188 34610
rect 48136 34546 48188 34552
rect 48148 34105 48176 34546
rect 48134 34096 48190 34105
rect 48134 34031 48190 34040
rect 47964 33425 47992 33934
rect 48056 33918 48176 33946
rect 48044 33856 48096 33862
rect 48044 33798 48096 33804
rect 48056 33658 48084 33798
rect 48044 33652 48096 33658
rect 48044 33594 48096 33600
rect 47950 33416 48006 33425
rect 47950 33351 48006 33360
rect 47860 33312 47912 33318
rect 47860 33254 47912 33260
rect 48148 32858 48176 33918
rect 47688 26206 47808 26234
rect 48056 32830 48176 32858
rect 47492 23860 47544 23866
rect 47492 23802 47544 23808
rect 47584 23724 47636 23730
rect 47584 23666 47636 23672
rect 47308 22704 47360 22710
rect 47308 22646 47360 22652
rect 47216 22568 47268 22574
rect 47216 22510 47268 22516
rect 47228 21554 47256 22510
rect 47320 22114 47348 22646
rect 47596 22438 47624 23666
rect 47584 22432 47636 22438
rect 47584 22374 47636 22380
rect 47320 22086 47440 22114
rect 47308 22024 47360 22030
rect 47308 21966 47360 21972
rect 47320 21865 47348 21966
rect 47306 21856 47362 21865
rect 47306 21791 47362 21800
rect 47216 21548 47268 21554
rect 47216 21490 47268 21496
rect 47228 20262 47256 21490
rect 47216 20256 47268 20262
rect 47216 20198 47268 20204
rect 47412 18290 47440 22086
rect 47492 21616 47544 21622
rect 47492 21558 47544 21564
rect 47400 18284 47452 18290
rect 47400 18226 47452 18232
rect 47136 18142 47440 18170
rect 47044 17870 47348 17898
rect 46768 17190 46888 17218
rect 46768 17134 46796 17190
rect 46756 17128 46808 17134
rect 46756 17070 46808 17076
rect 46940 16992 46992 16998
rect 46940 16934 46992 16940
rect 46952 16522 46980 16934
rect 46940 16516 46992 16522
rect 46940 16458 46992 16464
rect 47320 15638 47348 17870
rect 47308 15632 47360 15638
rect 47308 15574 47360 15580
rect 46664 15564 46716 15570
rect 46664 15506 46716 15512
rect 46572 3664 46624 3670
rect 46572 3606 46624 3612
rect 46018 3567 46074 3576
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 46676 3505 46704 15506
rect 47412 10674 47440 18142
rect 47400 10668 47452 10674
rect 47400 10610 47452 10616
rect 46846 8256 46902 8265
rect 46846 8191 46902 8200
rect 46860 8090 46888 8191
rect 46848 8084 46900 8090
rect 46848 8026 46900 8032
rect 47504 7954 47532 21558
rect 47688 19718 47716 26206
rect 47768 26036 47820 26042
rect 47768 25978 47820 25984
rect 47780 23798 47808 25978
rect 47768 23792 47820 23798
rect 47768 23734 47820 23740
rect 47780 22642 47808 23734
rect 48056 23594 48084 32830
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48148 31890 48176 32671
rect 48136 31884 48188 31890
rect 48136 31826 48188 31832
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48228 26308 48280 26314
rect 48228 26250 48280 26256
rect 48134 25936 48190 25945
rect 48134 25871 48190 25880
rect 48148 25362 48176 25871
rect 48136 25356 48188 25362
rect 48136 25298 48188 25304
rect 48240 25265 48268 26250
rect 48226 25256 48282 25265
rect 48226 25191 48282 25200
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48044 23588 48096 23594
rect 48044 23530 48096 23536
rect 48148 23186 48176 24511
rect 48136 23180 48188 23186
rect 48136 23122 48188 23128
rect 48136 22976 48188 22982
rect 48136 22918 48188 22924
rect 48148 22778 48176 22918
rect 48136 22772 48188 22778
rect 48136 22714 48188 22720
rect 47768 22636 47820 22642
rect 47768 22578 47820 22584
rect 47780 21690 47808 22578
rect 47860 22568 47912 22574
rect 47860 22510 47912 22516
rect 47768 21684 47820 21690
rect 47768 21626 47820 21632
rect 47872 21622 47900 22510
rect 47952 22500 48004 22506
rect 47952 22442 48004 22448
rect 47964 21690 47992 22442
rect 48044 21956 48096 21962
rect 48044 21898 48096 21904
rect 47952 21684 48004 21690
rect 47952 21626 48004 21632
rect 47860 21616 47912 21622
rect 47860 21558 47912 21564
rect 47964 20466 47992 21626
rect 48056 20602 48084 21898
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48044 20596 48096 20602
rect 48044 20538 48096 20544
rect 47952 20460 48004 20466
rect 47952 20402 48004 20408
rect 47676 19712 47728 19718
rect 47676 19654 47728 19660
rect 47964 19666 47992 20402
rect 47688 19378 47716 19654
rect 47964 19638 48084 19666
rect 48056 19514 48084 19638
rect 47952 19508 48004 19514
rect 47952 19450 48004 19456
rect 48044 19508 48096 19514
rect 48044 19450 48096 19456
rect 47676 19372 47728 19378
rect 47676 19314 47728 19320
rect 47860 19236 47912 19242
rect 47860 19178 47912 19184
rect 47676 18692 47728 18698
rect 47676 18634 47728 18640
rect 47688 18426 47716 18634
rect 47676 18420 47728 18426
rect 47676 18362 47728 18368
rect 47676 17604 47728 17610
rect 47676 17546 47728 17552
rect 47688 17338 47716 17546
rect 47872 17542 47900 19178
rect 47964 17746 47992 19450
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48148 18834 48176 19071
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 47952 17740 48004 17746
rect 47952 17682 48004 17688
rect 47860 17536 47912 17542
rect 47860 17478 47912 17484
rect 47676 17332 47728 17338
rect 47676 17274 47728 17280
rect 47584 17060 47636 17066
rect 47584 17002 47636 17008
rect 47492 7948 47544 7954
rect 47492 7890 47544 7896
rect 47308 7880 47360 7886
rect 47308 7822 47360 7828
rect 47320 7585 47348 7822
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47596 6914 47624 17002
rect 47768 16652 47820 16658
rect 47768 16594 47820 16600
rect 47780 16114 47808 16594
rect 47768 16108 47820 16114
rect 47768 16050 47820 16056
rect 47872 11778 47900 17478
rect 47504 6886 47624 6914
rect 47688 11750 47900 11778
rect 46848 4616 46900 4622
rect 46848 4558 46900 4564
rect 46860 4185 46888 4558
rect 46846 4176 46902 4185
rect 46756 4140 46808 4146
rect 46846 4111 46902 4120
rect 46756 4082 46808 4088
rect 46662 3496 46718 3505
rect 46662 3431 46718 3440
rect 45652 2848 45704 2854
rect 45652 2790 45704 2796
rect 46388 2372 46440 2378
rect 46388 2314 46440 2320
rect 46400 800 46428 2314
rect 2962 776 3018 785
rect 2962 711 3018 720
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46768 105 46796 4082
rect 47504 3466 47532 6886
rect 47492 3460 47544 3466
rect 47492 3402 47544 3408
rect 47688 3194 47716 11750
rect 47858 9616 47914 9625
rect 47858 9551 47860 9560
rect 47912 9551 47914 9560
rect 47860 9522 47912 9528
rect 47766 8936 47822 8945
rect 47766 8871 47768 8880
rect 47820 8871 47822 8880
rect 47768 8842 47820 8848
rect 47964 6914 47992 17682
rect 48136 17604 48188 17610
rect 48136 17546 48188 17552
rect 48148 17105 48176 17546
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48136 16516 48188 16522
rect 48136 16458 48188 16464
rect 48148 16425 48176 16458
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48136 13252 48188 13258
rect 48136 13194 48188 13200
rect 48148 12345 48176 13194
rect 48134 12336 48190 12345
rect 48134 12271 48190 12280
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 48228 7404 48280 7410
rect 48228 7346 48280 7352
rect 47872 6886 47992 6914
rect 48240 6905 48268 7346
rect 48226 6896 48282 6905
rect 47768 4208 47820 4214
rect 47768 4150 47820 4156
rect 47676 3188 47728 3194
rect 47676 3130 47728 3136
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 47044 800 47072 2382
rect 47688 800 47716 2926
rect 47780 1465 47808 4150
rect 47872 2514 47900 6886
rect 48226 6831 48282 6840
rect 47952 6316 48004 6322
rect 47952 6258 48004 6264
rect 47964 6225 47992 6258
rect 47950 6216 48006 6225
rect 47950 6151 48006 6160
rect 47952 5228 48004 5234
rect 47952 5170 48004 5176
rect 47964 3505 47992 5170
rect 47950 3496 48006 3505
rect 47950 3431 48006 3440
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48320 3052 48372 3058
rect 48320 2994 48372 3000
rect 47860 2508 47912 2514
rect 47860 2450 47912 2456
rect 48044 2440 48096 2446
rect 48044 2382 48096 2388
rect 47766 1456 47822 1465
rect 47766 1391 47822 1400
rect 46754 96 46810 105
rect 46754 31 46810 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48056 785 48084 2382
rect 48332 800 48360 2994
rect 48976 800 49004 3402
rect 48042 776 48098 785
rect 48042 711 48098 720
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1858 47640 1914 47696
rect 3422 46960 3478 47016
rect 1398 42880 1454 42936
rect 1398 40160 1454 40216
rect 1398 33360 1454 33416
rect 1858 41520 1914 41576
rect 1582 35400 1638 35456
rect 1582 32680 1638 32736
rect 1582 23588 1638 23624
rect 1582 23568 1584 23588
rect 1584 23568 1636 23588
rect 1636 23568 1638 23588
rect 1398 23160 1454 23216
rect 1858 25236 1860 25256
rect 1860 25236 1912 25256
rect 1912 25236 1914 25256
rect 1858 25200 1914 25236
rect 1398 17720 1454 17776
rect 1398 12280 1454 12336
rect 2778 46280 2834 46336
rect 2962 36760 3018 36816
rect 2778 32000 2834 32056
rect 3330 44920 3386 44976
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3606 43560 3662 43616
rect 3514 39480 3570 39536
rect 3882 31320 3938 31376
rect 3974 28600 4030 28656
rect 3054 19760 3110 19816
rect 2778 19080 2834 19136
rect 3330 18400 3386 18456
rect 3514 17040 3570 17096
rect 2778 16360 2834 16416
rect 2778 15000 2834 15056
rect 3146 10240 3202 10296
rect 3422 13640 3478 13696
rect 3330 7520 3386 7576
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3422 6860 3478 6896
rect 3422 6840 3424 6860
rect 3424 6840 3476 6860
rect 3476 6840 3478 6860
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3882 3576 3938 3632
rect 3422 3440 3478 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4066 1400 4122 1456
rect 16026 21548 16082 21584
rect 16026 21528 16028 21548
rect 16028 21528 16080 21548
rect 16080 21528 16082 21548
rect 17590 3440 17646 3496
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 28722 46980 28778 47016
rect 28722 46960 28724 46980
rect 28724 46960 28776 46980
rect 28776 46960 28778 46980
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 20626 26832 20682 26888
rect 21270 24828 21272 24848
rect 21272 24828 21324 24848
rect 21324 24828 21326 24848
rect 21270 24792 21326 24828
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 21730 28600 21786 28656
rect 21822 24132 21878 24168
rect 21822 24112 21824 24132
rect 21824 24112 21876 24132
rect 21876 24112 21878 24132
rect 25042 27376 25098 27432
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 24766 19352 24822 19408
rect 25594 19372 25650 19408
rect 25594 19352 25596 19372
rect 25596 19352 25648 19372
rect 25648 19352 25650 19372
rect 26974 27648 27030 27704
rect 27342 28600 27398 28656
rect 27710 28636 27712 28656
rect 27712 28636 27764 28656
rect 27764 28636 27766 28656
rect 27710 28600 27766 28636
rect 28170 26832 28226 26888
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 28906 32272 28962 32328
rect 28906 31864 28962 31920
rect 28538 27668 28594 27704
rect 28538 27648 28540 27668
rect 28540 27648 28592 27668
rect 28592 27648 28594 27668
rect 28722 27396 28778 27432
rect 28722 27376 28724 27396
rect 28724 27376 28776 27396
rect 28776 27376 28778 27396
rect 29366 25220 29422 25256
rect 29366 25200 29368 25220
rect 29368 25200 29420 25220
rect 29420 25200 29422 25220
rect 29642 25472 29698 25528
rect 29642 23724 29698 23760
rect 29642 23704 29644 23724
rect 29644 23704 29696 23724
rect 29696 23704 29698 23724
rect 28998 20984 29054 21040
rect 30102 23724 30158 23760
rect 30102 23704 30104 23724
rect 30104 23704 30156 23724
rect 30156 23704 30158 23724
rect 31574 31864 31630 31920
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 31850 31864 31906 31920
rect 32494 31864 32550 31920
rect 31850 25200 31906 25256
rect 31206 21004 31262 21040
rect 31206 20984 31208 21004
rect 31208 20984 31260 21004
rect 31260 20984 31262 21004
rect 31666 19760 31722 19816
rect 32126 21004 32182 21040
rect 32126 20984 32128 21004
rect 32128 20984 32180 21004
rect 32180 20984 32182 21004
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 33138 23568 33194 23624
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34242 25492 34298 25528
rect 34242 25472 34244 25492
rect 34244 25472 34296 25492
rect 34296 25472 34298 25492
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34518 21936 34574 21992
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 37278 24112 37334 24168
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 40038 24792 40094 24848
rect 45926 39480 45982 39536
rect 45282 26288 45338 26344
rect 46202 32000 46258 32056
rect 46018 22480 46074 22536
rect 45834 18400 45890 18456
rect 46386 29960 46442 30016
rect 48134 47640 48190 47696
rect 46846 28600 46902 28656
rect 46846 26152 46902 26208
rect 46294 15680 46350 15736
rect 46018 3576 46074 3632
rect 46662 23160 46718 23216
rect 46846 25744 46902 25800
rect 46846 23840 46902 23896
rect 47674 38800 47730 38856
rect 47398 29280 47454 29336
rect 47950 46280 48006 46336
rect 48134 45600 48190 45656
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 48134 41556 48136 41576
rect 48136 41556 48188 41576
rect 48188 41556 48190 41576
rect 48134 41520 48190 41556
rect 47950 40840 48006 40896
rect 48134 40160 48190 40216
rect 48134 38120 48190 38176
rect 48134 34720 48190 34776
rect 48134 34040 48190 34096
rect 47950 33360 48006 33416
rect 47306 21800 47362 21856
rect 46846 8200 46902 8256
rect 48134 32680 48190 32736
rect 48134 27920 48190 27976
rect 48134 25880 48190 25936
rect 48226 25200 48282 25256
rect 48134 24520 48190 24576
rect 48134 21120 48190 21176
rect 48134 19080 48190 19136
rect 47306 7520 47362 7576
rect 46846 4120 46902 4176
rect 46662 3440 46718 3496
rect 2962 720 3018 776
rect 47858 9580 47914 9616
rect 47858 9560 47860 9580
rect 47860 9560 47912 9580
rect 47912 9560 47914 9580
rect 47766 8900 47822 8936
rect 47766 8880 47768 8900
rect 47768 8880 47820 8900
rect 47820 8880 47822 8900
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 12280 48190 12336
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 48226 6840 48282 6896
rect 47950 6160 48006 6216
rect 47950 3440 48006 3496
rect 47766 1400 47822 1456
rect 46754 40 46810 96
rect 48042 720 48098 776
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1853 47698 1919 47701
rect 0 47696 1919 47698
rect 0 47640 1858 47696
rect 1914 47640 1919 47696
rect 0 47638 1919 47640
rect 0 47548 800 47638
rect 1853 47635 1919 47638
rect 48129 47698 48195 47701
rect 49200 47698 50000 47788
rect 48129 47696 50000 47698
rect 48129 47640 48134 47696
rect 48190 47640 50000 47696
rect 48129 47638 50000 47640
rect 48129 47635 48195 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3417 47018 3483 47021
rect 0 47016 3483 47018
rect 0 46960 3422 47016
rect 3478 46960 3483 47016
rect 0 46958 3483 46960
rect 0 46868 800 46958
rect 3417 46955 3483 46958
rect 28717 47020 28783 47021
rect 28717 47016 28764 47020
rect 28828 47018 28834 47020
rect 28717 46960 28722 47016
rect 28717 46956 28764 46960
rect 28828 46958 28874 47018
rect 28828 46956 28834 46958
rect 46054 46956 46060 47020
rect 46124 47018 46130 47020
rect 49200 47018 50000 47108
rect 46124 46958 50000 47018
rect 46124 46956 46130 46958
rect 28717 46955 28783 46956
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46188 800 46278
rect 2773 46275 2839 46278
rect 47945 46338 48011 46341
rect 49200 46338 50000 46428
rect 47945 46336 50000 46338
rect 47945 46280 47950 46336
rect 48006 46280 50000 46336
rect 47945 46278 50000 46280
rect 47945 46275 48011 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3325 44978 3391 44981
rect 0 44976 3391 44978
rect 0 44920 3330 44976
rect 3386 44920 3391 44976
rect 0 44918 3391 44920
rect 0 44828 800 44918
rect 3325 44915 3391 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3601 43618 3667 43621
rect 0 43616 3667 43618
rect 0 43560 3606 43616
rect 3662 43560 3667 43616
rect 0 43558 3667 43560
rect 0 43468 800 43558
rect 3601 43555 3667 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42788 800 42878
rect 1393 42875 1459 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 47945 40898 48011 40901
rect 49200 40898 50000 40988
rect 47945 40896 50000 40898
rect 47945 40840 47950 40896
rect 48006 40840 50000 40896
rect 47945 40838 50000 40840
rect 47945 40835 48011 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1393 40218 1459 40221
rect 0 40216 1459 40218
rect 0 40160 1398 40216
rect 1454 40160 1459 40216
rect 0 40158 1459 40160
rect 0 40068 800 40158
rect 1393 40155 1459 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40308
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3509 39538 3575 39541
rect 0 39536 3575 39538
rect 0 39480 3514 39536
rect 3570 39480 3575 39536
rect 0 39478 3575 39480
rect 0 39388 800 39478
rect 3509 39475 3575 39478
rect 45921 39538 45987 39541
rect 49200 39538 50000 39628
rect 45921 39536 50000 39538
rect 45921 39480 45926 39536
rect 45982 39480 50000 39536
rect 45921 39478 50000 39480
rect 45921 39475 45987 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47669 38858 47735 38861
rect 49200 38858 50000 38948
rect 47669 38856 50000 38858
rect 47669 38800 47674 38856
rect 47730 38800 50000 38856
rect 47669 38798 50000 38800
rect 47669 38795 47735 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2957 36818 3023 36821
rect 0 36816 3023 36818
rect 0 36760 2962 36816
rect 3018 36760 3023 36816
rect 0 36758 3023 36760
rect 0 36668 800 36758
rect 2957 36755 3023 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35458 800 35548
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 48129 34098 48195 34101
rect 49200 34098 50000 34188
rect 48129 34096 50000 34098
rect 48129 34040 48134 34096
rect 48190 34040 50000 34096
rect 48129 34038 50000 34040
rect 48129 34035 48195 34038
rect 49200 33948 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 47945 33418 48011 33421
rect 49200 33418 50000 33508
rect 47945 33416 50000 33418
rect 47945 33360 47950 33416
rect 48006 33360 50000 33416
rect 47945 33358 50000 33360
rect 47945 33355 48011 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32828
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32588 800 32678
rect 1577 32675 1643 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 49200 32588 50000 32678
rect 28901 32330 28967 32333
rect 28901 32328 29010 32330
rect 28901 32272 28906 32328
rect 28962 32272 29010 32328
rect 28901 32267 29010 32272
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 2773 32058 2839 32061
rect 0 32056 2839 32058
rect 0 32000 2778 32056
rect 2834 32000 2839 32056
rect 0 31998 2839 32000
rect 0 31908 800 31998
rect 2773 31995 2839 31998
rect 28950 31925 29010 32267
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 46197 32058 46263 32061
rect 49200 32058 50000 32148
rect 46197 32056 50000 32058
rect 46197 32000 46202 32056
rect 46258 32000 50000 32056
rect 46197 31998 50000 32000
rect 46197 31995 46263 31998
rect 28901 31920 29010 31925
rect 28901 31864 28906 31920
rect 28962 31864 29010 31920
rect 28901 31862 29010 31864
rect 31569 31922 31635 31925
rect 31845 31922 31911 31925
rect 32489 31922 32555 31925
rect 31569 31920 32555 31922
rect 31569 31864 31574 31920
rect 31630 31864 31850 31920
rect 31906 31864 32494 31920
rect 32550 31864 32555 31920
rect 49200 31908 50000 31998
rect 31569 31862 32555 31864
rect 28901 31859 28967 31862
rect 31569 31859 31635 31862
rect 31845 31859 31911 31862
rect 32489 31859 32555 31862
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3877 31378 3943 31381
rect 0 31376 3943 31378
rect 0 31320 3882 31376
rect 3938 31320 3943 31376
rect 0 31318 3943 31320
rect 0 31228 800 31318
rect 3877 31315 3943 31318
rect 46238 31316 46244 31380
rect 46308 31378 46314 31380
rect 49200 31378 50000 31468
rect 46308 31318 50000 31378
rect 46308 31316 46314 31318
rect 49200 31228 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 29868 800 30108
rect 46381 30018 46447 30021
rect 49200 30018 50000 30108
rect 46381 30016 50000 30018
rect 46381 29960 46386 30016
rect 46442 29960 50000 30016
rect 46381 29958 50000 29960
rect 46381 29955 46447 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 47393 29338 47459 29341
rect 49200 29338 50000 29428
rect 47393 29336 50000 29338
rect 47393 29280 47398 29336
rect 47454 29280 50000 29336
rect 47393 29278 50000 29280
rect 47393 29275 47459 29278
rect 49200 29188 50000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3969 28658 4035 28661
rect 0 28656 4035 28658
rect 0 28600 3974 28656
rect 4030 28600 4035 28656
rect 0 28598 4035 28600
rect 0 28508 800 28598
rect 3969 28595 4035 28598
rect 21725 28658 21791 28661
rect 27337 28658 27403 28661
rect 27705 28658 27771 28661
rect 21725 28656 27771 28658
rect 21725 28600 21730 28656
rect 21786 28600 27342 28656
rect 27398 28600 27710 28656
rect 27766 28600 27771 28656
rect 21725 28598 27771 28600
rect 21725 28595 21791 28598
rect 27337 28595 27403 28598
rect 27705 28595 27771 28598
rect 46841 28658 46907 28661
rect 49200 28658 50000 28748
rect 46841 28656 50000 28658
rect 46841 28600 46846 28656
rect 46902 28600 50000 28656
rect 46841 28598 50000 28600
rect 46841 28595 46907 28598
rect 49200 28508 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 49200 27828 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 26969 27706 27035 27709
rect 28533 27706 28599 27709
rect 26969 27704 28599 27706
rect 26969 27648 26974 27704
rect 27030 27648 28538 27704
rect 28594 27648 28599 27704
rect 26969 27646 28599 27648
rect 26969 27643 27035 27646
rect 28533 27643 28599 27646
rect 25037 27434 25103 27437
rect 28717 27434 28783 27437
rect 25037 27432 28783 27434
rect 0 27148 800 27388
rect 25037 27376 25042 27432
rect 25098 27376 28722 27432
rect 28778 27376 28783 27432
rect 25037 27374 28783 27376
rect 25037 27371 25103 27374
rect 28717 27371 28783 27374
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 20621 26890 20687 26893
rect 28165 26890 28231 26893
rect 20621 26888 28231 26890
rect 20621 26832 20626 26888
rect 20682 26832 28170 26888
rect 28226 26832 28231 26888
rect 20621 26830 28231 26832
rect 20621 26827 20687 26830
rect 28165 26827 28231 26830
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 49200 26618 50000 26708
rect 45510 26558 50000 26618
rect 45277 26346 45343 26349
rect 45510 26346 45570 26558
rect 49200 26468 50000 26558
rect 45277 26344 45570 26346
rect 45277 26288 45282 26344
rect 45338 26288 45570 26344
rect 45277 26286 45570 26288
rect 45277 26283 45343 26286
rect 46841 26210 46907 26213
rect 46798 26208 46907 26210
rect 46798 26152 46846 26208
rect 46902 26152 46907 26208
rect 46798 26147 46907 26152
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 46798 25805 46858 26147
rect 48129 25938 48195 25941
rect 49200 25938 50000 26028
rect 48129 25936 50000 25938
rect 48129 25880 48134 25936
rect 48190 25880 50000 25936
rect 48129 25878 50000 25880
rect 48129 25875 48195 25878
rect 46798 25800 46907 25805
rect 46798 25744 46846 25800
rect 46902 25744 46907 25800
rect 49200 25788 50000 25878
rect 46798 25742 46907 25744
rect 46841 25739 46907 25742
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 29637 25530 29703 25533
rect 34237 25530 34303 25533
rect 29637 25528 34303 25530
rect 29637 25472 29642 25528
rect 29698 25472 34242 25528
rect 34298 25472 34303 25528
rect 29637 25470 34303 25472
rect 29637 25467 29703 25470
rect 34237 25467 34303 25470
rect 0 25258 800 25348
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25108 800 25198
rect 1853 25195 1919 25198
rect 29361 25258 29427 25261
rect 31845 25258 31911 25261
rect 29361 25256 31911 25258
rect 29361 25200 29366 25256
rect 29422 25200 31850 25256
rect 31906 25200 31911 25256
rect 29361 25198 31911 25200
rect 29361 25195 29427 25198
rect 31845 25195 31911 25198
rect 48221 25258 48287 25261
rect 49200 25258 50000 25348
rect 48221 25256 50000 25258
rect 48221 25200 48226 25256
rect 48282 25200 50000 25256
rect 48221 25198 50000 25200
rect 48221 25195 48287 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 21265 24850 21331 24853
rect 40033 24850 40099 24853
rect 21265 24848 40099 24850
rect 21265 24792 21270 24848
rect 21326 24792 40038 24848
rect 40094 24792 40099 24848
rect 21265 24790 40099 24792
rect 21265 24787 21331 24790
rect 40033 24787 40099 24790
rect 0 24428 800 24668
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 21817 24170 21883 24173
rect 37273 24170 37339 24173
rect 21817 24168 37339 24170
rect 21817 24112 21822 24168
rect 21878 24112 37278 24168
rect 37334 24112 37339 24168
rect 21817 24110 37339 24112
rect 21817 24107 21883 24110
rect 37273 24107 37339 24110
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 46841 23898 46907 23901
rect 49200 23898 50000 23988
rect 46841 23896 50000 23898
rect 46841 23840 46846 23896
rect 46902 23840 50000 23896
rect 46841 23838 50000 23840
rect 46841 23835 46907 23838
rect 29637 23762 29703 23765
rect 30097 23762 30163 23765
rect 29637 23760 30163 23762
rect 29637 23704 29642 23760
rect 29698 23704 30102 23760
rect 30158 23704 30163 23760
rect 49200 23748 50000 23838
rect 29637 23702 30163 23704
rect 29637 23699 29703 23702
rect 30097 23699 30163 23702
rect 1577 23626 1643 23629
rect 33133 23626 33199 23629
rect 1577 23624 33199 23626
rect 1577 23568 1582 23624
rect 1638 23568 33138 23624
rect 33194 23568 33199 23624
rect 1577 23566 33199 23568
rect 1577 23563 1643 23566
rect 33133 23563 33199 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23068 800 23158
rect 1393 23155 1459 23158
rect 46657 23218 46723 23221
rect 49200 23218 50000 23308
rect 46657 23216 50000 23218
rect 46657 23160 46662 23216
rect 46718 23160 50000 23216
rect 46657 23158 50000 23160
rect 46657 23155 46723 23158
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 46013 22538 46079 22541
rect 49200 22538 50000 22628
rect 46013 22536 50000 22538
rect 46013 22480 46018 22536
rect 46074 22480 50000 22536
rect 46013 22478 50000 22480
rect 46013 22475 46079 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21708 800 21948
rect 28758 21932 28764 21996
rect 28828 21994 28834 21996
rect 34513 21994 34579 21997
rect 28828 21992 34579 21994
rect 28828 21936 34518 21992
rect 34574 21936 34579 21992
rect 28828 21934 34579 21936
rect 28828 21932 28834 21934
rect 34513 21931 34579 21934
rect 47301 21858 47367 21861
rect 49200 21858 50000 21948
rect 47301 21856 50000 21858
rect 47301 21800 47306 21856
rect 47362 21800 50000 21856
rect 47301 21798 50000 21800
rect 47301 21795 47367 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 16021 21586 16087 21589
rect 46238 21586 46244 21588
rect 16021 21584 46244 21586
rect 16021 21528 16026 21584
rect 16082 21528 46244 21584
rect 16021 21526 46244 21528
rect 16021 21523 16087 21526
rect 46238 21524 46244 21526
rect 46308 21524 46314 21588
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 28993 21042 29059 21045
rect 31201 21042 31267 21045
rect 32121 21042 32187 21045
rect 28993 21040 32187 21042
rect 28993 20984 28998 21040
rect 29054 20984 31206 21040
rect 31262 20984 32126 21040
rect 32182 20984 32187 21040
rect 49200 21028 50000 21118
rect 28993 20982 32187 20984
rect 28993 20979 29059 20982
rect 31201 20979 31267 20982
rect 32121 20979 32187 20982
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 3049 19818 3115 19821
rect 0 19816 3115 19818
rect 0 19760 3054 19816
rect 3110 19760 3115 19816
rect 0 19758 3115 19760
rect 0 19668 800 19758
rect 3049 19755 3115 19758
rect 31661 19818 31727 19821
rect 46054 19818 46060 19820
rect 31661 19816 46060 19818
rect 31661 19760 31666 19816
rect 31722 19760 46060 19816
rect 31661 19758 46060 19760
rect 31661 19755 31727 19758
rect 46054 19756 46060 19758
rect 46124 19756 46130 19820
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 24761 19410 24827 19413
rect 25589 19410 25655 19413
rect 24761 19408 25655 19410
rect 24761 19352 24766 19408
rect 24822 19352 25594 19408
rect 25650 19352 25655 19408
rect 24761 19350 25655 19352
rect 24761 19347 24827 19350
rect 25589 19347 25655 19350
rect 0 19138 800 19228
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 18988 800 19078
rect 2773 19075 2839 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3325 18458 3391 18461
rect 0 18456 3391 18458
rect 0 18400 3330 18456
rect 3386 18400 3391 18456
rect 0 18398 3391 18400
rect 0 18308 800 18398
rect 3325 18395 3391 18398
rect 45829 18458 45895 18461
rect 49200 18458 50000 18548
rect 45829 18456 50000 18458
rect 45829 18400 45834 18456
rect 45890 18400 50000 18456
rect 45829 18398 50000 18400
rect 45829 18395 45895 18398
rect 49200 18308 50000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17628 800 17718
rect 1393 17715 1459 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3509 17098 3575 17101
rect 0 17096 3575 17098
rect 0 17040 3514 17096
rect 3570 17040 3575 17096
rect 0 17038 3575 17040
rect 0 16948 800 17038
rect 3509 17035 3575 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 2773 16418 2839 16421
rect 0 16416 2839 16418
rect 0 16360 2778 16416
rect 2834 16360 2839 16416
rect 0 16358 2839 16360
rect 0 16268 800 16358
rect 2773 16355 2839 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16508
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 46289 15738 46355 15741
rect 49200 15738 50000 15828
rect 46289 15736 50000 15738
rect 46289 15680 46294 15736
rect 46350 15680 50000 15736
rect 46289 15678 50000 15680
rect 46289 15675 46355 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3417 13698 3483 13701
rect 0 13696 3483 13698
rect 0 13640 3422 13696
rect 3478 13640 3483 13696
rect 0 13638 3483 13640
rect 0 13548 800 13638
rect 3417 13635 3483 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 3141 10298 3207 10301
rect 0 10296 3207 10298
rect 0 10240 3146 10296
rect 3202 10240 3207 10296
rect 0 10238 3207 10240
rect 0 10148 800 10238
rect 3141 10235 3207 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 47853 9618 47919 9621
rect 49200 9618 50000 9708
rect 47853 9616 50000 9618
rect 47853 9560 47858 9616
rect 47914 9560 50000 9616
rect 47853 9558 50000 9560
rect 47853 9555 47919 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47761 8938 47827 8941
rect 49200 8938 50000 9028
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 46841 8258 46907 8261
rect 49200 8258 50000 8348
rect 46841 8256 50000 8258
rect 46841 8200 46846 8256
rect 46902 8200 50000 8256
rect 46841 8198 50000 8200
rect 46841 8195 46907 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3325 7578 3391 7581
rect 0 7576 3391 7578
rect 0 7520 3330 7576
rect 3386 7520 3391 7576
rect 0 7518 3391 7520
rect 0 7428 800 7518
rect 3325 7515 3391 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 3417 6898 3483 6901
rect 0 6896 3483 6898
rect 0 6840 3422 6896
rect 3478 6840 3483 6896
rect 0 6838 3483 6840
rect 0 6748 800 6838
rect 3417 6835 3483 6838
rect 48221 6898 48287 6901
rect 49200 6898 50000 6988
rect 48221 6896 50000 6898
rect 48221 6840 48226 6896
rect 48282 6840 50000 6896
rect 48221 6838 50000 6840
rect 48221 6835 48287 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 47945 6218 48011 6221
rect 49200 6218 50000 6308
rect 47945 6216 50000 6218
rect 47945 6160 47950 6216
rect 48006 6160 50000 6216
rect 47945 6158 50000 6160
rect 47945 6155 48011 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 46841 4178 46907 4181
rect 49200 4178 50000 4268
rect 46841 4176 50000 4178
rect 46841 4120 46846 4176
rect 46902 4120 50000 4176
rect 46841 4118 50000 4120
rect 46841 4115 46907 4118
rect 49200 4028 50000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 3877 3634 3943 3637
rect 46013 3634 46079 3637
rect 3877 3632 46079 3634
rect 0 3498 800 3588
rect 3877 3576 3882 3632
rect 3938 3576 46018 3632
rect 46074 3576 46079 3632
rect 3877 3574 46079 3576
rect 3877 3571 3943 3574
rect 46013 3571 46079 3574
rect 3417 3498 3483 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3348 800 3438
rect 3417 3435 3483 3438
rect 17585 3498 17651 3501
rect 46657 3498 46723 3501
rect 17585 3496 46723 3498
rect 17585 3440 17590 3496
rect 17646 3440 46662 3496
rect 46718 3440 46723 3496
rect 17585 3438 46723 3440
rect 17585 3435 17651 3438
rect 46657 3435 46723 3438
rect 47945 3498 48011 3501
rect 49200 3498 50000 3588
rect 47945 3496 50000 3498
rect 47945 3440 47950 3496
rect 48006 3440 50000 3496
rect 47945 3438 50000 3440
rect 47945 3435 48011 3438
rect 49200 3348 50000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 0 2668 800 2908
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 4061 1458 4127 1461
rect 0 1456 4127 1458
rect 0 1400 4066 1456
rect 4122 1400 4127 1456
rect 0 1398 4127 1400
rect 0 1308 800 1398
rect 4061 1395 4127 1398
rect 47761 1458 47827 1461
rect 49200 1458 50000 1548
rect 47761 1456 50000 1458
rect 47761 1400 47766 1456
rect 47822 1400 50000 1456
rect 47761 1398 50000 1400
rect 47761 1395 47827 1398
rect 49200 1308 50000 1398
rect 0 778 800 868
rect 2957 778 3023 781
rect 0 776 3023 778
rect 0 720 2962 776
rect 3018 720 3023 776
rect 0 718 3023 720
rect 0 628 800 718
rect 2957 715 3023 718
rect 48037 778 48103 781
rect 49200 778 50000 868
rect 48037 776 50000 778
rect 48037 720 48042 776
rect 48098 720 50000 776
rect 48037 718 50000 720
rect 48037 715 48103 718
rect 49200 628 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 188
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 28764 47016 28828 47020
rect 28764 46960 28778 47016
rect 28778 46960 28828 47016
rect 28764 46956 28828 46960
rect 46060 46956 46124 47020
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 46244 31316 46308 31380
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 28764 21932 28828 21996
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 46244 21524 46308 21588
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 46060 19756 46124 19820
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 28763 47020 28829 47021
rect 28763 46956 28764 47020
rect 28828 46956 28829 47020
rect 28763 46955 28829 46956
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 28766 21997 28826 46955
rect 34928 46272 35248 47296
rect 46059 47020 46125 47021
rect 46059 46956 46060 47020
rect 46124 46956 46125 47020
rect 46059 46955 46125 46956
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 28763 21996 28829 21997
rect 28763 21932 28764 21996
rect 28828 21932 28829 21996
rect 28763 21931 28829 21932
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 46062 19821 46122 46955
rect 46243 31380 46309 31381
rect 46243 31316 46244 31380
rect 46308 31316 46309 31380
rect 46243 31315 46309 31316
rect 46246 21589 46306 31315
rect 46243 21588 46309 21589
rect 46243 21524 46244 21588
rect 46308 21524 46309 21588
rect 46243 21523 46309 21524
rect 46059 19820 46125 19821
rect 46059 19756 46060 19820
rect 46124 19756 46125 19820
rect 46059 19755 46125 19756
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 40112 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 44528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform -1 0 29072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 29900 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 23736 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 33304 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 43792 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 38640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform 1 0 27876 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform 1 0 35604 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1644511149
transform 1 0 28888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1644511149
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_89
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1644511149
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1644511149
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_205
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1644511149
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 1644511149
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1644511149
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1644511149
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_314
timestamp 1644511149
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1644511149
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1644511149
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_430
timestamp 1644511149
transform 1 0 40664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1644511149
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1644511149
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_455
timestamp 1644511149
transform 1 0 42964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_9
timestamp 1644511149
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_31
timestamp 1644511149
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_43
timestamp 1644511149
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_63
timestamp 1644511149
transform 1 0 6900 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_71
timestamp 1644511149
transform 1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_95
timestamp 1644511149
transform 1 0 9844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1644511149
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_176
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_183
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_191
timestamp 1644511149
transform 1 0 18676 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1644511149
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_229
timestamp 1644511149
transform 1 0 22172 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_251
timestamp 1644511149
transform 1 0 24196 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_259
timestamp 1644511149
transform 1 0 24932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_284
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_296
timestamp 1644511149
transform 1 0 28336 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_308
timestamp 1644511149
transform 1 0 29440 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_320
timestamp 1644511149
transform 1 0 30544 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_345
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1644511149
transform 1 0 35972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_399
timestamp 1644511149
transform 1 0 37812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_411
timestamp 1644511149
transform 1 0 38916 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_415
timestamp 1644511149
transform 1 0 39284 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_422
timestamp 1644511149
transform 1 0 39928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_434
timestamp 1644511149
transform 1 0 41032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1644511149
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_453
timestamp 1644511149
transform 1 0 42780 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_475
timestamp 1644511149
transform 1 0 44804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1644511149
transform 1 0 5520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_117
timestamp 1644511149
transform 1 0 11868 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_156
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_172
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_176
timestamp 1644511149
transform 1 0 17296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_183
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1644511149
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1644511149
transform 1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1644511149
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_217
timestamp 1644511149
transform 1 0 21068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_224
timestamp 1644511149
transform 1 0 21712 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_230
timestamp 1644511149
transform 1 0 22264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1644511149
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_256
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_264
timestamp 1644511149
transform 1 0 25392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_286
timestamp 1644511149
transform 1 0 27416 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_298
timestamp 1644511149
transform 1 0 28520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1644511149
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_350
timestamp 1644511149
transform 1 0 33304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1644511149
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_430
timestamp 1644511149
transform 1 0 40664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_452
timestamp 1644511149
transform 1 0 42688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_459
timestamp 1644511149
transform 1 0 43332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_466
timestamp 1644511149
transform 1 0 43976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1644511149
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_14
timestamp 1644511149
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_18
timestamp 1644511149
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_22
timestamp 1644511149
transform 1 0 3128 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_34
timestamp 1644511149
transform 1 0 4232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_46
timestamp 1644511149
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1644511149
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_67
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_79
timestamp 1644511149
transform 1 0 8372 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_83
timestamp 1644511149
transform 1 0 8740 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_87
timestamp 1644511149
transform 1 0 9108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_95
timestamp 1644511149
transform 1 0 9844 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_100
timestamp 1644511149
transform 1 0 10304 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_116
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_128
timestamp 1644511149
transform 1 0 12880 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_136
timestamp 1644511149
transform 1 0 13616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_175
timestamp 1644511149
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1644511149
transform 1 0 17572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_186
timestamp 1644511149
transform 1 0 18216 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_197
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_204
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_211
timestamp 1644511149
transform 1 0 20516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1644511149
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_242
timestamp 1644511149
transform 1 0 23368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_257
timestamp 1644511149
transform 1 0 24748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_396
timestamp 1644511149
transform 1 0 37536 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_408
timestamp 1644511149
transform 1 0 38640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_424
timestamp 1644511149
transform 1 0 40112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_433
timestamp 1644511149
transform 1 0 40940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_445
timestamp 1644511149
transform 1 0 42044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_465
timestamp 1644511149
transform 1 0 43884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_477
timestamp 1644511149
transform 1 0 44988 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_492
timestamp 1644511149
transform 1 0 46368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_92
timestamp 1644511149
transform 1 0 9568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_104
timestamp 1644511149
transform 1 0 10672 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_116
timestamp 1644511149
transform 1 0 11776 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_128
timestamp 1644511149
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_183
timestamp 1644511149
transform 1 0 17940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_200
timestamp 1644511149
transform 1 0 19504 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_217
timestamp 1644511149
transform 1 0 21068 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_224
timestamp 1644511149
transform 1 0 21712 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_231
timestamp 1644511149
transform 1 0 22356 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_238
timestamp 1644511149
transform 1 0 23000 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_269
timestamp 1644511149
transform 1 0 25852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_281
timestamp 1644511149
transform 1 0 26956 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_293
timestamp 1644511149
transform 1 0 28060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1644511149
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_393
timestamp 1644511149
transform 1 0 37260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_407
timestamp 1644511149
transform 1 0 38548 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_416
timestamp 1644511149
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_446
timestamp 1644511149
transform 1 0 42136 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_453
timestamp 1644511149
transform 1 0 42780 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_465
timestamp 1644511149
transform 1 0 43884 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_473
timestamp 1644511149
transform 1 0 44620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_498
timestamp 1644511149
transform 1 0 46920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_190
timestamp 1644511149
transform 1 0 18584 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_202
timestamp 1644511149
transform 1 0 19688 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_214
timestamp 1644511149
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1644511149
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_228
timestamp 1644511149
transform 1 0 22080 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_235
timestamp 1644511149
transform 1 0 22724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_247
timestamp 1644511149
transform 1 0 23828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_259
timestamp 1644511149
transform 1 0 24932 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1644511149
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_406
timestamp 1644511149
transform 1 0 38456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_410
timestamp 1644511149
transform 1 0 38824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_421
timestamp 1644511149
transform 1 0 39836 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_428
timestamp 1644511149
transform 1 0 40480 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_436
timestamp 1644511149
transform 1 0 41216 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_462
timestamp 1644511149
transform 1 0 43608 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_466
timestamp 1644511149
transform 1 0 43976 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_478
timestamp 1644511149
transform 1 0 45080 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_490
timestamp 1644511149
transform 1 0 46184 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1644511149
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_427
timestamp 1644511149
transform 1 0 40388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_439
timestamp 1644511149
transform 1 0 41492 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_451
timestamp 1644511149
transform 1 0 42596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_463
timestamp 1644511149
transform 1 0 43700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_481
timestamp 1644511149
transform 1 0 45356 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_496
timestamp 1644511149
transform 1 0 46736 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1644511149
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_492
timestamp 1644511149
transform 1 0 46368 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_500
timestamp 1644511149
transform 1 0 47104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_469
timestamp 1644511149
transform 1 0 44252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_474
timestamp 1644511149
transform 1 0 44712 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_482
timestamp 1644511149
transform 1 0 45448 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_489
timestamp 1644511149
transform 1 0 46092 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_501
timestamp 1644511149
transform 1 0 47196 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1644511149
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_505
timestamp 1644511149
transform 1 0 47564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_512
timestamp 1644511149
transform 1 0 48208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_492
timestamp 1644511149
transform 1 0 46368 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_499
timestamp 1644511149
transform 1 0 47012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_191
timestamp 1644511149
transform 1 0 18676 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_203
timestamp 1644511149
transform 1 0 19780 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_215
timestamp 1644511149
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1644511149
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_229
timestamp 1644511149
transform 1 0 22172 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_234
timestamp 1644511149
transform 1 0 22632 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 1644511149
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_173
timestamp 1644511149
transform 1 0 17020 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_180
timestamp 1644511149
transform 1 0 17664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_184
timestamp 1644511149
transform 1 0 18032 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1644511149
transform 1 0 18400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_213
timestamp 1644511149
transform 1 0 20700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1644511149
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_246
timestamp 1644511149
transform 1 0 23736 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_258
timestamp 1644511149
transform 1 0 24840 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_270
timestamp 1644511149
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1644511149
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_493
timestamp 1644511149
transform 1 0 46460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1644511149
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1644511149
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_182
timestamp 1644511149
transform 1 0 17848 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1644511149
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_216
timestamp 1644511149
transform 1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1644511149
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_172
timestamp 1644511149
transform 1 0 16928 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_180
timestamp 1644511149
transform 1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_213
timestamp 1644511149
transform 1 0 20700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1644511149
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_265
timestamp 1644511149
transform 1 0 25484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1644511149
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1644511149
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_149
timestamp 1644511149
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_170
timestamp 1644511149
transform 1 0 16744 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_176
timestamp 1644511149
transform 1 0 17296 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_182
timestamp 1644511149
transform 1 0 17848 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1644511149
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_201
timestamp 1644511149
transform 1 0 19596 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_208
timestamp 1644511149
transform 1 0 20240 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_214
timestamp 1644511149
transform 1 0 20792 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_235
timestamp 1644511149
transform 1 0 22724 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_274
timestamp 1644511149
transform 1 0 26312 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_286
timestamp 1644511149
transform 1 0 27416 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_298
timestamp 1644511149
transform 1 0 28520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1644511149
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_465
timestamp 1644511149
transform 1 0 43884 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_498
timestamp 1644511149
transform 1 0 46920 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_510
timestamp 1644511149
transform 1 0 48024 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_144
timestamp 1644511149
transform 1 0 14352 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1644511149
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_173
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1644511149
transform 1 0 17572 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_204
timestamp 1644511149
transform 1 0 19872 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_214
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1644511149
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_235
timestamp 1644511149
transform 1 0 22724 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_242
timestamp 1644511149
transform 1 0 23368 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1644511149
transform 1 0 24748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1644511149
transform 1 0 25852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1644511149
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_486
timestamp 1644511149
transform 1 0 45816 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_498
timestamp 1644511149
transform 1 0 46920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_167
timestamp 1644511149
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_174
timestamp 1644511149
transform 1 0 17112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_185
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1644511149
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_204
timestamp 1644511149
transform 1 0 19872 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_216
timestamp 1644511149
transform 1 0 20976 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_224
timestamp 1644511149
transform 1 0 21712 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_228
timestamp 1644511149
transform 1 0 22080 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_241
timestamp 1644511149
transform 1 0 23276 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1644511149
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_259
timestamp 1644511149
transform 1 0 24932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_263
timestamp 1644511149
transform 1 0 25300 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_267
timestamp 1644511149
transform 1 0 25668 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_279
timestamp 1644511149
transform 1 0 26772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_285
timestamp 1644511149
transform 1 0 27324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_297
timestamp 1644511149
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1644511149
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_312
timestamp 1644511149
transform 1 0 29808 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_324
timestamp 1644511149
transform 1 0 30912 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_336
timestamp 1644511149
transform 1 0 32016 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_348
timestamp 1644511149
transform 1 0 33120 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1644511149
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_480
timestamp 1644511149
transform 1 0 45264 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_488
timestamp 1644511149
transform 1 0 46000 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_28
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_40
timestamp 1644511149
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_145
timestamp 1644511149
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_151
timestamp 1644511149
transform 1 0 14996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1644511149
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_186
timestamp 1644511149
transform 1 0 18216 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_198
timestamp 1644511149
transform 1 0 19320 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_206
timestamp 1644511149
transform 1 0 20056 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_212
timestamp 1644511149
transform 1 0 20608 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_248
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_275
timestamp 1644511149
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_294
timestamp 1644511149
transform 1 0 28152 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_327
timestamp 1644511149
transform 1 0 31188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_456
timestamp 1644511149
transform 1 0 43056 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_460
timestamp 1644511149
transform 1 0 43424 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_482
timestamp 1644511149
transform 1 0 45448 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_493
timestamp 1644511149
transform 1 0 46460 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_14
timestamp 1644511149
transform 1 0 2392 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1644511149
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_152
timestamp 1644511149
transform 1 0 15088 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_164
timestamp 1644511149
transform 1 0 16192 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_172
timestamp 1644511149
transform 1 0 16928 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1644511149
transform 1 0 21160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_226
timestamp 1644511149
transform 1 0 21896 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_238
timestamp 1644511149
transform 1 0 23000 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_260
timestamp 1644511149
transform 1 0 25024 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_268
timestamp 1644511149
transform 1 0 25760 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_280
timestamp 1644511149
transform 1 0 26864 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_286
timestamp 1644511149
transform 1 0 27416 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_315
timestamp 1644511149
transform 1 0 30084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_337
timestamp 1644511149
transform 1 0 32108 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_349
timestamp 1644511149
transform 1 0 33212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1644511149
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_439
timestamp 1644511149
transform 1 0 41492 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_453
timestamp 1644511149
transform 1 0 42780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_467
timestamp 1644511149
transform 1 0 44068 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_482
timestamp 1644511149
transform 1 0 45448 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_490
timestamp 1644511149
transform 1 0 46184 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_129
timestamp 1644511149
transform 1 0 12972 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_133
timestamp 1644511149
transform 1 0 13340 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_145
timestamp 1644511149
transform 1 0 14444 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_157
timestamp 1644511149
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1644511149
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_251
timestamp 1644511149
transform 1 0 24196 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_258
timestamp 1644511149
transform 1 0 24840 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_270
timestamp 1644511149
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1644511149
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_290
timestamp 1644511149
transform 1 0 27784 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_315
timestamp 1644511149
transform 1 0 30084 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_322
timestamp 1644511149
transform 1 0 30728 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_434
timestamp 1644511149
transform 1 0 41032 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_453
timestamp 1644511149
transform 1 0 42780 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_459
timestamp 1644511149
transform 1 0 43332 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1644511149
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1644511149
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_144
timestamp 1644511149
transform 1 0 14352 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_152
timestamp 1644511149
transform 1 0 15088 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_164
timestamp 1644511149
transform 1 0 16192 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_172
timestamp 1644511149
transform 1 0 16928 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1644511149
transform 1 0 17480 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1644511149
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_205
timestamp 1644511149
transform 1 0 19964 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1644511149
transform 1 0 20424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_235
timestamp 1644511149
transform 1 0 22724 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1644511149
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_258
timestamp 1644511149
transform 1 0 24840 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_285
timestamp 1644511149
transform 1 0 27324 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_297
timestamp 1644511149
transform 1 0 28428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_338
timestamp 1644511149
transform 1 0 32200 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_350
timestamp 1644511149
transform 1 0 33304 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1644511149
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_466
timestamp 1644511149
transform 1 0 43976 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_474
timestamp 1644511149
transform 1 0 44712 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_480
timestamp 1644511149
transform 1 0 45264 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_487
timestamp 1644511149
transform 1 0 45908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1644511149
transform 1 0 1932 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_31
timestamp 1644511149
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_43
timestamp 1644511149
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_121
timestamp 1644511149
transform 1 0 12236 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_134
timestamp 1644511149
transform 1 0 13432 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_145
timestamp 1644511149
transform 1 0 14444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_154
timestamp 1644511149
transform 1 0 15272 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_176
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_180
timestamp 1644511149
transform 1 0 17664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_188
timestamp 1644511149
transform 1 0 18400 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_196
timestamp 1644511149
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_201
timestamp 1644511149
transform 1 0 19596 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_212
timestamp 1644511149
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_228
timestamp 1644511149
transform 1 0 22080 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_235
timestamp 1644511149
transform 1 0 22724 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_243
timestamp 1644511149
transform 1 0 23460 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_260
timestamp 1644511149
transform 1 0 25024 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_267
timestamp 1644511149
transform 1 0 25668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_289
timestamp 1644511149
transform 1 0 27692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_300
timestamp 1644511149
transform 1 0 28704 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_309
timestamp 1644511149
transform 1 0 29532 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_316
timestamp 1644511149
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1644511149
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_457
timestamp 1644511149
transform 1 0 43148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_462
timestamp 1644511149
transform 1 0 43608 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_474
timestamp 1644511149
transform 1 0 44712 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_483
timestamp 1644511149
transform 1 0 45540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_499
timestamp 1644511149
transform 1 0 47012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_512
timestamp 1644511149
transform 1 0 48208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_125
timestamp 1644511149
transform 1 0 12604 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_129
timestamp 1644511149
transform 1 0 12972 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_225
timestamp 1644511149
transform 1 0 21804 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_237
timestamp 1644511149
transform 1 0 22908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1644511149
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_258
timestamp 1644511149
transform 1 0 24840 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_283
timestamp 1644511149
transform 1 0 27140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_295
timestamp 1644511149
transform 1 0 28244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_313
timestamp 1644511149
transform 1 0 29900 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_335
timestamp 1644511149
transform 1 0 31924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_347
timestamp 1644511149
transform 1 0 33028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1644511149
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_453
timestamp 1644511149
transform 1 0 42780 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_466
timestamp 1644511149
transform 1 0 43976 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1644511149
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_481
timestamp 1644511149
transform 1 0 45356 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_511
timestamp 1644511149
transform 1 0 48116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_515
timestamp 1644511149
transform 1 0 48484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_101
timestamp 1644511149
transform 1 0 10396 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1644511149
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1644511149
transform 1 0 13340 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_144
timestamp 1644511149
transform 1 0 14352 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_156
timestamp 1644511149
transform 1 0 15456 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_160
timestamp 1644511149
transform 1 0 15824 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_177
timestamp 1644511149
transform 1 0 17388 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_183
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_187
timestamp 1644511149
transform 1 0 18308 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_199
timestamp 1644511149
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_203
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_209
timestamp 1644511149
transform 1 0 20332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1644511149
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_243
timestamp 1644511149
transform 1 0 23460 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_255
timestamp 1644511149
transform 1 0 24564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_262
timestamp 1644511149
transform 1 0 25208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_269
timestamp 1644511149
transform 1 0 25852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_284
timestamp 1644511149
transform 1 0 27232 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_292
timestamp 1644511149
transform 1 0 27968 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_298
timestamp 1644511149
transform 1 0 28520 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_323
timestamp 1644511149
transform 1 0 30820 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_330
timestamp 1644511149
transform 1 0 31464 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1644511149
transform 1 0 32660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_355
timestamp 1644511149
transform 1 0 33764 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1644511149
transform 1 0 34868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_379
timestamp 1644511149
transform 1 0 35972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_452
timestamp 1644511149
transform 1 0 42688 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_469
timestamp 1644511149
transform 1 0 44252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_494
timestamp 1644511149
transform 1 0 46552 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_502
timestamp 1644511149
transform 1 0 47288 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_511
timestamp 1644511149
transform 1 0 48116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_515
timestamp 1644511149
transform 1 0 48484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_106
timestamp 1644511149
transform 1 0 10856 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_118
timestamp 1644511149
transform 1 0 11960 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_130
timestamp 1644511149
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1644511149
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_173
timestamp 1644511149
transform 1 0 17020 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_200
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_212
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_224
timestamp 1644511149
transform 1 0 21712 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_282
timestamp 1644511149
transform 1 0 27048 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_288
timestamp 1644511149
transform 1 0 27600 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_292
timestamp 1644511149
transform 1 0 27968 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_328
timestamp 1644511149
transform 1 0 31280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_369
timestamp 1644511149
transform 1 0 35052 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_379
timestamp 1644511149
transform 1 0 35972 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_391
timestamp 1644511149
transform 1 0 37076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_403
timestamp 1644511149
transform 1 0 38180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_415
timestamp 1644511149
transform 1 0 39284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_453
timestamp 1644511149
transform 1 0 42780 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_461
timestamp 1644511149
transform 1 0 43516 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_468
timestamp 1644511149
transform 1 0 44160 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_480
timestamp 1644511149
transform 1 0 45264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_487
timestamp 1644511149
transform 1 0 45908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_102
timestamp 1644511149
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1644511149
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_117
timestamp 1644511149
transform 1 0 11868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_129
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_138
timestamp 1644511149
transform 1 0 13800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_163
timestamp 1644511149
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_173
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_202
timestamp 1644511149
transform 1 0 19688 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_210
timestamp 1644511149
transform 1 0 20424 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_246
timestamp 1644511149
transform 1 0 23736 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_258
timestamp 1644511149
transform 1 0 24840 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1644511149
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1644511149
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_306
timestamp 1644511149
transform 1 0 29256 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_318
timestamp 1644511149
transform 1 0 30360 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1644511149
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_340
timestamp 1644511149
transform 1 0 32384 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_348
timestamp 1644511149
transform 1 0 33120 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_352
timestamp 1644511149
transform 1 0 33488 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_360
timestamp 1644511149
transform 1 0 34224 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_453
timestamp 1644511149
transform 1 0 42780 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_457
timestamp 1644511149
transform 1 0 43148 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_468
timestamp 1644511149
transform 1 0 44160 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_475
timestamp 1644511149
transform 1 0 44804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1644511149
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1644511149
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_88
timestamp 1644511149
transform 1 0 9200 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_96
timestamp 1644511149
transform 1 0 9936 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1644511149
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_126
timestamp 1644511149
transform 1 0 12696 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_132
timestamp 1644511149
transform 1 0 13248 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_162
timestamp 1644511149
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_170
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_176
timestamp 1644511149
transform 1 0 17296 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_184
timestamp 1644511149
transform 1 0 18032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1644511149
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1644511149
transform 1 0 20700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_235
timestamp 1644511149
transform 1 0 22724 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_242
timestamp 1644511149
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1644511149
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_281
timestamp 1644511149
transform 1 0 26956 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1644511149
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1644511149
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_368
timestamp 1644511149
transform 1 0 34960 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_380
timestamp 1644511149
transform 1 0 36064 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_392
timestamp 1644511149
transform 1 0 37168 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_404
timestamp 1644511149
transform 1 0 38272 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1644511149
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_430
timestamp 1644511149
transform 1 0 40664 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_442
timestamp 1644511149
transform 1 0 41768 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_450
timestamp 1644511149
transform 1 0 42504 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_455
timestamp 1644511149
transform 1 0 42964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_466
timestamp 1644511149
transform 1 0 43976 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_474
timestamp 1644511149
transform 1 0 44712 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_484
timestamp 1644511149
transform 1 0 45632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_498
timestamp 1644511149
transform 1 0 46920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_88
timestamp 1644511149
transform 1 0 9200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_99
timestamp 1644511149
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_106
timestamp 1644511149
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_116
timestamp 1644511149
transform 1 0 11776 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_143
timestamp 1644511149
transform 1 0 14260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_155
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_190
timestamp 1644511149
transform 1 0 18584 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_198
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_213
timestamp 1644511149
transform 1 0 20700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_229
timestamp 1644511149
transform 1 0 22172 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_258
timestamp 1644511149
transform 1 0 24840 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1644511149
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_284
timestamp 1644511149
transform 1 0 27232 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_292
timestamp 1644511149
transform 1 0 27968 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_296
timestamp 1644511149
transform 1 0 28336 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_309
timestamp 1644511149
transform 1 0 29532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_323
timestamp 1644511149
transform 1 0 30820 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1644511149
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_352
timestamp 1644511149
transform 1 0 33488 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_364
timestamp 1644511149
transform 1 0 34592 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_376
timestamp 1644511149
transform 1 0 35696 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1644511149
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_421
timestamp 1644511149
transform 1 0 39836 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_424
timestamp 1644511149
transform 1 0 40112 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_432
timestamp 1644511149
transform 1 0 40848 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1644511149
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_457
timestamp 1644511149
transform 1 0 43148 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_465
timestamp 1644511149
transform 1 0 43884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_478
timestamp 1644511149
transform 1 0 45080 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_493
timestamp 1644511149
transform 1 0 46460 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1644511149
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1644511149
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_144
timestamp 1644511149
transform 1 0 14352 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_173
timestamp 1644511149
transform 1 0 17020 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_180
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_205
timestamp 1644511149
transform 1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_213
timestamp 1644511149
transform 1 0 20700 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_236
timestamp 1644511149
transform 1 0 22816 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_261
timestamp 1644511149
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_282
timestamp 1644511149
transform 1 0 27048 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_298
timestamp 1644511149
transform 1 0 28520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1644511149
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_317
timestamp 1644511149
transform 1 0 30268 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_325
timestamp 1644511149
transform 1 0 31004 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_329
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_400
timestamp 1644511149
transform 1 0 37904 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_412
timestamp 1644511149
transform 1 0 39008 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_428
timestamp 1644511149
transform 1 0 40480 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_453
timestamp 1644511149
transform 1 0 42780 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_464
timestamp 1644511149
transform 1 0 43792 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_468
timestamp 1644511149
transform 1 0 44160 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_472
timestamp 1644511149
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_487
timestamp 1644511149
transform 1 0 45908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_19
timestamp 1644511149
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_31
timestamp 1644511149
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_43
timestamp 1644511149
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_85
timestamp 1644511149
transform 1 0 8924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_97
timestamp 1644511149
transform 1 0 10028 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1644511149
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_119
timestamp 1644511149
transform 1 0 12052 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_131
timestamp 1644511149
transform 1 0 13156 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_135
timestamp 1644511149
transform 1 0 13524 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_157
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1644511149
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_172
timestamp 1644511149
transform 1 0 16928 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_180
timestamp 1644511149
transform 1 0 17664 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_186
timestamp 1644511149
transform 1 0 18216 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_190
timestamp 1644511149
transform 1 0 18584 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_198
timestamp 1644511149
transform 1 0 19320 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_204
timestamp 1644511149
transform 1 0 19872 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1644511149
transform 1 0 20240 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_229
timestamp 1644511149
transform 1 0 22172 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_255
timestamp 1644511149
transform 1 0 24564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_267
timestamp 1644511149
transform 1 0 25668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_289
timestamp 1644511149
transform 1 0 27692 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_297
timestamp 1644511149
transform 1 0 28428 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_309
timestamp 1644511149
transform 1 0 29532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_314
timestamp 1644511149
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_323
timestamp 1644511149
transform 1 0 30820 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_331
timestamp 1644511149
transform 1 0 31556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_343
timestamp 1644511149
transform 1 0 32660 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_347
timestamp 1644511149
transform 1 0 33028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_355
timestamp 1644511149
transform 1 0 33764 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_367
timestamp 1644511149
transform 1 0 34868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_371
timestamp 1644511149
transform 1 0 35236 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1644511149
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_425
timestamp 1644511149
transform 1 0 40204 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_434
timestamp 1644511149
transform 1 0 41032 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_446
timestamp 1644511149
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_458
timestamp 1644511149
transform 1 0 43240 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_475
timestamp 1644511149
transform 1 0 44804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_510
timestamp 1644511149
transform 1 0 48024 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_108
timestamp 1644511149
transform 1 0 11040 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1644511149
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_127
timestamp 1644511149
transform 1 0 12788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1644511149
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 1644511149
transform 1 0 14444 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_161
timestamp 1644511149
transform 1 0 15916 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_169
timestamp 1644511149
transform 1 0 16652 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_175
timestamp 1644511149
transform 1 0 17204 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_183
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_201
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_226
timestamp 1644511149
transform 1 0 21896 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_238
timestamp 1644511149
transform 1 0 23000 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_274
timestamp 1644511149
transform 1 0 26312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_285
timestamp 1644511149
transform 1 0 27324 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_293
timestamp 1644511149
transform 1 0 28060 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_312
timestamp 1644511149
transform 1 0 29808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_320
timestamp 1644511149
transform 1 0 30544 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_328
timestamp 1644511149
transform 1 0 31280 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_350
timestamp 1644511149
transform 1 0 33304 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1644511149
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_373
timestamp 1644511149
transform 1 0 35420 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_397
timestamp 1644511149
transform 1 0 37628 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_409
timestamp 1644511149
transform 1 0 38732 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_417
timestamp 1644511149
transform 1 0 39468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_428
timestamp 1644511149
transform 1 0 40480 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_432
timestamp 1644511149
transform 1 0 40848 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_440
timestamp 1644511149
transform 1 0 41584 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_452
timestamp 1644511149
transform 1 0 42688 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_458
timestamp 1644511149
transform 1 0 43240 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_462
timestamp 1644511149
transform 1 0 43608 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_472
timestamp 1644511149
transform 1 0 44528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_486
timestamp 1644511149
transform 1 0 45816 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1644511149
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_515
timestamp 1644511149
transform 1 0 48484 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_77
timestamp 1644511149
transform 1 0 8188 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_100
timestamp 1644511149
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_118
timestamp 1644511149
transform 1 0 11960 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_126
timestamp 1644511149
transform 1 0 12696 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_155
timestamp 1644511149
transform 1 0 15364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_195
timestamp 1644511149
transform 1 0 19044 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_241
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_253
timestamp 1644511149
transform 1 0 24380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_260
timestamp 1644511149
transform 1 0 25024 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_268
timestamp 1644511149
transform 1 0 25760 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_285
timestamp 1644511149
transform 1 0 27324 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_291
timestamp 1644511149
transform 1 0 27876 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_298
timestamp 1644511149
transform 1 0 28520 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_304
timestamp 1644511149
transform 1 0 29072 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_309
timestamp 1644511149
transform 1 0 29532 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_321
timestamp 1644511149
transform 1 0 30636 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1644511149
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_368
timestamp 1644511149
transform 1 0 34960 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_374
timestamp 1644511149
transform 1 0 35512 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_377
timestamp 1644511149
transform 1 0 35788 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_444
timestamp 1644511149
transform 1 0 41952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_457
timestamp 1644511149
transform 1 0 43148 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_463
timestamp 1644511149
transform 1 0 43700 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_471
timestamp 1644511149
transform 1 0 44436 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_476
timestamp 1644511149
transform 1 0 44896 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_13
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1644511149
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_113
timestamp 1644511149
transform 1 0 11500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_128
timestamp 1644511149
transform 1 0 12880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_132
timestamp 1644511149
transform 1 0 13248 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_146
timestamp 1644511149
transform 1 0 14536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_154
timestamp 1644511149
transform 1 0 15272 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_161
timestamp 1644511149
transform 1 0 15916 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_171
timestamp 1644511149
transform 1 0 16836 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_179
timestamp 1644511149
transform 1 0 17572 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_183
timestamp 1644511149
transform 1 0 17940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_227
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_257
timestamp 1644511149
transform 1 0 24748 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_263
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_270
timestamp 1644511149
transform 1 0 25944 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_287
timestamp 1644511149
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_303
timestamp 1644511149
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_317
timestamp 1644511149
transform 1 0 30268 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1644511149
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_335
timestamp 1644511149
transform 1 0 31924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_347
timestamp 1644511149
transform 1 0 33028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_355
timestamp 1644511149
transform 1 0 33764 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1644511149
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_385
timestamp 1644511149
transform 1 0 36524 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_397
timestamp 1644511149
transform 1 0 37628 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_409
timestamp 1644511149
transform 1 0 38732 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_417
timestamp 1644511149
transform 1 0 39468 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_485
timestamp 1644511149
transform 1 0 45724 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_99
timestamp 1644511149
transform 1 0 10212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_117
timestamp 1644511149
transform 1 0 11868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_133
timestamp 1644511149
transform 1 0 13340 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_141
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_146
timestamp 1644511149
transform 1 0 14536 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_157
timestamp 1644511149
transform 1 0 15548 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_179
timestamp 1644511149
transform 1 0 17572 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_187
timestamp 1644511149
transform 1 0 18308 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_199
timestamp 1644511149
transform 1 0 19412 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_207
timestamp 1644511149
transform 1 0 20148 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_233
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_238
timestamp 1644511149
transform 1 0 23000 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_251
timestamp 1644511149
transform 1 0 24196 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_259
timestamp 1644511149
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_271
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_285
timestamp 1644511149
transform 1 0 27324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_297
timestamp 1644511149
transform 1 0 28428 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_303
timestamp 1644511149
transform 1 0 28980 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_320
timestamp 1644511149
transform 1 0 30544 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_344
timestamp 1644511149
transform 1 0 32752 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_376
timestamp 1644511149
transform 1 0 35696 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1644511149
transform 1 0 36800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_492
timestamp 1644511149
transform 1 0 46368 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_499
timestamp 1644511149
transform 1 0 47012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_123
timestamp 1644511149
transform 1 0 12420 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1644511149
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_147
timestamp 1644511149
transform 1 0 14628 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_151
timestamp 1644511149
transform 1 0 14996 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_172
timestamp 1644511149
transform 1 0 16928 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_184
timestamp 1644511149
transform 1 0 18032 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_220
timestamp 1644511149
transform 1 0 21344 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_227
timestamp 1644511149
transform 1 0 21988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_239
timestamp 1644511149
transform 1 0 23092 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_261
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_273
timestamp 1644511149
transform 1 0 26220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_285
timestamp 1644511149
transform 1 0 27324 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_293
timestamp 1644511149
transform 1 0 28060 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_317
timestamp 1644511149
transform 1 0 30268 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_341
timestamp 1644511149
transform 1 0 32476 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_349
timestamp 1644511149
transform 1 0 33212 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1644511149
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_512
timestamp 1644511149
transform 1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_101
timestamp 1644511149
transform 1 0 10396 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_106
timestamp 1644511149
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_117
timestamp 1644511149
transform 1 0 11868 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_129
timestamp 1644511149
transform 1 0 12972 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_143
timestamp 1644511149
transform 1 0 14260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_151
timestamp 1644511149
transform 1 0 14996 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_156
timestamp 1644511149
transform 1 0 15456 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_173
timestamp 1644511149
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_177
timestamp 1644511149
transform 1 0 17388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_203
timestamp 1644511149
transform 1 0 19780 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_211
timestamp 1644511149
transform 1 0 20516 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1644511149
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_234
timestamp 1644511149
transform 1 0 22632 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_246
timestamp 1644511149
transform 1 0 23736 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_254
timestamp 1644511149
transform 1 0 24472 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_266
timestamp 1644511149
transform 1 0 25576 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_271
timestamp 1644511149
transform 1 0 26036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_287
timestamp 1644511149
transform 1 0 27508 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 1644511149
transform 1 0 28796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_308
timestamp 1644511149
transform 1 0 29440 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_320
timestamp 1644511149
transform 1 0 30544 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_344
timestamp 1644511149
transform 1 0 32752 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_350
timestamp 1644511149
transform 1 0 33304 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_360
timestamp 1644511149
transform 1 0 34224 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_372
timestamp 1644511149
transform 1 0 35328 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_384
timestamp 1644511149
transform 1 0 36432 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_508
timestamp 1644511149
transform 1 0 47840 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1644511149
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_95
timestamp 1644511149
transform 1 0 9844 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_103
timestamp 1644511149
transform 1 0 10580 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_117
timestamp 1644511149
transform 1 0 11868 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_162
timestamp 1644511149
transform 1 0 16008 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_170
timestamp 1644511149
transform 1 0 16744 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_185
timestamp 1644511149
transform 1 0 18124 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1644511149
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_216
timestamp 1644511149
transform 1 0 20976 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_227
timestamp 1644511149
transform 1 0 21988 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_236
timestamp 1644511149
transform 1 0 22816 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_261
timestamp 1644511149
transform 1 0 25116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_269
timestamp 1644511149
transform 1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_275
timestamp 1644511149
transform 1 0 26404 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_283
timestamp 1644511149
transform 1 0 27140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_287
timestamp 1644511149
transform 1 0 27508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_303
timestamp 1644511149
transform 1 0 28980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_316
timestamp 1644511149
transform 1 0 30176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_324
timestamp 1644511149
transform 1 0 30912 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_338
timestamp 1644511149
transform 1 0 32200 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_350
timestamp 1644511149
transform 1 0 33304 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1644511149
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1644511149
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_117
timestamp 1644511149
transform 1 0 11868 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_129
timestamp 1644511149
transform 1 0 12972 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_133
timestamp 1644511149
transform 1 0 13340 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_138
timestamp 1644511149
transform 1 0 13800 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_151
timestamp 1644511149
transform 1 0 14996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_175
timestamp 1644511149
transform 1 0 17204 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_183
timestamp 1644511149
transform 1 0 17940 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_209
timestamp 1644511149
transform 1 0 20332 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1644511149
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1644511149
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_231
timestamp 1644511149
transform 1 0 22356 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_241
timestamp 1644511149
transform 1 0 23276 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_253
timestamp 1644511149
transform 1 0 24380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_260
timestamp 1644511149
transform 1 0 25024 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_264
timestamp 1644511149
transform 1 0 25392 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_268
timestamp 1644511149
transform 1 0 25760 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_272
timestamp 1644511149
transform 1 0 26128 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_285
timestamp 1644511149
transform 1 0 27324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_300
timestamp 1644511149
transform 1 0 28704 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_307
timestamp 1644511149
transform 1 0 29348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_315
timestamp 1644511149
transform 1 0 30084 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_321
timestamp 1644511149
transform 1 0 30636 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_331
timestamp 1644511149
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_345
timestamp 1644511149
transform 1 0 32844 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_366
timestamp 1644511149
transform 1 0 34776 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_93
timestamp 1644511149
transform 1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_103
timestamp 1644511149
transform 1 0 10580 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_130
timestamp 1644511149
transform 1 0 13064 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1644511149
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_146
timestamp 1644511149
transform 1 0 14536 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_157
timestamp 1644511149
transform 1 0 15548 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_161
timestamp 1644511149
transform 1 0 15916 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_182
timestamp 1644511149
transform 1 0 17848 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_217
timestamp 1644511149
transform 1 0 21068 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_228
timestamp 1644511149
transform 1 0 22080 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_238
timestamp 1644511149
transform 1 0 23000 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1644511149
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_262
timestamp 1644511149
transform 1 0 25208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_266
timestamp 1644511149
transform 1 0 25576 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_271
timestamp 1644511149
transform 1 0 26036 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_283
timestamp 1644511149
transform 1 0 27140 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_293
timestamp 1644511149
transform 1 0 28060 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_297
timestamp 1644511149
transform 1 0 28428 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_316
timestamp 1644511149
transform 1 0 30176 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_324
timestamp 1644511149
transform 1 0 30912 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_335
timestamp 1644511149
transform 1 0 31924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_342
timestamp 1644511149
transform 1 0 32568 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_354
timestamp 1644511149
transform 1 0 33672 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1644511149
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_369
timestamp 1644511149
transform 1 0 35052 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_376
timestamp 1644511149
transform 1 0 35696 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_388
timestamp 1644511149
transform 1 0 36800 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_400
timestamp 1644511149
transform 1 0 37904 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_412
timestamp 1644511149
transform 1 0 39008 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_507
timestamp 1644511149
transform 1 0 47748 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_515
timestamp 1644511149
transform 1 0 48484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_89
timestamp 1644511149
transform 1 0 9292 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_95
timestamp 1644511149
transform 1 0 9844 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_107
timestamp 1644511149
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_145
timestamp 1644511149
transform 1 0 14444 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_160
timestamp 1644511149
transform 1 0 15824 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_174
timestamp 1644511149
transform 1 0 17112 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_186
timestamp 1644511149
transform 1 0 18216 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_198
timestamp 1644511149
transform 1 0 19320 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_210
timestamp 1644511149
transform 1 0 20424 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1644511149
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_230
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_242
timestamp 1644511149
transform 1 0 23368 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_250
timestamp 1644511149
transform 1 0 24104 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_289
timestamp 1644511149
transform 1 0 27692 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_311
timestamp 1644511149
transform 1 0 29716 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_319
timestamp 1644511149
transform 1 0 30452 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_326
timestamp 1644511149
transform 1 0 31096 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1644511149
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_341
timestamp 1644511149
transform 1 0 32476 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_347
timestamp 1644511149
transform 1 0 33028 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_354
timestamp 1644511149
transform 1 0 33672 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_380
timestamp 1644511149
transform 1 0 36064 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_110
timestamp 1644511149
transform 1 0 11224 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_122
timestamp 1644511149
transform 1 0 12328 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_134
timestamp 1644511149
transform 1 0 13432 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_159
timestamp 1644511149
transform 1 0 15732 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_183
timestamp 1644511149
transform 1 0 17940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_217
timestamp 1644511149
transform 1 0 21068 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_227
timestamp 1644511149
transform 1 0 21988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_239
timestamp 1644511149
transform 1 0 23092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_264
timestamp 1644511149
transform 1 0 25392 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_274
timestamp 1644511149
transform 1 0 26312 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_282
timestamp 1644511149
transform 1 0 27048 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1644511149
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_331
timestamp 1644511149
transform 1 0 31556 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_335
timestamp 1644511149
transform 1 0 31924 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_343
timestamp 1644511149
transform 1 0 32660 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_356
timestamp 1644511149
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_371
timestamp 1644511149
transform 1 0 35236 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_380
timestamp 1644511149
transform 1 0 36064 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_392
timestamp 1644511149
transform 1 0 37168 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_404
timestamp 1644511149
transform 1 0 38272 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_416
timestamp 1644511149
transform 1 0 39376 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_101
timestamp 1644511149
transform 1 0 10396 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1644511149
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_117
timestamp 1644511149
transform 1 0 11868 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_128
timestamp 1644511149
transform 1 0 12880 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_140
timestamp 1644511149
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_144
timestamp 1644511149
transform 1 0 14352 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_156
timestamp 1644511149
transform 1 0 15456 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_219
timestamp 1644511149
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_235
timestamp 1644511149
transform 1 0 22724 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_243
timestamp 1644511149
transform 1 0 23460 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_248
timestamp 1644511149
transform 1 0 23920 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_258
timestamp 1644511149
transform 1 0 24840 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_262
timestamp 1644511149
transform 1 0 25208 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_267
timestamp 1644511149
transform 1 0 25668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1644511149
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_292
timestamp 1644511149
transform 1 0 27968 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_308
timestamp 1644511149
transform 1 0 29440 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_345
timestamp 1644511149
transform 1 0 32844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_353
timestamp 1644511149
transform 1 0 33580 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_364
timestamp 1644511149
transform 1 0 34592 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1644511149
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_125
timestamp 1644511149
transform 1 0 12604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_136
timestamp 1644511149
transform 1 0 13616 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_145
timestamp 1644511149
transform 1 0 14444 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_157
timestamp 1644511149
transform 1 0 15548 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_179
timestamp 1644511149
transform 1 0 17572 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_191
timestamp 1644511149
transform 1 0 18676 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_217
timestamp 1644511149
transform 1 0 21068 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_225
timestamp 1644511149
transform 1 0 21804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_243
timestamp 1644511149
transform 1 0 23460 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_258
timestamp 1644511149
transform 1 0 24840 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_269
timestamp 1644511149
transform 1 0 25852 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_276
timestamp 1644511149
transform 1 0 26496 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_288
timestamp 1644511149
transform 1 0 27600 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_299
timestamp 1644511149
transform 1 0 28612 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_315
timestamp 1644511149
transform 1 0 30084 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_319
timestamp 1644511149
transform 1 0 30452 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_323
timestamp 1644511149
transform 1 0 30820 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_340
timestamp 1644511149
transform 1 0 32384 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_352
timestamp 1644511149
transform 1 0 33488 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1644511149
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_376
timestamp 1644511149
transform 1 0 35696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_388
timestamp 1644511149
transform 1 0 36800 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_400
timestamp 1644511149
transform 1 0 37904 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_412
timestamp 1644511149
transform 1 0 39008 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_9
timestamp 1644511149
transform 1 0 1932 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_31
timestamp 1644511149
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_43
timestamp 1644511149
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_101
timestamp 1644511149
transform 1 0 10396 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1644511149
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_124
timestamp 1644511149
transform 1 0 12512 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_136
timestamp 1644511149
transform 1 0 13616 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_157
timestamp 1644511149
transform 1 0 15548 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1644511149
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_172
timestamp 1644511149
transform 1 0 16928 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_184
timestamp 1644511149
transform 1 0 18032 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_192
timestamp 1644511149
transform 1 0 18768 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_213
timestamp 1644511149
transform 1 0 20700 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_236
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_246
timestamp 1644511149
transform 1 0 23736 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_270
timestamp 1644511149
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1644511149
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_345
timestamp 1644511149
transform 1 0 32844 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1644511149
transform 1 0 34868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1644511149
transform 1 0 35972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_500
timestamp 1644511149
transform 1 0 47104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_6
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_18
timestamp 1644511149
transform 1 0 2760 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_22
timestamp 1644511149
transform 1 0 3128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_96
timestamp 1644511149
transform 1 0 9936 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_107
timestamp 1644511149
transform 1 0 10948 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_118
timestamp 1644511149
transform 1 0 11960 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_127
timestamp 1644511149
transform 1 0 12788 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_134
timestamp 1644511149
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_147
timestamp 1644511149
transform 1 0 14628 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_154
timestamp 1644511149
transform 1 0 15272 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_166
timestamp 1644511149
transform 1 0 16376 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_178
timestamp 1644511149
transform 1 0 17480 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1644511149
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_208
timestamp 1644511149
transform 1 0 20240 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_216
timestamp 1644511149
transform 1 0 20976 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_224
timestamp 1644511149
transform 1 0 21712 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_230
timestamp 1644511149
transform 1 0 22264 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_238
timestamp 1644511149
transform 1 0 23000 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1644511149
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_260
timestamp 1644511149
transform 1 0 25024 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_266
timestamp 1644511149
transform 1 0 25576 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_274
timestamp 1644511149
transform 1 0 26312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_282
timestamp 1644511149
transform 1 0 27048 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_290
timestamp 1644511149
transform 1 0 27784 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_327
timestamp 1644511149
transform 1 0 31188 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_331
timestamp 1644511149
transform 1 0 31556 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_335
timestamp 1644511149
transform 1 0 31924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_368
timestamp 1644511149
transform 1 0 34960 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_380
timestamp 1644511149
transform 1 0 36064 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_392
timestamp 1644511149
transform 1 0 37168 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_404
timestamp 1644511149
transform 1 0 38272 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_416
timestamp 1644511149
transform 1 0 39376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_12
timestamp 1644511149
transform 1 0 2208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_37
timestamp 1644511149
transform 1 0 4508 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_49
timestamp 1644511149
transform 1 0 5612 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1644511149
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_134
timestamp 1644511149
transform 1 0 13432 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_143
timestamp 1644511149
transform 1 0 14260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_155
timestamp 1644511149
transform 1 0 15364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_213
timestamp 1644511149
transform 1 0 20700 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_230
timestamp 1644511149
transform 1 0 22264 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_242
timestamp 1644511149
transform 1 0 23368 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_254
timestamp 1644511149
transform 1 0 24472 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_260
timestamp 1644511149
transform 1 0 25024 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_268
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_286
timestamp 1644511149
transform 1 0 27416 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_294
timestamp 1644511149
transform 1 0 28152 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_299
timestamp 1644511149
transform 1 0 28612 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_307
timestamp 1644511149
transform 1 0 29348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_320
timestamp 1644511149
transform 1 0 30544 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_324
timestamp 1644511149
transform 1 0 30912 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_344
timestamp 1644511149
transform 1 0 32752 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_353
timestamp 1644511149
transform 1 0 33580 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_371
timestamp 1644511149
transform 1 0 35236 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_383
timestamp 1644511149
transform 1 0 36340 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_489
timestamp 1644511149
transform 1 0 46092 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_508
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_13
timestamp 1644511149
transform 1 0 2300 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_23
timestamp 1644511149
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1644511149
transform 1 0 4048 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1644511149
transform 1 0 5152 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1644511149
transform 1 0 6256 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_68
timestamp 1644511149
transform 1 0 7360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1644511149
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1644511149
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_162
timestamp 1644511149
transform 1 0 16008 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_174
timestamp 1644511149
transform 1 0 17112 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_186
timestamp 1644511149
transform 1 0 18216 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1644511149
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_222
timestamp 1644511149
transform 1 0 21528 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_235
timestamp 1644511149
transform 1 0 22724 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_247
timestamp 1644511149
transform 1 0 23828 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_262
timestamp 1644511149
transform 1 0 25208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_266
timestamp 1644511149
transform 1 0 25576 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_274
timestamp 1644511149
transform 1 0 26312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_285
timestamp 1644511149
transform 1 0 27324 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_291
timestamp 1644511149
transform 1 0 27876 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_297
timestamp 1644511149
transform 1 0 28428 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_315
timestamp 1644511149
transform 1 0 30084 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_326
timestamp 1644511149
transform 1 0 31096 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_338
timestamp 1644511149
transform 1 0 32200 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_346
timestamp 1644511149
transform 1 0 32936 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_354
timestamp 1644511149
transform 1 0 33672 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1644511149
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_385
timestamp 1644511149
transform 1 0 36524 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_397
timestamp 1644511149
transform 1 0 37628 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_409
timestamp 1644511149
transform 1 0 38732 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_417
timestamp 1644511149
transform 1 0 39468 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_495
timestamp 1644511149
transform 1 0 46644 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_30
timestamp 1644511149
transform 1 0 3864 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_42
timestamp 1644511149
transform 1 0 4968 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1644511149
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_199
timestamp 1644511149
transform 1 0 19412 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_234
timestamp 1644511149
transform 1 0 22632 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_246
timestamp 1644511149
transform 1 0 23736 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_260
timestamp 1644511149
transform 1 0 25024 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_271
timestamp 1644511149
transform 1 0 26036 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_298
timestamp 1644511149
transform 1 0 28520 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_314
timestamp 1644511149
transform 1 0 29992 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_323
timestamp 1644511149
transform 1 0 30820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_343
timestamp 1644511149
transform 1 0 32660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_351
timestamp 1644511149
transform 1 0 33396 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_363
timestamp 1644511149
transform 1 0 34500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_371
timestamp 1644511149
transform 1 0 35236 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_375
timestamp 1644511149
transform 1 0 35604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_387
timestamp 1644511149
transform 1 0 36708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_511
timestamp 1644511149
transform 1 0 48116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_515
timestamp 1644511149
transform 1 0 48484 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_214
timestamp 1644511149
transform 1 0 20792 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_240
timestamp 1644511149
transform 1 0 23184 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_258
timestamp 1644511149
transform 1 0 24840 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_266
timestamp 1644511149
transform 1 0 25576 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_274
timestamp 1644511149
transform 1 0 26312 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_286
timestamp 1644511149
transform 1 0 27416 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_298
timestamp 1644511149
transform 1 0 28520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1644511149
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_315
timestamp 1644511149
transform 1 0 30084 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_339
timestamp 1644511149
transform 1 0 32292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_351
timestamp 1644511149
transform 1 0 33396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_368
timestamp 1644511149
transform 1 0 34960 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_380
timestamp 1644511149
transform 1 0 36064 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_392
timestamp 1644511149
transform 1 0 37168 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_404
timestamp 1644511149
transform 1 0 38272 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_416
timestamp 1644511149
transform 1 0 39376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_507
timestamp 1644511149
transform 1 0 47748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_231
timestamp 1644511149
transform 1 0 22356 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_263
timestamp 1644511149
transform 1 0 25300 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_301
timestamp 1644511149
transform 1 0 28796 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_304
timestamp 1644511149
transform 1 0 29072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_314
timestamp 1644511149
transform 1 0 29992 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_327
timestamp 1644511149
transform 1 0 31188 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_345
timestamp 1644511149
transform 1 0 32844 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1644511149
transform 1 0 34868 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_379
timestamp 1644511149
transform 1 0 35972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_512
timestamp 1644511149
transform 1 0 48208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_215
timestamp 1644511149
transform 1 0 20884 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_227
timestamp 1644511149
transform 1 0 21988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_239
timestamp 1644511149
transform 1 0 23092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_259
timestamp 1644511149
transform 1 0 24932 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_267
timestamp 1644511149
transform 1 0 25668 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_286
timestamp 1644511149
transform 1 0 27416 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_290
timestamp 1644511149
transform 1 0 27784 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_297
timestamp 1644511149
transform 1 0 28428 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1644511149
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_317
timestamp 1644511149
transform 1 0 30268 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_328
timestamp 1644511149
transform 1 0 31280 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_340
timestamp 1644511149
transform 1 0 32384 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_353
timestamp 1644511149
transform 1 0 33580 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_361
timestamp 1644511149
transform 1 0 34316 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_236
timestamp 1644511149
transform 1 0 22816 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_248
timestamp 1644511149
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_252
timestamp 1644511149
transform 1 0 24288 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_257
timestamp 1644511149
transform 1 0 24748 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_265
timestamp 1644511149
transform 1 0 25484 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_303
timestamp 1644511149
transform 1 0 28980 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_327
timestamp 1644511149
transform 1 0 31188 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_359
timestamp 1644511149
transform 1 0 34132 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_371
timestamp 1644511149
transform 1 0 35236 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_383
timestamp 1644511149
transform 1 0 36340 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1644511149
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1644511149
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_227
timestamp 1644511149
transform 1 0 21988 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1644511149
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_273
timestamp 1644511149
transform 1 0 26220 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_285
timestamp 1644511149
transform 1 0 27324 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_297
timestamp 1644511149
transform 1 0 28428 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_352
timestamp 1644511149
transform 1 0 33488 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_30
timestamp 1644511149
transform 1 0 3864 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_42
timestamp 1644511149
transform 1 0 4968 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1644511149
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_241
timestamp 1644511149
transform 1 0 23276 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_253
timestamp 1644511149
transform 1 0 24380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_265
timestamp 1644511149
transform 1 0 25484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_290
timestamp 1644511149
transform 1 0 27784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_302
timestamp 1644511149
transform 1 0 28888 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_314
timestamp 1644511149
transform 1 0 29992 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_326
timestamp 1644511149
transform 1 0 31096 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1644511149
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_9
timestamp 1644511149
transform 1 0 1932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_13
timestamp 1644511149
transform 1 0 2300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp 1644511149
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_272
timestamp 1644511149
transform 1 0 26128 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_284
timestamp 1644511149
transform 1 0 27232 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_296
timestamp 1644511149
transform 1 0 28336 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_432
timestamp 1644511149
transform 1 0 40848 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_444
timestamp 1644511149
transform 1 0 41952 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_456
timestamp 1644511149
transform 1 0 43056 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_468
timestamp 1644511149
transform 1 0 44160 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_507
timestamp 1644511149
transform 1 0 47748 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_515
timestamp 1644511149
transform 1 0 48484 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_435
timestamp 1644511149
transform 1 0 41124 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_409
timestamp 1644511149
transform 1 0 38732 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_416
timestamp 1644511149
transform 1 0 39376 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_435
timestamp 1644511149
transform 1 0 41124 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_500
timestamp 1644511149
transform 1 0 47104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_428
timestamp 1644511149
transform 1 0 40480 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_440
timestamp 1644511149
transform 1 0 41584 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_452
timestamp 1644511149
transform 1 0 42688 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_464
timestamp 1644511149
transform 1 0 43792 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_7
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 1644511149
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_14
timestamp 1644511149
transform 1 0 2392 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_26
timestamp 1644511149
transform 1 0 3496 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_38
timestamp 1644511149
transform 1 0 4600 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_50
timestamp 1644511149
transform 1 0 5704 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_500
timestamp 1644511149
transform 1 0 47104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1644511149
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_9
timestamp 1644511149
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_21
timestamp 1644511149
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_437
timestamp 1644511149
transform 1 0 41308 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_442
timestamp 1644511149
transform 1 0 41768 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_481
timestamp 1644511149
transform 1 0 45356 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_485
timestamp 1644511149
transform 1 0 45724 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_489
timestamp 1644511149
transform 1 0 46092 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_297
timestamp 1644511149
transform 1 0 28428 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_303
timestamp 1644511149
transform 1 0 28980 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_412
timestamp 1644511149
transform 1 0 39008 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_437
timestamp 1644511149
transform 1 0 41308 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_459
timestamp 1644511149
transform 1 0 43332 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_467
timestamp 1644511149
transform 1 0 44068 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_9
timestamp 1644511149
transform 1 0 1932 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_31
timestamp 1644511149
transform 1 0 3956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_43
timestamp 1644511149
transform 1 0 5060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_101
timestamp 1644511149
transform 1 0 10396 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_106
timestamp 1644511149
transform 1 0 10856 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_211
timestamp 1644511149
transform 1 0 20516 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_218
timestamp 1644511149
transform 1 0 21160 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_266
timestamp 1644511149
transform 1 0 25576 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1644511149
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_352
timestamp 1644511149
transform 1 0 33488 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_364
timestamp 1644511149
transform 1 0 34592 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_376
timestamp 1644511149
transform 1 0 35696 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1644511149
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_436
timestamp 1644511149
transform 1 0 41216 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_443
timestamp 1644511149
transform 1 0 41860 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1644511149
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_461
timestamp 1644511149
transform 1 0 43516 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_467
timestamp 1644511149
transform 1 0 44068 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_492
timestamp 1644511149
transform 1 0 46368 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1644511149
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_508
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_22
timestamp 1644511149
transform 1 0 3128 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_32
timestamp 1644511149
transform 1 0 4048 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_39
timestamp 1644511149
transform 1 0 4692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_51
timestamp 1644511149
transform 1 0 5796 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_63
timestamp 1644511149
transform 1 0 6900 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_75
timestamp 1644511149
transform 1 0 8004 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_101
timestamp 1644511149
transform 1 0 10396 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_123
timestamp 1644511149
transform 1 0 12420 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1644511149
transform 1 0 13524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_205
timestamp 1644511149
transform 1 0 19964 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_210
timestamp 1644511149
transform 1 0 20424 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_235
timestamp 1644511149
transform 1 0 22724 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_247
timestamp 1644511149
transform 1 0 23828 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_258
timestamp 1644511149
transform 1 0 24840 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_283
timestamp 1644511149
transform 1 0 27140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_295
timestamp 1644511149
transform 1 0 28244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_344
timestamp 1644511149
transform 1 0 32752 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_356
timestamp 1644511149
transform 1 0 33856 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_407
timestamp 1644511149
transform 1 0 38548 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1644511149
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_437
timestamp 1644511149
transform 1 0 41308 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_459
timestamp 1644511149
transform 1 0 43332 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_466
timestamp 1644511149
transform 1 0 43976 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_474
timestamp 1644511149
transform 1 0 44712 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_13
timestamp 1644511149
transform 1 0 2300 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_20
timestamp 1644511149
transform 1 0 2944 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_24
timestamp 1644511149
transform 1 0 3312 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_46
timestamp 1644511149
transform 1 0 5336 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1644511149
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_101
timestamp 1644511149
transform 1 0 10396 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_106
timestamp 1644511149
transform 1 0 10856 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_131
timestamp 1644511149
transform 1 0 13156 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_156
timestamp 1644511149
transform 1 0 15456 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_228
timestamp 1644511149
transform 1 0 22080 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_240
timestamp 1644511149
transform 1 0 23184 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_252
timestamp 1644511149
transform 1 0 24288 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_424
timestamp 1644511149
transform 1 0 40112 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_436
timestamp 1644511149
transform 1 0 41216 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1644511149
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_449
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_473
timestamp 1644511149
transform 1 0 44620 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1644511149
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_63
timestamp 1644511149
transform 1 0 6900 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_71
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_117
timestamp 1644511149
transform 1 0 11868 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1644511149
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_149
timestamp 1644511149
transform 1 0 14812 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_161
timestamp 1644511149
transform 1 0 15916 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_185
timestamp 1644511149
transform 1 0 18124 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_192
timestamp 1644511149
transform 1 0 18768 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_216
timestamp 1644511149
transform 1 0 20976 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_259
timestamp 1644511149
transform 1 0 24932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_266
timestamp 1644511149
transform 1 0 25576 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1644511149
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1644511149
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_323
timestamp 1644511149
transform 1 0 30820 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_329
timestamp 1644511149
transform 1 0 31372 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_335
timestamp 1644511149
transform 1 0 31924 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_406
timestamp 1644511149
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_418
timestamp 1644511149
transform 1 0 39560 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_441
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_447
timestamp 1644511149
transform 1 0 42228 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_453
timestamp 1644511149
transform 1 0 42780 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_461
timestamp 1644511149
transform 1 0 43516 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1644511149
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1644511149
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_512
timestamp 1644511149
transform 1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0591_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13432 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31372 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0597_
timestamp 1644511149
transform 1 0 26036 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0598_
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0599_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0600_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0601_
timestamp 1644511149
transform 1 0 25668 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0602_
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0603_
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21252 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0605_
timestamp 1644511149
transform 1 0 22356 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0606_
timestamp 1644511149
transform 1 0 23460 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0607_
timestamp 1644511149
transform 1 0 21344 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0608_
timestamp 1644511149
transform 1 0 26772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1644511149
transform 1 0 28704 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0611_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18676 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0613_
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0614_
timestamp 1644511149
transform 1 0 12880 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0615_
timestamp 1644511149
transform 1 0 22816 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0616_
timestamp 1644511149
transform 1 0 17112 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22172 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0618_
timestamp 1644511149
transform 1 0 12972 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0619_
timestamp 1644511149
transform 1 0 14904 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0620_
timestamp 1644511149
transform 1 0 14904 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _0621_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _0622_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19412 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0623_
timestamp 1644511149
transform 1 0 20700 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22172 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0626_
timestamp 1644511149
transform 1 0 19872 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0627_
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1644511149
transform 1 0 22448 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0629_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0630_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1644511149
transform 1 0 18032 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0632_
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0634_
timestamp 1644511149
transform 1 0 18308 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0635_
timestamp 1644511149
transform 1 0 18952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0636_
timestamp 1644511149
transform 1 0 18400 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0637_
timestamp 1644511149
transform 1 0 16468 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0639_
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1644511149
transform 1 0 17664 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0641_
timestamp 1644511149
transform 1 0 17572 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0642_
timestamp 1644511149
transform 1 0 17940 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0644_
timestamp 1644511149
transform 1 0 14536 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0646_
timestamp 1644511149
transform 1 0 14168 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0647_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0648_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0649_
timestamp 1644511149
transform 1 0 13340 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0650_
timestamp 1644511149
transform 1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1644511149
transform 1 0 15640 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1644511149
transform 1 0 17112 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0653_
timestamp 1644511149
transform 1 0 14352 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15364 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0655_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0656_
timestamp 1644511149
transform 1 0 14076 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1644511149
transform 1 0 16836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0658_
timestamp 1644511149
transform 1 0 15180 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0661_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14536 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1644511149
transform 1 0 14996 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0663_
timestamp 1644511149
transform 1 0 12236 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0664_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1644511149
transform 1 0 12236 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0666_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10580 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0667_
timestamp 1644511149
transform 1 0 11592 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1644511149
transform 1 0 12512 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0669_
timestamp 1644511149
transform 1 0 13156 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0670_
timestamp 1644511149
transform 1 0 11316 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0671_
timestamp 1644511149
transform 1 0 13156 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1644511149
transform 1 0 11960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0673_
timestamp 1644511149
transform 1 0 9936 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1644511149
transform 1 0 11592 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0675_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0676_
timestamp 1644511149
transform 1 0 12328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0677_
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0678_
timestamp 1644511149
transform 1 0 10856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0680_
timestamp 1644511149
transform 1 0 12328 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0681_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10304 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1644511149
transform 1 0 12328 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0683_
timestamp 1644511149
transform 1 0 11408 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0684_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0687_
timestamp 1644511149
transform 1 0 9568 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0688_
timestamp 1644511149
transform 1 0 15088 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1644511149
transform 1 0 12696 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1644511149
transform 1 0 14628 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0691_
timestamp 1644511149
transform 1 0 13800 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0692_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1644511149
transform 1 0 13064 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0694_
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0695_
timestamp 1644511149
transform 1 0 12788 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1644511149
transform 1 0 15640 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0697_
timestamp 1644511149
transform 1 0 14720 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0698_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1644511149
transform 1 0 15364 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0700_
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1644511149
transform 1 0 16836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0702_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0703_
timestamp 1644511149
transform 1 0 23276 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0704_
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0705_
timestamp 1644511149
transform 1 0 15456 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0706_
timestamp 1644511149
transform 1 0 24656 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0707_
timestamp 1644511149
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1644511149
transform 1 0 19964 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0709_
timestamp 1644511149
transform 1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0710_
timestamp 1644511149
transform 1 0 17848 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1644511149
transform 1 0 19596 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0712_
timestamp 1644511149
transform 1 0 17480 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1644511149
transform 1 0 21804 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0714_
timestamp 1644511149
transform 1 0 23276 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0715_
timestamp 1644511149
transform 1 0 22356 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0716_
timestamp 1644511149
transform 1 0 23092 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1644511149
transform 1 0 25208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0718_
timestamp 1644511149
transform 1 0 23276 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1644511149
transform 1 0 25392 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0720_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0721_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0722_
timestamp 1644511149
transform 1 0 24564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0723_
timestamp 1644511149
transform 1 0 26680 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0725_
timestamp 1644511149
transform 1 0 25392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0726_
timestamp 1644511149
transform 1 0 24380 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0729_
timestamp 1644511149
transform 1 0 23552 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0730_
timestamp 1644511149
transform 1 0 25576 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1644511149
transform 1 0 28428 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0732_
timestamp 1644511149
transform 1 0 21896 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0733_
timestamp 1644511149
transform 1 0 23184 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23828 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1644511149
transform 1 0 29072 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0736_
timestamp 1644511149
transform 1 0 27692 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0737_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0738_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0739_
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0740_
timestamp 1644511149
transform 1 0 29900 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0741_
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0742_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0743_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0745_
timestamp 1644511149
transform 1 0 28612 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0746_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0747_
timestamp 1644511149
transform 1 0 24472 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0748_
timestamp 1644511149
transform 1 0 25668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0749_
timestamp 1644511149
transform 1 0 28244 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0750_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27600 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0751_
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0752_
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1644511149
transform 1 0 21712 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0754_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0755_
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0756_
timestamp 1644511149
transform 1 0 27600 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0757_
timestamp 1644511149
transform 1 0 28612 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _0758_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0759_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0760_
timestamp 1644511149
transform 1 0 33304 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _0761_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0762_
timestamp 1644511149
transform 1 0 30544 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0763_
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0764_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0765_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0766_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26680 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0767_
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0768_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0769_
timestamp 1644511149
transform 1 0 22908 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0770_
timestamp 1644511149
transform 1 0 21896 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0771_
timestamp 1644511149
transform 1 0 21896 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0772_
timestamp 1644511149
transform 1 0 28980 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0773_
timestamp 1644511149
transform 1 0 28612 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0774_
timestamp 1644511149
transform 1 0 31004 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0775_
timestamp 1644511149
transform 1 0 20884 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0776_
timestamp 1644511149
transform 1 0 20884 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0777_
timestamp 1644511149
transform 1 0 21896 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0778_
timestamp 1644511149
transform 1 0 23184 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0779_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0780_
timestamp 1644511149
transform 1 0 21252 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0782_
timestamp 1644511149
transform 1 0 26680 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0783_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0784_
timestamp 1644511149
transform 1 0 24656 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0785_
timestamp 1644511149
transform 1 0 22356 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0786_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _0787_
timestamp 1644511149
transform 1 0 25668 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0788_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0789_
timestamp 1644511149
transform 1 0 26956 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0790_
timestamp 1644511149
transform 1 0 25852 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0792_
timestamp 1644511149
transform 1 0 23000 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0793_
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0794_
timestamp 1644511149
transform 1 0 25852 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1644511149
transform 1 0 25668 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0796_
timestamp 1644511149
transform 1 0 26036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0797_
timestamp 1644511149
transform 1 0 25576 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0798_
timestamp 1644511149
transform 1 0 27416 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0799_
timestamp 1644511149
transform 1 0 26680 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0800_
timestamp 1644511149
transform 1 0 27968 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0801_
timestamp 1644511149
transform 1 0 27692 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0802_
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0803_
timestamp 1644511149
transform 1 0 28152 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0804_
timestamp 1644511149
transform 1 0 24104 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0805_
timestamp 1644511149
transform 1 0 24288 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0806_
timestamp 1644511149
transform 1 0 32476 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0807_
timestamp 1644511149
transform 1 0 30360 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0808_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29900 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0809_
timestamp 1644511149
transform 1 0 30268 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0810_
timestamp 1644511149
transform 1 0 29808 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0811_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29256 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0812_
timestamp 1644511149
transform 1 0 29256 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0813_
timestamp 1644511149
transform 1 0 33028 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0814_
timestamp 1644511149
transform 1 0 33304 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0815_
timestamp 1644511149
transform 1 0 33764 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0816_
timestamp 1644511149
transform 1 0 34408 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0817_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0818_
timestamp 1644511149
transform 1 0 31280 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0819_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0820_
timestamp 1644511149
transform 1 0 28520 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0821_
timestamp 1644511149
transform 1 0 33120 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28520 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0823_
timestamp 1644511149
transform 1 0 31004 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1644511149
transform 1 0 32292 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0825_
timestamp 1644511149
transform 1 0 30728 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0826_
timestamp 1644511149
transform 1 0 32936 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp 1644511149
transform 1 0 33304 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0828_
timestamp 1644511149
transform 1 0 33212 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0829_
timestamp 1644511149
transform 1 0 31464 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0830_
timestamp 1644511149
transform 1 0 31004 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0831_
timestamp 1644511149
transform 1 0 31464 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0832_
timestamp 1644511149
transform 1 0 30636 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0833_
timestamp 1644511149
transform 1 0 33120 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0834_
timestamp 1644511149
transform 1 0 32016 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0835_
timestamp 1644511149
transform 1 0 33028 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0836_
timestamp 1644511149
transform 1 0 33948 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1644511149
transform 1 0 33764 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0838_
timestamp 1644511149
transform 1 0 34868 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0839_
timestamp 1644511149
transform 1 0 30544 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0840_
timestamp 1644511149
transform 1 0 30544 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1644511149
transform 1 0 29716 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0842_
timestamp 1644511149
transform 1 0 29808 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0843_
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0844_
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0845_
timestamp 1644511149
transform 1 0 27324 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0846_
timestamp 1644511149
transform 1 0 25760 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0847_
timestamp 1644511149
transform 1 0 24748 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0848_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0849_
timestamp 1644511149
transform 1 0 25208 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0850_
timestamp 1644511149
transform 1 0 25668 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0851_
timestamp 1644511149
transform 1 0 24472 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0852_
timestamp 1644511149
transform 1 0 30360 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0853_
timestamp 1644511149
transform 1 0 31004 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0854_
timestamp 1644511149
transform 1 0 30912 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1644511149
transform 1 0 26128 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0856_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0857_
timestamp 1644511149
transform 1 0 33304 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0858_
timestamp 1644511149
transform 1 0 30084 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0859_
timestamp 1644511149
transform 1 0 30636 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29624 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0861_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0862_
timestamp 1644511149
transform 1 0 30176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0863_
timestamp 1644511149
transform 1 0 29624 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0864_
timestamp 1644511149
transform 1 0 30084 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0865_
timestamp 1644511149
transform 1 0 29716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0866_
timestamp 1644511149
transform 1 0 31188 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0867_
timestamp 1644511149
transform 1 0 30360 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0868_
timestamp 1644511149
transform 1 0 31188 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0869_
timestamp 1644511149
transform 1 0 31464 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0870_
timestamp 1644511149
transform 1 0 27968 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1644511149
transform 1 0 27968 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0872_
timestamp 1644511149
transform 1 0 28152 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0873_
timestamp 1644511149
transform 1 0 33396 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0874_
timestamp 1644511149
transform 1 0 26680 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0875_
timestamp 1644511149
transform 1 0 25852 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0876_
timestamp 1644511149
transform 1 0 25760 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0877_
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0878_
timestamp 1644511149
transform 1 0 28152 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0879_
timestamp 1644511149
transform 1 0 28888 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0880_
timestamp 1644511149
transform 1 0 28612 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1644511149
transform 1 0 27968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0882_
timestamp 1644511149
transform 1 0 26680 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0883_
timestamp 1644511149
transform 1 0 25392 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0884_
timestamp 1644511149
transform 1 0 35972 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _0885_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35972 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1644511149
transform 1 0 46736 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1644511149
transform 1 0 23092 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1644511149
transform 1 0 21896 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36156 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 43792 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform 1 0 2760 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0897_
timestamp 1644511149
transform 1 0 35328 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 2944 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1644511149
transform 1 0 20240 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0903_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 2116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0909_
timestamp 1644511149
transform 1 0 45356 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45264 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1644511149
transform 1 0 43700 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45448 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  _0917_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 41492 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1644511149
transform 1 0 43976 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0922_
timestamp 1644511149
transform 1 0 45080 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 27508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 28244 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45264 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1644511149
transform 1 0 46644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 46736 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1644511149
transform 1 0 45080 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0934_
timestamp 1644511149
transform 1 0 43976 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 40204 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 38732 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 46736 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1644511149
transform 1 0 39008 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0941_
timestamp 1644511149
transform 1 0 40020 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 20884 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0947_
timestamp 1644511149
transform 1 0 40020 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 10580 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 25300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 2852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0953_
timestamp 1644511149
transform 1 0 40204 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 2852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 43056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0959_
timestamp 1644511149
transform 1 0 40020 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 45632 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 46828 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 38272 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0965_
timestamp 1644511149
transform 1 0 39928 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 40940 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 31188 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 22356 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 20700 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0971_
timestamp 1644511149
transform 1 0 17940 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0972_
timestamp 1644511149
transform 1 0 17112 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 16744 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 17388 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0978_
timestamp 1644511149
transform 1 0 13892 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 8648 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 8924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform 1 0 13524 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0984_
timestamp 1644511149
transform 1 0 13892 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 9568 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 13984 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 9568 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1644511149
transform 1 0 9660 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0990_
timestamp 1644511149
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 17848 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1644511149
transform 1 0 18216 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0996_
timestamp 1644511149
transform 1 0 16744 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 19320 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 20424 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1644511149
transform 1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 35512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1003_
timestamp 1644511149
transform 1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1004_
timestamp 1644511149
transform 1 0 21528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__or2b_1  _1007_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31096 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1644511149
transform 1 0 30452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43240 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_2  _1010_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _1011_
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1012_
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1644511149
transform 1 0 45356 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1014_
timestamp 1644511149
transform 1 0 44804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1644511149
transform 1 0 44528 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1017_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1019_
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1020_
timestamp 1644511149
transform 1 0 40296 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1644511149
transform 1 0 40204 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1022_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40204 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1644511149
transform 1 0 40480 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1644511149
transform 1 0 40204 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1025_
timestamp 1644511149
transform 1 0 40020 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1644511149
transform 1 0 39652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1027_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1028_
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1030_
timestamp 1644511149
transform 1 0 25208 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1032_
timestamp 1644511149
transform 1 0 2668 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1034_
timestamp 1644511149
transform 1 0 44896 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1644511149
transform 1 0 45816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1036_
timestamp 1644511149
transform 1 0 33672 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1038_
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1040_
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1644511149
transform 1 0 42504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1042_
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1044_
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1045_
timestamp 1644511149
transform 1 0 28244 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1046_
timestamp 1644511149
transform 1 0 29072 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1644511149
transform 1 0 29900 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1049_
timestamp 1644511149
transform 1 0 27784 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1050_
timestamp 1644511149
transform 1 0 26864 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_4  _1051_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27508 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1052_
timestamp 1644511149
transform 1 0 40756 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1053_
timestamp 1644511149
transform 1 0 41400 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1054_
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1055_
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1056_
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1057_
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1058_
timestamp 1644511149
transform 1 0 43700 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1059_
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43424 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1061_
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1062_
timestamp 1644511149
transform 1 0 43056 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1063_
timestamp 1644511149
transform 1 0 43884 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_2  _1064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41860 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1065_
timestamp 1644511149
transform 1 0 43332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1066_
timestamp 1644511149
transform 1 0 43056 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1067_
timestamp 1644511149
transform 1 0 42688 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1068_
timestamp 1644511149
transform 1 0 42872 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1069_
timestamp 1644511149
transform 1 0 43332 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_2  _1070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43056 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _1071_
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1072_
timestamp 1644511149
transform 1 0 43332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1073_
timestamp 1644511149
transform 1 0 43332 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1074_
timestamp 1644511149
transform 1 0 43424 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1075_
timestamp 1644511149
transform 1 0 43332 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1076_
timestamp 1644511149
transform 1 0 43608 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _1077_
timestamp 1644511149
transform 1 0 42504 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1078_
timestamp 1644511149
transform 1 0 40388 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1079_
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1644511149
transform 1 0 27324 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1083_
timestamp 1644511149
transform 1 0 33396 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1644511149
transform 1 0 34684 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1644511149
transform 1 0 32752 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1644511149
transform 1 0 32476 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1089_
timestamp 1644511149
transform 1 0 25668 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1644511149
transform 1 0 26220 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1644511149
transform 1 0 25484 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1644511149
transform 1 0 32108 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1095_
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1644511149
transform 1 0 35420 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1644511149
transform 1 0 35144 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1099_
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1644511149
transform 1 0 35328 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1101_
timestamp 1644511149
transform 1 0 24380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1644511149
transform 1 0 30360 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1644511149
transform 1 0 24564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1105_
timestamp 1644511149
transform 1 0 28520 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1644511149
transform 1 0 24656 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1107_
timestamp 1644511149
transform 1 0 20516 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1644511149
transform 1 0 22540 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1644511149
transform 1 0 22080 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1644511149
transform 1 0 19964 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1111_
timestamp 1644511149
transform 1 0 20516 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1113_
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1644511149
transform 1 0 20424 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1644511149
transform 1 0 20700 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1644511149
transform 1 0 23368 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1644511149
transform 1 0 23000 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1644511149
transform 1 0 21896 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1119_
timestamp 1644511149
transform 1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1120_
timestamp 1644511149
transform 1 0 24472 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1121_
timestamp 1644511149
transform 1 0 24380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1644511149
transform 1 0 23736 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1123_
timestamp 1644511149
transform 1 0 20240 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1124_
timestamp 1644511149
transform 1 0 20424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1125_
timestamp 1644511149
transform 1 0 17848 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1126_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1127_
timestamp 1644511149
transform 1 0 14720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1128_
timestamp 1644511149
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1129_
timestamp 1644511149
transform 1 0 12328 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1130_
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1131_
timestamp 1644511149
transform 1 0 11868 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1132_
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1644511149
transform 1 0 10580 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1134_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1135_
timestamp 1644511149
transform 1 0 11868 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1644511149
transform 1 0 9936 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1137_
timestamp 1644511149
transform 1 0 10488 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1138_
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1644511149
transform 1 0 10672 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1140_
timestamp 1644511149
transform 1 0 10672 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1141_
timestamp 1644511149
transform 1 0 14904 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1142_
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1143_
timestamp 1644511149
transform 1 0 15548 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1144_
timestamp 1644511149
transform 1 0 15364 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1145_
timestamp 1644511149
transform 1 0 16376 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1146_
timestamp 1644511149
transform 1 0 15824 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1147_
timestamp 1644511149
transform 1 0 16376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1148_
timestamp 1644511149
transform 1 0 15548 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1149_
timestamp 1644511149
transform 1 0 16928 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1150_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1644511149
transform 1 0 17112 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1152_
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1153_
timestamp 1644511149
transform 1 0 20700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1154_
timestamp 1644511149
transform 1 0 19228 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1155_
timestamp 1644511149
transform 1 0 21344 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1157_
timestamp 1644511149
transform 1 0 27416 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1644511149
transform 1 0 25208 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1159_
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 1644511149
transform 1 0 32108 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 1644511149
transform 1 0 31464 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1162_
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1163_
timestamp 1644511149
transform 1 0 33856 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1164_
timestamp 1644511149
transform 1 0 24104 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1165_
timestamp 1644511149
transform 1 0 24288 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1166_
timestamp 1644511149
transform 1 0 27232 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1644511149
transform 1 0 34960 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1644511149
transform 1 0 34224 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1170_
timestamp 1644511149
transform 1 0 32936 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1644511149
transform 1 0 33028 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32936 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1173_
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 1644511149
transform 1 0 29348 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1175_
timestamp 1644511149
transform 1 0 30452 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1644511149
transform 1 0 23460 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 1644511149
transform 1 0 27140 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1178_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1179_
timestamp 1644511149
transform 1 0 22080 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1180_
timestamp 1644511149
transform 1 0 21344 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1181_
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 1644511149
transform 1 0 19504 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 1644511149
transform 1 0 19504 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 1644511149
transform 1 0 22724 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1187_
timestamp 1644511149
transform 1 0 22080 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1188_
timestamp 1644511149
transform 1 0 20884 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1189_
timestamp 1644511149
transform 1 0 25208 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1190_
timestamp 1644511149
transform 1 0 25392 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1191_
timestamp 1644511149
transform 1 0 24472 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1192_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1644511149
transform 1 0 20884 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1194_
timestamp 1644511149
transform 1 0 17940 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1196_
timestamp 1644511149
transform 1 0 14904 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14352 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 1644511149
transform 1 0 14444 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1199_
timestamp 1644511149
transform 1 0 11776 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1200_
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1201_
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1202_
timestamp 1644511149
transform 1 0 11408 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1203_
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1204_
timestamp 1644511149
transform 1 0 10580 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1205_
timestamp 1644511149
transform 1 0 10948 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1206_
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1644511149
transform 1 0 10764 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1208_
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1209_
timestamp 1644511149
transform 1 0 15640 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1210_
timestamp 1644511149
transform 1 0 16100 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1211_
timestamp 1644511149
transform 1 0 16008 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1644511149
transform 1 0 15088 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1213_
timestamp 1644511149
transform 1 0 15088 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1214_
timestamp 1644511149
transform 1 0 17204 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1215_
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1216_
timestamp 1644511149
transform 1 0 17848 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1217_
timestamp 1644511149
transform 1 0 16836 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1218_
timestamp 1644511149
transform 1 0 20792 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1644511149
transform 1 0 19964 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1220_
timestamp 1644511149
transform 1 0 22080 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _1221__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1222__82
timestamp 1644511149
transform 1 0 32476 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1223__83
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1224__84
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1225__85
timestamp 1644511149
transform 1 0 47472 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1226__86
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1227__87
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1228__88
timestamp 1644511149
transform 1 0 24656 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1229__89
timestamp 1644511149
transform 1 0 10580 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1230__90
timestamp 1644511149
transform 1 0 25300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1231__91
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1232__92
timestamp 1644511149
transform 1 0 2668 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1233__93
timestamp 1644511149
transform 1 0 33672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1234__94
timestamp 1644511149
transform 1 0 4416 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1235__95
timestamp 1644511149
transform 1 0 1932 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1236__96
timestamp 1644511149
transform 1 0 43700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1237__97
timestamp 1644511149
transform 1 0 45448 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1238__98
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1239__99
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1240__100
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1241__101
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1242__102
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1243__103
timestamp 1644511149
transform 1 0 41400 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1244__104
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1245__105
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1246__106
timestamp 1644511149
transform 1 0 22356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1247__107
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1248__108
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1249__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1250__110
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1251__111
timestamp 1644511149
transform 1 0 1472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1252__112
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1253__113
timestamp 1644511149
transform 1 0 41584 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1254__114
timestamp 1644511149
transform 1 0 45264 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1255__115
timestamp 1644511149
transform 1 0 25576 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1256__116
timestamp 1644511149
transform 1 0 42504 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1257__117
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1258__118
timestamp 1644511149
transform 1 0 12880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1259__119
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1260__120
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1261__121
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1262__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1263__123
timestamp 1644511149
transform 1 0 46368 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1264__124
timestamp 1644511149
transform 1 0 1472 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1265__125
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1266__126
timestamp 1644511149
transform 1 0 20148 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1267__127
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1268__128
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1269__129
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1270__130
timestamp 1644511149
transform 1 0 46092 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1271__131
timestamp 1644511149
transform 1 0 2024 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1272__132
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1273__133
timestamp 1644511149
transform 1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1274__134
timestamp 1644511149
transform 1 0 46184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1275__135
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28888 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1277_
timestamp 1644511149
transform 1 0 28152 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1278_
timestamp 1644511149
transform 1 0 43884 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1279_
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1280_
timestamp 1644511149
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1281_
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1282_
timestamp 1644511149
transform 1 0 46184 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1283_
timestamp 1644511149
transform 1 0 40020 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1284_
timestamp 1644511149
transform 1 0 38640 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1285_
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1286_
timestamp 1644511149
transform 1 0 32384 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1644511149
transform 1 0 20792 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1644511149
transform 1 0 10488 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1644511149
transform 1 0 25208 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1644511149
transform 1 0 2024 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1644511149
transform 1 0 32936 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1644511149
transform 1 0 3404 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1644511149
transform 1 0 2024 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1644511149
transform 1 0 42872 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1644511149
transform 1 0 38180 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 7912 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1644511149
transform 1 0 41400 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1644511149
transform 1 0 35972 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1309_
timestamp 1644511149
transform 1 0 29992 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1310_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1311_
timestamp 1644511149
transform 1 0 21988 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1312_
timestamp 1644511149
transform 1 0 22080 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1313_
timestamp 1644511149
transform 1 0 18768 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1314_
timestamp 1644511149
transform 1 0 16560 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1315_
timestamp 1644511149
transform 1 0 15916 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1316_
timestamp 1644511149
transform 1 0 16744 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1317_
timestamp 1644511149
transform 1 0 16928 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1318_
timestamp 1644511149
transform 1 0 14168 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1319_
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1320_
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1321_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1322_
timestamp 1644511149
transform 1 0 8372 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1323_
timestamp 1644511149
transform 1 0 9108 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1324_
timestamp 1644511149
transform 1 0 13984 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1325_
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1326_
timestamp 1644511149
transform 1 0 9292 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1327_
timestamp 1644511149
transform 1 0 9108 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1328_
timestamp 1644511149
transform 1 0 13432 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1329_
timestamp 1644511149
transform 1 0 17848 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1330_
timestamp 1644511149
transform 1 0 18032 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1331_
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1332_
timestamp 1644511149
transform 1 0 13616 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1333_
timestamp 1644511149
transform 1 0 19412 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1334_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1335_
timestamp 1644511149
transform 1 0 19964 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1336_
timestamp 1644511149
transform 1 0 20792 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1337_
timestamp 1644511149
transform 1 0 29256 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1338_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1339_
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1340_
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1341_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1342_
timestamp 1644511149
transform 1 0 22264 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1343_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1344_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1345_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1346_
timestamp 1644511149
transform 1 0 46276 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1347_
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1348_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1349_
timestamp 1644511149
transform 1 0 41400 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1350_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1351_
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1352_
timestamp 1644511149
transform 1 0 42688 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1353_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1354_
timestamp 1644511149
transform 1 0 13524 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1355_
timestamp 1644511149
transform 1 0 5888 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1356_
timestamp 1644511149
transform 1 0 2024 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1357_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1358_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1359_
timestamp 1644511149
transform 1 0 46276 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1360_
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1361_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1362_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1363_
timestamp 1644511149
transform 1 0 13800 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1364_
timestamp 1644511149
transform 1 0 46276 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1365_
timestamp 1644511149
transform 1 0 2024 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1366_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1367_
timestamp 1644511149
transform 1 0 1932 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1368_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1369_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1370_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1371_
timestamp 1644511149
transform 1 0 44436 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 27876 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 25300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 24472 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 31372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1644511149
transform 1 0 47656 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 47932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1644511149
transform 1 0 18216 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1644511149
transform 1 0 47288 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input18
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 46092 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 39008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1644511149
transform 1 0 47840 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 47656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1644511149
transform 1 0 47840 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 1644511149
transform 1 0 46736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1644511149
transform 1 0 46184 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 47656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1644511149
transform 1 0 47288 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1644511149
transform 1 0 20056 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 14444 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 24472 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform 1 0 31004 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1644511149
transform 1 0 43148 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 46000 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input66
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 45632 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 47840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1644511149
transform 1 0 46736 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 23368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40296 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 40756 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 39376 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 40204 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 40020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 39560 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 40112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 17940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 17020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 18032 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 17296 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 19596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 20792 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 22080 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 22724 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[0\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31648 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 25024 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 1932 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45540 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  instrumented_adder.tristate_ext_inputs\[4\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34592 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 30084 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 25024 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2576 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45172 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35144 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 45908 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42688 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37352 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 30268 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 30176 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 46184 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 40848 0 1 22848
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
