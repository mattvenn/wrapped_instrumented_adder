magic
tech sky130A
magscale 1 2
timestamp 1654176699
<< viali >>
rect 28457 47209 28491 47243
rect 19441 47141 19475 47175
rect 47961 47141 47995 47175
rect 12357 47073 12391 47107
rect 14105 47073 14139 47107
rect 20085 47073 20119 47107
rect 30757 47073 30791 47107
rect 44465 47073 44499 47107
rect 47041 47073 47075 47107
rect 1961 47005 1995 47039
rect 2697 47005 2731 47039
rect 3801 47005 3835 47039
rect 4813 47005 4847 47039
rect 6837 47005 6871 47039
rect 7757 47005 7791 47039
rect 9413 47005 9447 47039
rect 12633 47005 12667 47039
rect 14381 47005 14415 47039
rect 16681 47005 16715 47039
rect 16957 47005 16991 47039
rect 19257 47005 19291 47039
rect 20361 47005 20395 47039
rect 28641 47005 28675 47039
rect 29745 47005 29779 47039
rect 31033 47005 31067 47039
rect 38393 47005 38427 47039
rect 42625 47005 42659 47039
rect 45201 47005 45235 47039
rect 47777 47005 47811 47039
rect 4077 46937 4111 46971
rect 5181 46937 5215 46971
rect 7941 46937 7975 46971
rect 9597 46937 9631 46971
rect 40325 46937 40359 46971
rect 40509 46937 40543 46971
rect 42809 46937 42843 46971
rect 45385 46937 45419 46971
rect 2145 46869 2179 46903
rect 2881 46869 2915 46903
rect 6929 46869 6963 46903
rect 29929 46869 29963 46903
rect 29469 46597 29503 46631
rect 1409 46529 1443 46563
rect 11713 46529 11747 46563
rect 29285 46529 29319 46563
rect 38117 46529 38151 46563
rect 47869 46529 47903 46563
rect 3985 46461 4019 46495
rect 4169 46461 4203 46495
rect 5089 46461 5123 46495
rect 11989 46461 12023 46495
rect 13185 46461 13219 46495
rect 13645 46461 13679 46495
rect 13829 46461 13863 46495
rect 14289 46461 14323 46495
rect 19441 46461 19475 46495
rect 19625 46461 19659 46495
rect 20637 46461 20671 46495
rect 26157 46461 26191 46495
rect 26985 46461 27019 46495
rect 27169 46461 27203 46495
rect 27721 46461 27755 46495
rect 31125 46461 31159 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 41889 46461 41923 46495
rect 42441 46461 42475 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46857 46461 46891 46495
rect 1593 46325 1627 46359
rect 2329 46325 2363 46359
rect 10793 46325 10827 46359
rect 25513 46325 25547 46359
rect 32321 46325 32355 46359
rect 41245 46325 41279 46359
rect 48053 46325 48087 46359
rect 4353 46121 4387 46155
rect 4997 46121 5031 46155
rect 14197 46121 14231 46155
rect 19349 46121 19383 46155
rect 20085 46121 20119 46155
rect 27629 46121 27663 46155
rect 38393 46121 38427 46155
rect 1409 45985 1443 46019
rect 2789 45985 2823 46019
rect 10609 45985 10643 46019
rect 11069 45985 11103 46019
rect 21373 45985 21407 46019
rect 25237 45985 25271 46019
rect 25697 45985 25731 46019
rect 31677 45985 31711 46019
rect 32229 45985 32263 46019
rect 41337 45985 41371 46019
rect 41889 45985 41923 46019
rect 47041 45985 47075 46019
rect 4905 45917 4939 45951
rect 13093 45917 13127 45951
rect 14105 45917 14139 45951
rect 19257 45917 19291 45951
rect 20913 45917 20947 45951
rect 27537 45917 27571 45951
rect 38301 45917 38335 45951
rect 43913 45917 43947 45951
rect 45661 45917 45695 45951
rect 46305 45917 46339 45951
rect 1593 45849 1627 45883
rect 10793 45849 10827 45883
rect 13461 45849 13495 45883
rect 21097 45849 21131 45883
rect 25421 45849 25455 45883
rect 31861 45849 31895 45883
rect 41521 45849 41555 45883
rect 46489 45849 46523 45883
rect 44097 45781 44131 45815
rect 45753 45781 45787 45815
rect 2237 45577 2271 45611
rect 10793 45577 10827 45611
rect 32229 45577 32263 45611
rect 41797 45577 41831 45611
rect 45937 45577 45971 45611
rect 41153 45509 41187 45543
rect 46581 45509 46615 45543
rect 2145 45441 2179 45475
rect 10701 45441 10735 45475
rect 21097 45441 21131 45475
rect 32137 45441 32171 45475
rect 41061 45441 41095 45475
rect 41705 45441 41739 45475
rect 45293 45441 45327 45475
rect 45845 45441 45879 45475
rect 47593 45441 47627 45475
rect 42625 45373 42659 45407
rect 42809 45373 42843 45407
rect 43177 45373 43211 45407
rect 45109 45237 45143 45271
rect 46673 45237 46707 45271
rect 47685 45237 47719 45271
rect 21189 45033 21223 45067
rect 42625 45033 42659 45067
rect 43269 45033 43303 45067
rect 44465 45033 44499 45067
rect 46489 44897 46523 44931
rect 48145 44897 48179 44931
rect 21097 44829 21131 44863
rect 24777 44829 24811 44863
rect 42533 44829 42567 44863
rect 43177 44829 43211 44863
rect 45477 44829 45511 44863
rect 46305 44829 46339 44863
rect 45661 44761 45695 44795
rect 24869 44693 24903 44727
rect 45293 44489 45327 44523
rect 46949 44489 46983 44523
rect 24685 44421 24719 44455
rect 23765 44353 23799 44387
rect 42901 44353 42935 44387
rect 45201 44353 45235 44387
rect 46397 44353 46431 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 24501 44285 24535 44319
rect 24961 44285 24995 44319
rect 44097 44285 44131 44319
rect 23857 44149 23891 44183
rect 47685 44149 47719 44183
rect 24593 43809 24627 43843
rect 26249 43809 26283 43843
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 23673 43741 23707 43775
rect 23765 43741 23799 43775
rect 24409 43741 24443 43775
rect 45845 43741 45879 43775
rect 46305 43741 46339 43775
rect 1869 43265 1903 43299
rect 46397 43265 46431 43299
rect 47041 43265 47075 43299
rect 1961 43061 1995 43095
rect 47777 43061 47811 43095
rect 46305 42721 46339 42755
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 47685 42313 47719 42347
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 27629 41633 27663 41667
rect 46305 41633 46339 41667
rect 25789 41565 25823 41599
rect 26433 41565 26467 41599
rect 48145 41565 48179 41599
rect 1593 41497 1627 41531
rect 25881 41497 25915 41531
rect 26617 41497 26651 41531
rect 46489 41497 46523 41531
rect 2145 41225 2179 41259
rect 46949 41225 46983 41259
rect 2053 41089 2087 41123
rect 46857 41089 46891 41123
rect 47777 41089 47811 41123
rect 46305 40613 46339 40647
rect 25605 40545 25639 40579
rect 1409 40477 1443 40511
rect 1685 40477 1719 40511
rect 45937 40477 45971 40511
rect 46121 40477 46155 40511
rect 47685 40477 47719 40511
rect 25789 40409 25823 40443
rect 27445 40409 27479 40443
rect 47961 40137 47995 40171
rect 44833 40001 44867 40035
rect 45477 40001 45511 40035
rect 46765 40001 46799 40035
rect 48145 40001 48179 40035
rect 44741 39933 44775 39967
rect 46857 39797 46891 39831
rect 46305 39457 46339 39491
rect 46489 39457 46523 39491
rect 48145 39457 48179 39491
rect 20177 39049 20211 39083
rect 20545 39049 20579 39083
rect 24593 39049 24627 39083
rect 19533 38913 19567 38947
rect 23949 38913 23983 38947
rect 24961 38913 24995 38947
rect 46857 38913 46891 38947
rect 47777 38913 47811 38947
rect 19901 38845 19935 38879
rect 20637 38845 20671 38879
rect 20821 38845 20855 38879
rect 24317 38845 24351 38879
rect 25053 38845 25087 38879
rect 25145 38845 25179 38879
rect 47961 38777 47995 38811
rect 19349 38709 19383 38743
rect 23765 38709 23799 38743
rect 46949 38709 46983 38743
rect 24961 38505 24995 38539
rect 17785 38369 17819 38403
rect 19257 38369 19291 38403
rect 24501 38369 24535 38403
rect 46489 38369 46523 38403
rect 48145 38369 48179 38403
rect 23213 38301 23247 38335
rect 24593 38301 24627 38335
rect 46305 38301 46339 38335
rect 19533 38233 19567 38267
rect 17141 38165 17175 38199
rect 17509 38165 17543 38199
rect 17601 38165 17635 38199
rect 21005 38165 21039 38199
rect 23305 38165 23339 38199
rect 17601 37961 17635 37995
rect 20269 37961 20303 37995
rect 21189 37961 21223 37995
rect 17969 37893 18003 37927
rect 15945 37825 15979 37859
rect 16865 37825 16899 37859
rect 19349 37825 19383 37859
rect 20177 37825 20211 37859
rect 21005 37825 21039 37859
rect 21833 37825 21867 37859
rect 47593 37825 47627 37859
rect 18061 37757 18095 37791
rect 18245 37757 18279 37791
rect 19441 37757 19475 37791
rect 19717 37757 19751 37791
rect 22937 37757 22971 37791
rect 23213 37757 23247 37791
rect 16681 37689 16715 37723
rect 16037 37621 16071 37655
rect 22017 37621 22051 37655
rect 24685 37621 24719 37655
rect 47041 37621 47075 37655
rect 47685 37621 47719 37655
rect 17325 37417 17359 37451
rect 18245 37417 18279 37451
rect 15853 37281 15887 37315
rect 18061 37281 18095 37315
rect 20361 37281 20395 37315
rect 21557 37281 21591 37315
rect 48145 37281 48179 37315
rect 2053 37213 2087 37247
rect 15577 37213 15611 37247
rect 17969 37213 18003 37247
rect 20545 37213 20579 37247
rect 20729 37213 20763 37247
rect 20821 37213 20855 37247
rect 21281 37213 21315 37247
rect 25513 37213 25547 37247
rect 28549 37213 28583 37247
rect 46305 37213 46339 37247
rect 25789 37145 25823 37179
rect 46489 37145 46523 37179
rect 23029 37077 23063 37111
rect 27261 37077 27295 37111
rect 28641 37077 28675 37111
rect 22017 36873 22051 36907
rect 22661 36873 22695 36907
rect 23305 36873 23339 36907
rect 25789 36873 25823 36907
rect 27077 36873 27111 36907
rect 18337 36805 18371 36839
rect 1777 36737 1811 36771
rect 17417 36737 17451 36771
rect 17693 36737 17727 36771
rect 18153 36737 18187 36771
rect 21833 36737 21867 36771
rect 22569 36737 22603 36771
rect 23857 36737 23891 36771
rect 24041 36737 24075 36771
rect 24777 36737 24811 36771
rect 24961 36737 24995 36771
rect 25973 36737 26007 36771
rect 26985 36737 27019 36771
rect 27905 36737 27939 36771
rect 1961 36669 1995 36703
rect 2789 36669 2823 36703
rect 14381 36669 14415 36703
rect 14657 36669 14691 36703
rect 17601 36669 17635 36703
rect 23581 36669 23615 36703
rect 23765 36669 23799 36703
rect 25145 36669 25179 36703
rect 26249 36669 26283 36703
rect 28181 36669 28215 36703
rect 16129 36601 16163 36635
rect 17233 36533 17267 36567
rect 18521 36533 18555 36567
rect 23673 36533 23707 36567
rect 26157 36533 26191 36567
rect 29653 36533 29687 36567
rect 2237 36329 2271 36363
rect 15209 36329 15243 36363
rect 16497 36329 16531 36363
rect 17509 36329 17543 36363
rect 23305 36329 23339 36363
rect 25329 36329 25363 36363
rect 25973 36329 26007 36363
rect 28457 36329 28491 36363
rect 18613 36261 18647 36295
rect 16037 36193 16071 36227
rect 16129 36193 16163 36227
rect 17417 36193 17451 36227
rect 23121 36193 23155 36227
rect 28089 36193 28123 36227
rect 2145 36125 2179 36159
rect 15117 36125 15151 36159
rect 15761 36125 15795 36159
rect 15933 36123 15967 36157
rect 16313 36125 16347 36159
rect 17141 36125 17175 36159
rect 18429 36125 18463 36159
rect 19257 36125 19291 36159
rect 20085 36125 20119 36159
rect 20269 36125 20303 36159
rect 20361 36125 20395 36159
rect 23581 36125 23615 36159
rect 24593 36125 24627 36159
rect 25237 36125 25271 36159
rect 25421 36125 25455 36159
rect 25881 36125 25915 36159
rect 26065 36125 26099 36159
rect 27721 36125 27755 36159
rect 27905 36125 27939 36159
rect 27997 36125 28031 36159
rect 28273 36125 28307 36159
rect 29561 36125 29595 36159
rect 19349 36057 19383 36091
rect 24409 36057 24443 36091
rect 17693 35989 17727 36023
rect 19901 35989 19935 36023
rect 23489 35989 23523 36023
rect 24777 35989 24811 36023
rect 29653 35989 29687 36023
rect 24133 35785 24167 35819
rect 24685 35785 24719 35819
rect 19349 35717 19383 35751
rect 23765 35717 23799 35751
rect 23981 35717 24015 35751
rect 1593 35649 1627 35683
rect 15301 35649 15335 35683
rect 24593 35649 24627 35683
rect 24777 35649 24811 35683
rect 25789 35649 25823 35683
rect 27629 35649 27663 35683
rect 31217 35649 31251 35683
rect 19073 35581 19107 35615
rect 27905 35581 27939 35615
rect 1409 35445 1443 35479
rect 15393 35445 15427 35479
rect 20821 35445 20855 35479
rect 23949 35445 23983 35479
rect 25881 35445 25915 35479
rect 29377 35445 29411 35479
rect 31309 35445 31343 35479
rect 20545 35241 20579 35275
rect 21005 35241 21039 35275
rect 27905 35241 27939 35275
rect 28365 35241 28399 35275
rect 19809 35173 19843 35207
rect 21741 35173 21775 35207
rect 17969 35105 18003 35139
rect 19349 35105 19383 35139
rect 24685 35105 24719 35139
rect 30205 35105 30239 35139
rect 14197 35037 14231 35071
rect 17785 35037 17819 35071
rect 18061 35037 18095 35071
rect 19441 35037 19475 35071
rect 20729 35037 20763 35071
rect 20821 35037 20855 35071
rect 21097 35037 21131 35071
rect 21557 35037 21591 35071
rect 22385 35037 22419 35071
rect 27813 35037 27847 35071
rect 28181 35037 28215 35071
rect 48145 35037 48179 35071
rect 14473 34969 14507 35003
rect 24961 34969 24995 35003
rect 27169 34969 27203 35003
rect 30481 34969 30515 35003
rect 15945 34901 15979 34935
rect 17601 34901 17635 34935
rect 22477 34901 22511 34935
rect 26433 34901 26467 34935
rect 27261 34901 27295 34935
rect 31953 34901 31987 34935
rect 47961 34901 47995 34935
rect 16129 34697 16163 34731
rect 25789 34697 25823 34731
rect 29285 34697 29319 34731
rect 30941 34697 30975 34731
rect 24409 34629 24443 34663
rect 25329 34629 25363 34663
rect 15393 34561 15427 34595
rect 15577 34561 15611 34595
rect 15669 34561 15703 34595
rect 15945 34561 15979 34595
rect 17417 34561 17451 34595
rect 17693 34561 17727 34595
rect 18429 34561 18463 34595
rect 18705 34561 18739 34595
rect 19349 34561 19383 34595
rect 19533 34561 19567 34595
rect 21833 34561 21867 34595
rect 24685 34561 24719 34595
rect 25605 34561 25639 34595
rect 27629 34561 27663 34595
rect 27813 34561 27847 34595
rect 27905 34561 27939 34595
rect 28181 34561 28215 34595
rect 28365 34561 28399 34595
rect 28825 34561 28859 34595
rect 29101 34561 29135 34595
rect 30113 34561 30147 34595
rect 31125 34561 31159 34595
rect 31401 34561 31435 34595
rect 48145 34561 48179 34595
rect 15761 34493 15795 34527
rect 18521 34493 18555 34527
rect 19717 34493 19751 34527
rect 22109 34493 22143 34527
rect 24593 34493 24627 34527
rect 25421 34493 25455 34527
rect 27997 34493 28031 34527
rect 29009 34493 29043 34527
rect 30021 34493 30055 34527
rect 17969 34425 18003 34459
rect 18889 34425 18923 34459
rect 30481 34425 30515 34459
rect 31309 34425 31343 34459
rect 17785 34357 17819 34391
rect 18429 34357 18463 34391
rect 23581 34357 23615 34391
rect 24685 34357 24719 34391
rect 24869 34357 24903 34391
rect 25329 34357 25363 34391
rect 28825 34357 28859 34391
rect 47961 34357 47995 34391
rect 17325 34153 17359 34187
rect 17601 34153 17635 34187
rect 18245 34153 18279 34187
rect 22017 34153 22051 34187
rect 22661 34153 22695 34187
rect 23765 34153 23799 34187
rect 26157 34153 26191 34187
rect 27537 34153 27571 34187
rect 28549 34153 28583 34187
rect 30297 34153 30331 34187
rect 24961 34085 24995 34119
rect 17325 34017 17359 34051
rect 18245 34017 18279 34051
rect 21649 34017 21683 34051
rect 25881 34017 25915 34051
rect 28917 34017 28951 34051
rect 30757 34017 30791 34051
rect 47133 34017 47167 34051
rect 47409 34017 47443 34051
rect 1593 33949 1627 33983
rect 14197 33949 14231 33983
rect 16405 33949 16439 33983
rect 17141 33949 17175 33983
rect 17417 33949 17451 33983
rect 18061 33949 18095 33983
rect 18337 33949 18371 33983
rect 19257 33949 19291 33983
rect 21281 33949 21315 33983
rect 21465 33949 21499 33983
rect 21557 33949 21591 33983
rect 21833 33949 21867 33983
rect 22569 33949 22603 33983
rect 23581 33949 23615 33983
rect 23857 33949 23891 33983
rect 24590 33949 24624 33983
rect 25053 33949 25087 33983
rect 25973 33949 26007 33983
rect 26893 33949 26927 33983
rect 27077 33949 27111 33983
rect 27721 33949 27755 33983
rect 27813 33949 27847 33983
rect 27997 33949 28031 33983
rect 28089 33949 28123 33983
rect 28733 33949 28767 33983
rect 29009 33949 29043 33983
rect 30481 33949 30515 33983
rect 30573 33949 30607 33983
rect 30849 33949 30883 33983
rect 14473 33881 14507 33915
rect 16497 33881 16531 33915
rect 25513 33881 25547 33915
rect 47225 33881 47259 33915
rect 1409 33813 1443 33847
rect 15945 33813 15979 33847
rect 18521 33813 18555 33847
rect 19441 33813 19475 33847
rect 23397 33813 23431 33847
rect 24409 33813 24443 33847
rect 24593 33813 24627 33847
rect 25329 33813 25363 33847
rect 26985 33813 27019 33847
rect 15669 33609 15703 33643
rect 17693 33609 17727 33643
rect 18981 33609 19015 33643
rect 19901 33609 19935 33643
rect 22385 33609 22419 33643
rect 27261 33609 27295 33643
rect 28733 33609 28767 33643
rect 29561 33609 29595 33643
rect 18613 33541 18647 33575
rect 18813 33541 18847 33575
rect 23857 33541 23891 33575
rect 25053 33541 25087 33575
rect 25789 33541 25823 33575
rect 29377 33541 29411 33575
rect 15853 33473 15887 33507
rect 16037 33473 16071 33507
rect 16129 33473 16163 33507
rect 17325 33473 17359 33507
rect 17509 33473 17543 33507
rect 17785 33473 17819 33507
rect 19809 33473 19843 33507
rect 20729 33473 20763 33507
rect 21833 33473 21867 33507
rect 24133 33473 24167 33507
rect 24869 33473 24903 33507
rect 26985 33473 27019 33507
rect 27077 33473 27111 33507
rect 28365 33473 28399 33507
rect 28549 33473 28583 33507
rect 29193 33473 29227 33507
rect 30021 33473 30055 33507
rect 30205 33473 30239 33507
rect 47869 33473 47903 33507
rect 1409 33405 1443 33439
rect 1685 33405 1719 33439
rect 20453 33405 20487 33439
rect 22109 33405 22143 33439
rect 23949 33405 23983 33439
rect 25973 33405 26007 33439
rect 27261 33405 27295 33439
rect 24317 33337 24351 33371
rect 25237 33337 25271 33371
rect 18797 33269 18831 33303
rect 22201 33269 22235 33303
rect 24133 33269 24167 33303
rect 28549 33269 28583 33303
rect 30113 33269 30147 33303
rect 48053 33269 48087 33303
rect 16957 33065 16991 33099
rect 17969 33065 18003 33099
rect 23397 33065 23431 33099
rect 26709 33065 26743 33099
rect 27905 33065 27939 33099
rect 1409 32929 1443 32963
rect 1593 32929 1627 32963
rect 27169 32929 27203 32963
rect 30573 32929 30607 32963
rect 16405 32861 16439 32895
rect 16681 32861 16715 32895
rect 16773 32861 16807 32895
rect 17969 32861 18003 32895
rect 18153 32861 18187 32895
rect 20729 32861 20763 32895
rect 22661 32861 22695 32895
rect 23581 32861 23615 32895
rect 23857 32861 23891 32895
rect 26893 32861 26927 32895
rect 26985 32861 27019 32895
rect 27261 32861 27295 32895
rect 29561 32861 29595 32895
rect 29745 32861 29779 32895
rect 46305 32861 46339 32895
rect 3249 32793 3283 32827
rect 16589 32793 16623 32827
rect 19717 32793 19751 32827
rect 27813 32793 27847 32827
rect 30849 32793 30883 32827
rect 46489 32793 46523 32827
rect 48145 32793 48179 32827
rect 19809 32725 19843 32759
rect 20821 32725 20855 32759
rect 22753 32725 22787 32759
rect 23765 32725 23799 32759
rect 29745 32725 29779 32759
rect 32321 32725 32355 32759
rect 23413 32521 23447 32555
rect 24317 32521 24351 32555
rect 30573 32521 30607 32555
rect 31401 32521 31435 32555
rect 47685 32521 47719 32555
rect 2513 32453 2547 32487
rect 22109 32453 22143 32487
rect 23213 32453 23247 32487
rect 26065 32453 26099 32487
rect 26433 32453 26467 32487
rect 30297 32453 30331 32487
rect 15393 32385 15427 32419
rect 17141 32385 17175 32419
rect 17785 32385 17819 32419
rect 17969 32385 18003 32419
rect 20453 32385 20487 32419
rect 20545 32385 20579 32419
rect 20913 32385 20947 32419
rect 21927 32385 21961 32419
rect 22569 32385 22603 32419
rect 24225 32385 24259 32419
rect 24961 32385 24995 32419
rect 28089 32385 28123 32419
rect 29929 32385 29963 32419
rect 30022 32385 30056 32419
rect 30205 32385 30239 32419
rect 30394 32385 30428 32419
rect 31309 32385 31343 32419
rect 47041 32385 47075 32419
rect 47593 32385 47627 32419
rect 2329 32317 2363 32351
rect 3985 32317 4019 32351
rect 20637 32317 20671 32351
rect 20729 32317 20763 32351
rect 1869 32181 1903 32215
rect 15485 32181 15519 32215
rect 17233 32181 17267 32215
rect 17785 32181 17819 32215
rect 20269 32181 20303 32215
rect 22661 32181 22695 32215
rect 23397 32181 23431 32215
rect 23581 32181 23615 32215
rect 25145 32181 25179 32215
rect 28181 32181 28215 32215
rect 16037 31977 16071 32011
rect 17969 31977 18003 32011
rect 18613 31977 18647 32011
rect 21373 31977 21407 32011
rect 27353 31977 27387 32011
rect 30021 31977 30055 32011
rect 16865 31909 16899 31943
rect 17417 31909 17451 31943
rect 25697 31909 25731 31943
rect 1409 31841 1443 31875
rect 1869 31841 1903 31875
rect 14289 31841 14323 31875
rect 14565 31841 14599 31875
rect 16773 31841 16807 31875
rect 16957 31841 16991 31875
rect 18061 31841 18095 31875
rect 19901 31841 19935 31875
rect 21833 31841 21867 31875
rect 23581 31841 23615 31875
rect 47593 31841 47627 31875
rect 16681 31773 16715 31807
rect 17598 31773 17632 31807
rect 18521 31773 18555 31807
rect 18705 31773 18739 31807
rect 19625 31773 19659 31807
rect 22017 31773 22051 31807
rect 22201 31773 22235 31807
rect 22293 31773 22327 31807
rect 23489 31773 23523 31807
rect 24409 31773 24443 31807
rect 24593 31773 24627 31807
rect 24961 31773 24995 31807
rect 25513 31773 25547 31807
rect 26249 31773 26283 31807
rect 27261 31773 27295 31807
rect 28089 31773 28123 31807
rect 28181 31773 28215 31807
rect 28365 31773 28399 31807
rect 28457 31773 28491 31807
rect 29653 31773 29687 31807
rect 29837 31773 29871 31807
rect 47317 31773 47351 31807
rect 1593 31705 1627 31739
rect 17601 31637 17635 31671
rect 24593 31637 24627 31671
rect 26433 31637 26467 31671
rect 27905 31637 27939 31671
rect 2237 31433 2271 31467
rect 19349 31433 19383 31467
rect 21281 31433 21315 31467
rect 20913 31365 20947 31399
rect 22109 31365 22143 31399
rect 28365 31365 28399 31399
rect 30113 31365 30147 31399
rect 2145 31297 2179 31331
rect 16865 31297 16899 31331
rect 16957 31297 16991 31331
rect 17233 31297 17267 31331
rect 17969 31297 18003 31331
rect 19165 31297 19199 31331
rect 20637 31297 20671 31331
rect 20730 31297 20764 31331
rect 21005 31297 21039 31331
rect 21102 31297 21136 31331
rect 24041 31297 24075 31331
rect 27353 31297 27387 31331
rect 28089 31297 28123 31331
rect 28825 31297 28859 31331
rect 29009 31297 29043 31331
rect 29101 31297 29135 31331
rect 29929 31297 29963 31331
rect 30205 31297 30239 31331
rect 30297 31297 30331 31331
rect 14381 31229 14415 31263
rect 14657 31229 14691 31263
rect 16681 31229 16715 31263
rect 17785 31229 17819 31263
rect 18061 31229 18095 31263
rect 18153 31229 18187 31263
rect 18245 31229 18279 31263
rect 21833 31229 21867 31263
rect 25789 31229 25823 31263
rect 27629 31229 27663 31263
rect 28365 31229 28399 31263
rect 16129 31161 16163 31195
rect 28825 31161 28859 31195
rect 17141 31093 17175 31127
rect 23581 31093 23615 31127
rect 27169 31093 27203 31127
rect 27537 31093 27571 31127
rect 28181 31093 28215 31127
rect 30481 31093 30515 31127
rect 15577 30889 15611 30923
rect 17877 30889 17911 30923
rect 22753 30889 22787 30923
rect 28181 30889 28215 30923
rect 28825 30889 28859 30923
rect 21741 30821 21775 30855
rect 21833 30821 21867 30855
rect 23857 30821 23891 30855
rect 20821 30753 20855 30787
rect 25237 30753 25271 30787
rect 26433 30753 26467 30787
rect 30205 30753 30239 30787
rect 15485 30685 15519 30719
rect 16865 30685 16899 30719
rect 17049 30685 17083 30719
rect 17233 30685 17267 30719
rect 18061 30685 18095 30719
rect 18245 30685 18279 30719
rect 18337 30685 18371 30719
rect 21005 30685 21039 30719
rect 21281 30685 21315 30719
rect 21741 30685 21775 30719
rect 22661 30685 22695 30719
rect 23673 30685 23707 30719
rect 24961 30685 24995 30719
rect 28641 30685 28675 30719
rect 28733 30685 28767 30719
rect 17141 30617 17175 30651
rect 22017 30617 22051 30651
rect 26709 30617 26743 30651
rect 30481 30617 30515 30651
rect 17417 30549 17451 30583
rect 21189 30549 21223 30583
rect 29009 30549 29043 30583
rect 31953 30549 31987 30583
rect 24593 30345 24627 30379
rect 30849 30345 30883 30379
rect 19717 30277 19751 30311
rect 20545 30277 20579 30311
rect 22201 30277 22235 30311
rect 27077 30277 27111 30311
rect 27261 30277 27295 30311
rect 27721 30277 27755 30311
rect 29101 30277 29135 30311
rect 31217 30277 31251 30311
rect 20361 30209 20395 30243
rect 21833 30209 21867 30243
rect 22017 30209 22051 30243
rect 23765 30209 23799 30243
rect 24777 30209 24811 30243
rect 25421 30209 25455 30243
rect 25697 30209 25731 30243
rect 27905 30209 27939 30243
rect 28917 30209 28951 30243
rect 30021 30209 30055 30243
rect 31033 30209 31067 30243
rect 31309 30209 31343 30243
rect 13001 30141 13035 30175
rect 13185 30141 13219 30175
rect 13553 30141 13587 30175
rect 24409 30141 24443 30175
rect 25605 30141 25639 30175
rect 29285 30141 29319 30175
rect 29929 30141 29963 30175
rect 28089 30073 28123 30107
rect 30389 30073 30423 30107
rect 19809 30005 19843 30039
rect 20729 30005 20763 30039
rect 23857 30005 23891 30039
rect 24961 30005 24995 30039
rect 25697 30005 25731 30039
rect 25881 30005 25915 30039
rect 20913 29801 20947 29835
rect 21557 29801 21591 29835
rect 21925 29801 21959 29835
rect 25513 29801 25547 29835
rect 26157 29801 26191 29835
rect 27077 29801 27111 29835
rect 27721 29801 27755 29835
rect 31125 29801 31159 29835
rect 26433 29733 26467 29767
rect 14197 29597 14231 29631
rect 14841 29597 14875 29631
rect 17325 29597 17359 29631
rect 17601 29597 17635 29631
rect 20545 29597 20579 29631
rect 20821 29597 20855 29631
rect 21741 29597 21775 29631
rect 22017 29597 22051 29631
rect 22477 29597 22511 29631
rect 24409 29597 24443 29631
rect 26065 29597 26099 29631
rect 26157 29597 26191 29631
rect 26985 29597 27019 29631
rect 27629 29597 27663 29631
rect 28457 29597 28491 29631
rect 28641 29597 28675 29631
rect 31033 29597 31067 29631
rect 47317 29597 47351 29631
rect 47593 29597 47627 29631
rect 17509 29529 17543 29563
rect 25421 29529 25455 29563
rect 14289 29461 14323 29495
rect 14933 29461 14967 29495
rect 17141 29461 17175 29495
rect 21097 29461 21131 29495
rect 22569 29461 22603 29495
rect 24593 29461 24627 29495
rect 28549 29461 28583 29495
rect 13461 29257 13495 29291
rect 17601 29257 17635 29291
rect 30389 29257 30423 29291
rect 14289 29189 14323 29223
rect 15945 29189 15979 29223
rect 28641 29189 28675 29223
rect 13369 29121 13403 29155
rect 17233 29121 17267 29155
rect 18061 29121 18095 29155
rect 18245 29121 18279 29155
rect 18337 29121 18371 29155
rect 18613 29121 18647 29155
rect 19441 29121 19475 29155
rect 19625 29121 19659 29155
rect 20545 29121 20579 29155
rect 20729 29121 20763 29155
rect 20821 29121 20855 29155
rect 21097 29121 21131 29155
rect 21833 29121 21867 29155
rect 22017 29121 22051 29155
rect 25329 29121 25363 29155
rect 28181 29121 28215 29155
rect 28549 29121 28583 29155
rect 29101 29121 29135 29155
rect 29285 29121 29319 29155
rect 29377 29121 29411 29155
rect 29653 29121 29687 29155
rect 30297 29121 30331 29155
rect 14105 29053 14139 29087
rect 17141 29053 17175 29087
rect 18429 29053 18463 29087
rect 19717 29053 19751 29087
rect 20913 29053 20947 29087
rect 25605 29053 25639 29087
rect 28457 29053 28491 29087
rect 29469 29053 29503 29087
rect 19257 28985 19291 29019
rect 22201 28985 22235 29019
rect 25881 28985 25915 29019
rect 28273 28985 28307 29019
rect 18797 28917 18831 28951
rect 21281 28917 21315 28951
rect 22017 28917 22051 28951
rect 25421 28917 25455 28951
rect 29837 28917 29871 28951
rect 13001 28713 13035 28747
rect 18153 28713 18187 28747
rect 19349 28713 19383 28747
rect 19809 28713 19843 28747
rect 22661 28713 22695 28747
rect 25421 28713 25455 28747
rect 31677 28645 31711 28679
rect 10517 28577 10551 28611
rect 14105 28577 14139 28611
rect 14289 28577 14323 28611
rect 16405 28577 16439 28611
rect 16681 28577 16715 28611
rect 20913 28577 20947 28611
rect 21189 28577 21223 28611
rect 23581 28577 23615 28611
rect 23765 28577 23799 28611
rect 25881 28577 25915 28611
rect 26801 28577 26835 28611
rect 30205 28577 30239 28611
rect 46489 28577 46523 28611
rect 47869 28577 47903 28611
rect 10425 28509 10459 28543
rect 11253 28509 11287 28543
rect 19257 28509 19291 28543
rect 19625 28509 19659 28543
rect 24409 28509 24443 28543
rect 24777 28509 24811 28543
rect 25605 28509 25639 28543
rect 25789 28509 25823 28543
rect 26433 28509 26467 28543
rect 26617 28509 26651 28543
rect 26709 28509 26743 28543
rect 26985 28509 27019 28543
rect 28181 28509 28215 28543
rect 28365 28509 28399 28543
rect 29929 28509 29963 28543
rect 46305 28509 46339 28543
rect 11529 28441 11563 28475
rect 15945 28441 15979 28475
rect 23489 28441 23523 28475
rect 24593 28441 24627 28475
rect 24685 28441 24719 28475
rect 10793 28373 10827 28407
rect 23121 28373 23155 28407
rect 24961 28373 24995 28407
rect 27169 28373 27203 28407
rect 28549 28373 28583 28407
rect 10885 28169 10919 28203
rect 11621 28169 11655 28203
rect 12541 28169 12575 28203
rect 20913 28169 20947 28203
rect 23121 28169 23155 28203
rect 24869 28169 24903 28203
rect 25881 28169 25915 28203
rect 28733 28169 28767 28203
rect 30941 28169 30975 28203
rect 17785 28101 17819 28135
rect 19717 28101 19751 28135
rect 27261 28101 27295 28135
rect 10793 28033 10827 28067
rect 11529 28033 11563 28067
rect 11713 28033 11747 28067
rect 12449 28033 12483 28067
rect 17509 28033 17543 28067
rect 19901 28033 19935 28067
rect 20085 28033 20119 28067
rect 20545 28033 20579 28067
rect 20637 28033 20671 28067
rect 21833 28033 21867 28067
rect 22937 28033 22971 28067
rect 23213 28033 23247 28067
rect 24501 28033 24535 28067
rect 25421 28033 25455 28067
rect 25697 28033 25731 28067
rect 26985 28033 27019 28067
rect 29193 28033 29227 28067
rect 30849 28033 30883 28067
rect 47593 28033 47627 28067
rect 14289 27965 14323 27999
rect 14473 27965 14507 27999
rect 14749 27965 14783 27999
rect 19257 27965 19291 27999
rect 24593 27965 24627 27999
rect 25605 27965 25639 27999
rect 29285 27965 29319 27999
rect 20545 27829 20579 27863
rect 22017 27829 22051 27863
rect 22753 27829 22787 27863
rect 25421 27829 25455 27863
rect 29193 27829 29227 27863
rect 29561 27829 29595 27863
rect 47041 27829 47075 27863
rect 47685 27829 47719 27863
rect 14841 27625 14875 27659
rect 20545 27625 20579 27659
rect 22372 27625 22406 27659
rect 25973 27625 26007 27659
rect 17509 27557 17543 27591
rect 18521 27557 18555 27591
rect 21005 27557 21039 27591
rect 20637 27489 20671 27523
rect 22109 27489 22143 27523
rect 23857 27489 23891 27523
rect 26985 27489 27019 27523
rect 28641 27489 28675 27523
rect 46305 27489 46339 27523
rect 48145 27489 48179 27523
rect 11161 27421 11195 27455
rect 11345 27421 11379 27455
rect 11989 27421 12023 27455
rect 14105 27421 14139 27455
rect 14749 27421 14783 27455
rect 17417 27421 17451 27455
rect 18429 27421 18463 27455
rect 20821 27421 20855 27455
rect 24777 27421 24811 27455
rect 25145 27421 25179 27455
rect 25605 27421 25639 27455
rect 25881 27421 25915 27455
rect 26709 27421 26743 27455
rect 26801 27421 26835 27455
rect 27445 27421 27479 27455
rect 28273 27399 28307 27433
rect 28445 27423 28479 27457
rect 28549 27421 28583 27455
rect 28825 27421 28859 27455
rect 30205 27421 30239 27455
rect 20545 27353 20579 27387
rect 24961 27353 24995 27387
rect 46489 27353 46523 27387
rect 11253 27285 11287 27319
rect 12081 27285 12115 27319
rect 14197 27285 14231 27319
rect 26157 27285 26191 27319
rect 27629 27285 27663 27319
rect 29009 27285 29043 27319
rect 30297 27285 30331 27319
rect 11989 27081 12023 27115
rect 12173 27081 12207 27115
rect 14657 27081 14691 27115
rect 27997 27081 28031 27115
rect 30849 27081 30883 27115
rect 11897 27013 11931 27047
rect 18245 27013 18279 27047
rect 22293 27013 22327 27047
rect 22477 27013 22511 27047
rect 29377 27013 29411 27047
rect 10517 26945 10551 26979
rect 11805 26945 11839 26979
rect 15761 26945 15795 26979
rect 15945 26945 15979 26979
rect 20269 26945 20303 26979
rect 20453 26945 20487 26979
rect 20729 26945 20763 26979
rect 25697 26945 25731 26979
rect 25881 26945 25915 26979
rect 26249 26945 26283 26979
rect 27905 26945 27939 26979
rect 29101 26945 29135 26979
rect 46121 26945 46155 26979
rect 12909 26877 12943 26911
rect 13185 26877 13219 26911
rect 19993 26877 20027 26911
rect 25973 26877 26007 26911
rect 26065 26877 26099 26911
rect 46397 26877 46431 26911
rect 11621 26809 11655 26843
rect 20361 26809 20395 26843
rect 10517 26741 10551 26775
rect 16129 26741 16163 26775
rect 18337 26741 18371 26775
rect 20545 26741 20579 26775
rect 26433 26741 26467 26775
rect 12265 26537 12299 26571
rect 23673 26537 23707 26571
rect 16221 26469 16255 26503
rect 21741 26469 21775 26503
rect 22477 26469 22511 26503
rect 26249 26469 26283 26503
rect 10517 26401 10551 26435
rect 10793 26401 10827 26435
rect 22661 26401 22695 26435
rect 45477 26401 45511 26435
rect 48053 26401 48087 26435
rect 13185 26333 13219 26367
rect 13277 26333 13311 26367
rect 14105 26333 14139 26367
rect 14289 26333 14323 26367
rect 15577 26333 15611 26367
rect 15761 26333 15795 26367
rect 16497 26333 16531 26367
rect 16957 26333 16991 26367
rect 17141 26333 17175 26367
rect 21557 26333 21591 26367
rect 21649 26333 21683 26367
rect 21833 26333 21867 26367
rect 22385 26333 22419 26367
rect 23581 26333 23615 26367
rect 45109 26333 45143 26367
rect 46213 26333 46247 26367
rect 13001 26265 13035 26299
rect 14197 26265 14231 26299
rect 16221 26265 16255 26299
rect 21373 26265 21407 26299
rect 26065 26265 26099 26299
rect 46397 26265 46431 26299
rect 13369 26197 13403 26231
rect 13553 26197 13587 26231
rect 16405 26197 16439 26231
rect 17049 26197 17083 26231
rect 22661 26197 22695 26231
rect 11805 25993 11839 26027
rect 12817 25993 12851 26027
rect 13829 25993 13863 26027
rect 15945 25993 15979 26027
rect 21281 25993 21315 26027
rect 22293 25993 22327 26027
rect 44741 25993 44775 26027
rect 46765 25993 46799 26027
rect 11621 25925 11655 25959
rect 15853 25925 15887 25959
rect 16129 25925 16163 25959
rect 16957 25925 16991 25959
rect 21097 25925 21131 25959
rect 9505 25857 9539 25891
rect 11529 25857 11563 25891
rect 11897 25857 11931 25891
rect 13001 25857 13035 25891
rect 13185 25857 13219 25891
rect 13737 25857 13771 25891
rect 15761 25857 15795 25891
rect 18889 25857 18923 25891
rect 19809 25857 19843 25891
rect 20269 25857 20303 25891
rect 20913 25857 20947 25891
rect 22201 25857 22235 25891
rect 24501 25857 24535 25891
rect 25513 25857 25547 25891
rect 44649 25857 44683 25891
rect 45293 25857 45327 25891
rect 47593 25857 47627 25891
rect 11713 25789 11747 25823
rect 13277 25789 13311 25823
rect 16681 25789 16715 25823
rect 22385 25789 22419 25823
rect 47777 25789 47811 25823
rect 15577 25721 15611 25755
rect 19073 25721 19107 25755
rect 21833 25721 21867 25755
rect 9505 25653 9539 25687
rect 18429 25653 18463 25687
rect 19625 25653 19659 25687
rect 20361 25653 20395 25687
rect 24593 25653 24627 25687
rect 25605 25653 25639 25687
rect 16589 25449 16623 25483
rect 21005 25449 21039 25483
rect 21649 25449 21683 25483
rect 27077 25449 27111 25483
rect 22661 25381 22695 25415
rect 45845 25381 45879 25415
rect 9413 25313 9447 25347
rect 15577 25313 15611 25347
rect 19257 25313 19291 25347
rect 19533 25313 19567 25347
rect 21833 25313 21867 25347
rect 25329 25313 25363 25347
rect 48145 25313 48179 25347
rect 1409 25245 1443 25279
rect 13369 25245 13403 25279
rect 14105 25245 14139 25279
rect 15761 25245 15795 25279
rect 16405 25245 16439 25279
rect 21557 25245 21591 25279
rect 22017 25245 22051 25279
rect 22937 25245 22971 25279
rect 24593 25245 24627 25279
rect 24869 25245 24903 25279
rect 45661 25245 45695 25279
rect 46305 25245 46339 25279
rect 1685 25177 1719 25211
rect 9689 25177 9723 25211
rect 11437 25177 11471 25211
rect 13553 25177 13587 25211
rect 22661 25177 22695 25211
rect 22845 25177 22879 25211
rect 24777 25177 24811 25211
rect 25605 25177 25639 25211
rect 46489 25177 46523 25211
rect 14197 25109 14231 25143
rect 15945 25109 15979 25143
rect 22201 25109 22235 25143
rect 24409 25109 24443 25143
rect 22385 24905 22419 24939
rect 25237 24905 25271 24939
rect 23765 24837 23799 24871
rect 9873 24769 9907 24803
rect 17693 24769 17727 24803
rect 17785 24769 17819 24803
rect 19165 24769 19199 24803
rect 19993 24769 20027 24803
rect 22201 24769 22235 24803
rect 22477 24769 22511 24803
rect 23489 24769 23523 24803
rect 47593 24769 47627 24803
rect 47685 24769 47719 24803
rect 9965 24701 9999 24735
rect 13093 24701 13127 24735
rect 13369 24701 13403 24735
rect 45201 24701 45235 24735
rect 45385 24701 45419 24735
rect 46857 24701 46891 24735
rect 10241 24633 10275 24667
rect 14841 24565 14875 24599
rect 19349 24565 19383 24599
rect 20085 24565 20119 24599
rect 22017 24565 22051 24599
rect 10517 24361 10551 24395
rect 13185 24361 13219 24395
rect 21373 24361 21407 24395
rect 14105 24293 14139 24327
rect 12817 24225 12851 24259
rect 19625 24225 19659 24259
rect 19901 24225 19935 24259
rect 48145 24225 48179 24259
rect 10425 24157 10459 24191
rect 12081 24157 12115 24191
rect 12909 24157 12943 24191
rect 14105 24157 14139 24191
rect 15025 24157 15059 24191
rect 16037 24157 16071 24191
rect 16405 24157 16439 24191
rect 16497 24157 16531 24191
rect 16957 24157 16991 24191
rect 17969 24157 18003 24191
rect 24409 24157 24443 24191
rect 26525 24157 26559 24191
rect 27261 24157 27295 24191
rect 29561 24157 29595 24191
rect 45845 24157 45879 24191
rect 46305 24157 46339 24191
rect 29745 24089 29779 24123
rect 31401 24089 31435 24123
rect 46489 24089 46523 24123
rect 12173 24021 12207 24055
rect 15209 24021 15243 24055
rect 16313 24021 16347 24055
rect 17141 24021 17175 24055
rect 18061 24021 18095 24055
rect 24593 24021 24627 24055
rect 26709 24021 26743 24055
rect 27353 24021 27387 24055
rect 15945 23817 15979 23851
rect 16129 23817 16163 23851
rect 40785 23817 40819 23851
rect 46949 23817 46983 23851
rect 47685 23817 47719 23851
rect 13001 23749 13035 23783
rect 15853 23749 15887 23783
rect 16957 23749 16991 23783
rect 21005 23749 21039 23783
rect 31585 23749 31619 23783
rect 1869 23681 1903 23715
rect 7481 23681 7515 23715
rect 10333 23681 10367 23715
rect 12081 23681 12115 23715
rect 12817 23681 12851 23715
rect 15761 23681 15795 23715
rect 16681 23681 16715 23715
rect 22109 23681 22143 23715
rect 23121 23681 23155 23715
rect 23673 23681 23707 23715
rect 24685 23681 24719 23715
rect 25513 23681 25547 23715
rect 25697 23681 25731 23715
rect 26157 23681 26191 23715
rect 26341 23681 26375 23715
rect 26433 23681 26467 23715
rect 26985 23681 27019 23715
rect 41153 23681 41187 23715
rect 42441 23681 42475 23715
rect 46857 23681 46891 23715
rect 47593 23681 47627 23715
rect 7665 23613 7699 23647
rect 7941 23613 7975 23647
rect 13829 23613 13863 23647
rect 19165 23613 19199 23647
rect 19349 23613 19383 23647
rect 22201 23613 22235 23647
rect 25605 23613 25639 23647
rect 27261 23613 27295 23647
rect 28733 23613 28767 23647
rect 29745 23613 29779 23647
rect 29929 23613 29963 23647
rect 42717 23613 42751 23647
rect 15577 23545 15611 23579
rect 26157 23545 26191 23579
rect 1961 23477 1995 23511
rect 10333 23477 10367 23511
rect 12265 23477 12299 23511
rect 18429 23477 18463 23511
rect 22477 23477 22511 23511
rect 22937 23477 22971 23511
rect 23765 23477 23799 23511
rect 24501 23477 24535 23511
rect 41429 23477 41463 23511
rect 7757 23273 7791 23307
rect 16497 23273 16531 23307
rect 28089 23273 28123 23307
rect 28917 23273 28951 23307
rect 15485 23205 15519 23239
rect 21373 23137 21407 23171
rect 22017 23137 22051 23171
rect 22293 23137 22327 23171
rect 24593 23137 24627 23171
rect 47317 23137 47351 23171
rect 7665 23069 7699 23103
rect 8953 23069 8987 23103
rect 9689 23069 9723 23103
rect 9873 23069 9907 23103
rect 10333 23069 10367 23103
rect 12541 23069 12575 23103
rect 13369 23069 13403 23103
rect 14473 23069 14507 23103
rect 15853 23069 15887 23103
rect 16681 23069 16715 23103
rect 16957 23069 16991 23103
rect 18061 23069 18095 23103
rect 19349 23069 19383 23103
rect 20729 23069 20763 23103
rect 27261 23069 27295 23103
rect 28825 23069 28859 23103
rect 47593 23069 47627 23103
rect 9781 23001 9815 23035
rect 10609 23001 10643 23035
rect 12633 23001 12667 23035
rect 15669 23001 15703 23035
rect 18613 23001 18647 23035
rect 19717 23001 19751 23035
rect 24869 23001 24903 23035
rect 26893 23001 26927 23035
rect 27169 23001 27203 23035
rect 27905 23001 27939 23035
rect 30021 23001 30055 23035
rect 9045 22933 9079 22967
rect 12081 22933 12115 22967
rect 13461 22933 13495 22967
rect 14657 22933 14691 22967
rect 15761 22933 15795 22967
rect 16037 22933 16071 22967
rect 16865 22933 16899 22967
rect 23765 22933 23799 22967
rect 26341 22933 26375 22967
rect 27077 22933 27111 22967
rect 27445 22933 27479 22967
rect 28105 22933 28139 22967
rect 28273 22933 28307 22967
rect 30113 22933 30147 22967
rect 10885 22729 10919 22763
rect 16129 22729 16163 22763
rect 19809 22729 19843 22763
rect 7021 22661 7055 22695
rect 7757 22661 7791 22695
rect 25605 22661 25639 22695
rect 29653 22661 29687 22695
rect 6929 22593 6963 22627
rect 9413 22593 9447 22627
rect 9873 22593 9907 22627
rect 10701 22593 10735 22627
rect 14381 22593 14415 22627
rect 17417 22593 17451 22627
rect 19717 22593 19751 22627
rect 20177 22593 20211 22627
rect 20729 22593 20763 22627
rect 21005 22593 21039 22627
rect 21925 22593 21959 22627
rect 23029 22593 23063 22627
rect 24685 22593 24719 22627
rect 25513 22593 25547 22627
rect 26157 22593 26191 22627
rect 26341 22593 26375 22627
rect 26433 22593 26467 22627
rect 27169 22593 27203 22627
rect 27261 22593 27295 22627
rect 29561 22593 29595 22627
rect 46489 22593 46523 22627
rect 47777 22593 47811 22627
rect 7573 22525 7607 22559
rect 11529 22525 11563 22559
rect 11713 22525 11747 22559
rect 11989 22525 12023 22559
rect 14657 22525 14691 22559
rect 17601 22525 17635 22559
rect 19165 22525 19199 22559
rect 22477 22525 22511 22559
rect 24777 22525 24811 22559
rect 25053 22525 25087 22559
rect 46213 22525 46247 22559
rect 9965 22389 9999 22423
rect 20269 22389 20303 22423
rect 21189 22389 21223 22423
rect 23213 22389 23247 22423
rect 26157 22389 26191 22423
rect 27445 22389 27479 22423
rect 11253 22185 11287 22219
rect 13277 22185 13311 22219
rect 14289 22185 14323 22219
rect 17601 22185 17635 22219
rect 22845 22185 22879 22219
rect 8953 22049 8987 22083
rect 15485 22049 15519 22083
rect 15945 22049 15979 22083
rect 29009 22049 29043 22083
rect 46489 22049 46523 22083
rect 47133 22049 47167 22083
rect 7573 21981 7607 22015
rect 11161 21981 11195 22015
rect 11805 21981 11839 22015
rect 14105 21981 14139 22015
rect 15577 21981 15611 22015
rect 17509 21981 17543 22015
rect 19717 21981 19751 22015
rect 20453 21981 20487 22015
rect 24777 21981 24811 22015
rect 26617 21981 26651 22015
rect 26801 21981 26835 22015
rect 27261 21981 27295 22015
rect 46305 21981 46339 22015
rect 9229 21913 9263 21947
rect 13093 21913 13127 21947
rect 13309 21913 13343 21947
rect 20729 21913 20763 21947
rect 21373 21913 21407 21947
rect 26709 21913 26743 21947
rect 27537 21913 27571 21947
rect 7665 21845 7699 21879
rect 10701 21845 10735 21879
rect 11989 21845 12023 21879
rect 13461 21845 13495 21879
rect 19901 21845 19935 21879
rect 24961 21845 24995 21879
rect 9597 21641 9631 21675
rect 9781 21641 9815 21675
rect 21189 21641 21223 21675
rect 27537 21641 27571 21675
rect 28549 21641 28583 21675
rect 7481 21573 7515 21607
rect 10701 21573 10735 21607
rect 21097 21573 21131 21607
rect 47961 21573 47995 21607
rect 7297 21505 7331 21539
rect 9778 21505 9812 21539
rect 10885 21505 10919 21539
rect 10977 21505 11011 21539
rect 16681 21505 16715 21539
rect 18613 21505 18647 21539
rect 21833 21505 21867 21539
rect 23949 21505 23983 21539
rect 24961 21505 24995 21539
rect 27353 21505 27387 21539
rect 28457 21505 28491 21539
rect 7757 21437 7791 21471
rect 10149 21437 10183 21471
rect 10241 21437 10275 21471
rect 16957 21437 16991 21471
rect 18889 21437 18923 21471
rect 22569 21437 22603 21471
rect 25053 21437 25087 21471
rect 10701 21369 10735 21403
rect 20361 21301 20395 21335
rect 24041 21301 24075 21335
rect 25329 21301 25363 21335
rect 48053 21301 48087 21335
rect 9965 21097 9999 21131
rect 10793 21097 10827 21131
rect 11621 21097 11655 21131
rect 14933 21097 14967 21131
rect 18613 21097 18647 21131
rect 22937 21097 22971 21131
rect 10149 21029 10183 21063
rect 20453 21029 20487 21063
rect 24869 20961 24903 20995
rect 27445 20961 27479 20995
rect 27905 20961 27939 20995
rect 32229 20961 32263 20995
rect 46305 20961 46339 20995
rect 48145 20961 48179 20995
rect 14105 20893 14139 20927
rect 18521 20893 18555 20927
rect 19257 20893 19291 20927
rect 20269 20893 20303 20927
rect 21097 20893 21131 20927
rect 22753 20893 22787 20927
rect 23489 20893 23523 20927
rect 24409 20893 24443 20927
rect 26709 20893 26743 20927
rect 27537 20893 27571 20927
rect 30389 20893 30423 20927
rect 9781 20825 9815 20859
rect 10609 20825 10643 20859
rect 10825 20825 10859 20859
rect 11529 20825 11563 20859
rect 14749 20825 14783 20859
rect 14965 20825 14999 20859
rect 21925 20825 21959 20859
rect 22293 20825 22327 20859
rect 24593 20825 24627 20859
rect 30573 20825 30607 20859
rect 46489 20825 46523 20859
rect 9981 20757 10015 20791
rect 10977 20757 11011 20791
rect 14197 20757 14231 20791
rect 15117 20757 15151 20791
rect 19441 20757 19475 20791
rect 21281 20757 21315 20791
rect 23581 20757 23615 20791
rect 26801 20757 26835 20791
rect 29561 20553 29595 20587
rect 30573 20553 30607 20587
rect 46857 20553 46891 20587
rect 24409 20485 24443 20519
rect 28089 20485 28123 20519
rect 10057 20417 10091 20451
rect 10241 20417 10275 20451
rect 10333 20417 10367 20451
rect 14289 20417 14323 20451
rect 15945 20417 15979 20451
rect 17417 20417 17451 20451
rect 18061 20417 18095 20451
rect 18613 20417 18647 20451
rect 20637 20417 20671 20451
rect 21925 20417 21959 20451
rect 24225 20417 24259 20451
rect 26985 20417 27019 20451
rect 27813 20417 27847 20451
rect 30481 20417 30515 20451
rect 45109 20417 45143 20451
rect 45293 20417 45327 20451
rect 45753 20417 45787 20451
rect 45937 20417 45971 20451
rect 46765 20417 46799 20451
rect 47777 20417 47811 20451
rect 12081 20349 12115 20383
rect 12357 20349 12391 20383
rect 21189 20349 21223 20383
rect 22109 20349 22143 20383
rect 22385 20349 22419 20383
rect 26065 20349 26099 20383
rect 9873 20213 9907 20247
rect 13829 20213 13863 20247
rect 14473 20213 14507 20247
rect 16037 20213 16071 20247
rect 17233 20213 17267 20247
rect 17877 20213 17911 20247
rect 18705 20213 18739 20247
rect 27077 20213 27111 20247
rect 45201 20213 45235 20247
rect 45753 20213 45787 20247
rect 11621 20009 11655 20043
rect 12173 20009 12207 20043
rect 14657 20009 14691 20043
rect 26157 20009 26191 20043
rect 27537 20009 27571 20043
rect 28641 20009 28675 20043
rect 9965 19941 9999 19975
rect 14105 19941 14139 19975
rect 19901 19941 19935 19975
rect 45661 19941 45695 19975
rect 15945 19873 15979 19907
rect 17601 19873 17635 19907
rect 18337 19873 18371 19907
rect 23397 19873 23431 19907
rect 24685 19873 24719 19907
rect 45385 19873 45419 19907
rect 46305 19873 46339 19907
rect 2053 19805 2087 19839
rect 9689 19805 9723 19839
rect 11437 19805 11471 19839
rect 12357 19805 12391 19839
rect 12633 19805 12667 19839
rect 12817 19805 12851 19839
rect 15761 19805 15795 19839
rect 18245 19805 18279 19839
rect 18429 19805 18463 19839
rect 18521 19805 18555 19839
rect 19717 19805 19751 19839
rect 20453 19805 20487 19839
rect 21189 19805 21223 19839
rect 21833 19805 21867 19839
rect 24409 19805 24443 19839
rect 27261 19805 27295 19839
rect 28549 19805 28583 19839
rect 14381 19737 14415 19771
rect 21281 19737 21315 19771
rect 22017 19737 22051 19771
rect 26985 19737 27019 19771
rect 27169 19737 27203 19771
rect 46489 19737 46523 19771
rect 48145 19737 48179 19771
rect 10149 19669 10183 19703
rect 14289 19669 14323 19703
rect 14473 19669 14507 19703
rect 18061 19669 18095 19703
rect 20637 19669 20671 19703
rect 27353 19669 27387 19703
rect 45845 19669 45879 19703
rect 10609 19465 10643 19499
rect 12173 19465 12207 19499
rect 22293 19465 22327 19499
rect 27629 19465 27663 19499
rect 13645 19397 13679 19431
rect 17785 19397 17819 19431
rect 47685 19397 47719 19431
rect 1777 19329 1811 19363
rect 9045 19329 9079 19363
rect 9873 19329 9907 19363
rect 10793 19329 10827 19363
rect 11989 19329 12023 19363
rect 12725 19329 12759 19363
rect 13737 19329 13771 19363
rect 13829 19329 13863 19363
rect 17509 19329 17543 19363
rect 20545 19329 20579 19363
rect 22201 19329 22235 19363
rect 22845 19329 22879 19363
rect 27445 19329 27479 19363
rect 27721 19329 27755 19363
rect 45569 19329 45603 19363
rect 45753 19329 45787 19363
rect 46213 19329 46247 19363
rect 47593 19329 47627 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 9137 19261 9171 19295
rect 14013 19261 14047 19295
rect 23029 19261 23063 19295
rect 23305 19261 23339 19295
rect 13461 19193 13495 19227
rect 46213 19193 46247 19227
rect 9413 19125 9447 19159
rect 10057 19125 10091 19159
rect 12909 19125 12943 19159
rect 19257 19125 19291 19159
rect 20361 19125 20395 19159
rect 27445 19125 27479 19159
rect 2237 18921 2271 18955
rect 18613 18921 18647 18955
rect 19717 18921 19751 18955
rect 22293 18921 22327 18955
rect 22937 18921 22971 18955
rect 24409 18921 24443 18955
rect 27537 18921 27571 18955
rect 18429 18853 18463 18887
rect 9321 18785 9355 18819
rect 11345 18785 11379 18819
rect 11621 18785 11655 18819
rect 14105 18785 14139 18819
rect 17141 18785 17175 18819
rect 25329 18785 25363 18819
rect 25789 18785 25823 18819
rect 47501 18785 47535 18819
rect 2145 18717 2179 18751
rect 9045 18717 9079 18751
rect 16681 18717 16715 18751
rect 17693 18717 17727 18751
rect 18153 18717 18187 18751
rect 19349 18717 19383 18751
rect 19533 18717 19567 18751
rect 20545 18717 20579 18751
rect 22845 18717 22879 18751
rect 23673 18717 23707 18751
rect 24409 18717 24443 18751
rect 25421 18717 25455 18751
rect 26249 18717 26283 18751
rect 28181 18717 28215 18751
rect 28365 18717 28399 18751
rect 45937 18717 45971 18751
rect 46305 18717 46339 18751
rect 14381 18649 14415 18683
rect 17325 18649 17359 18683
rect 20821 18649 20855 18683
rect 27353 18649 27387 18683
rect 10793 18581 10827 18615
rect 13093 18581 13127 18615
rect 15853 18581 15887 18615
rect 16497 18581 16531 18615
rect 17417 18581 17451 18615
rect 17509 18581 17543 18615
rect 23765 18581 23799 18615
rect 26341 18581 26375 18615
rect 27553 18581 27587 18615
rect 27721 18581 27755 18615
rect 28273 18581 28307 18615
rect 9597 18377 9631 18411
rect 10241 18377 10275 18411
rect 11621 18377 11655 18411
rect 14381 18377 14415 18411
rect 16865 18377 16899 18411
rect 18521 18377 18555 18411
rect 20085 18377 20119 18411
rect 22017 18377 22051 18411
rect 22661 18377 22695 18411
rect 47685 18377 47719 18411
rect 2053 18309 2087 18343
rect 17049 18309 17083 18343
rect 18153 18309 18187 18343
rect 24225 18309 24259 18343
rect 27261 18309 27295 18343
rect 1869 18241 1903 18275
rect 9597 18241 9631 18275
rect 10149 18241 10183 18275
rect 11529 18241 11563 18275
rect 13277 18241 13311 18275
rect 14289 18241 14323 18275
rect 15485 18241 15519 18275
rect 16957 18241 16991 18275
rect 18337 18241 18371 18275
rect 19717 18241 19751 18275
rect 20729 18241 20763 18275
rect 21833 18241 21867 18275
rect 22569 18241 22603 18275
rect 23213 18241 23247 18275
rect 46397 18241 46431 18275
rect 47041 18241 47075 18275
rect 47593 18241 47627 18275
rect 13369 18173 13403 18207
rect 13645 18173 13679 18207
rect 15301 18173 15335 18207
rect 17233 18173 17267 18207
rect 19625 18173 19659 18207
rect 24041 18173 24075 18207
rect 24869 18173 24903 18207
rect 26985 18173 27019 18207
rect 16681 18105 16715 18139
rect 15669 18037 15703 18071
rect 20729 18037 20763 18071
rect 23305 18037 23339 18071
rect 28733 18037 28767 18071
rect 46213 18037 46247 18071
rect 14289 17833 14323 17867
rect 16129 17833 16163 17867
rect 19349 17833 19383 17867
rect 26985 17833 27019 17867
rect 28089 17833 28123 17867
rect 14473 17765 14507 17799
rect 16313 17765 16347 17799
rect 16773 17697 16807 17731
rect 20913 17697 20947 17731
rect 25513 17697 25547 17731
rect 12449 17629 12483 17663
rect 13277 17629 13311 17663
rect 13461 17629 13495 17663
rect 17141 17629 17175 17663
rect 18337 17629 18371 17663
rect 19257 17629 19291 17663
rect 19441 17629 19475 17663
rect 25237 17629 25271 17663
rect 27997 17629 28031 17663
rect 45845 17629 45879 17663
rect 46305 17629 46339 17663
rect 14105 17561 14139 17595
rect 14305 17561 14339 17595
rect 15945 17561 15979 17595
rect 17325 17561 17359 17595
rect 21189 17561 21223 17595
rect 22937 17561 22971 17595
rect 29653 17561 29687 17595
rect 29745 17561 29779 17595
rect 30665 17561 30699 17595
rect 46489 17561 46523 17595
rect 48145 17561 48179 17595
rect 12541 17493 12575 17527
rect 13369 17493 13403 17527
rect 16155 17493 16189 17527
rect 16957 17493 16991 17527
rect 17049 17493 17083 17527
rect 18429 17493 18463 17527
rect 25329 17289 25363 17323
rect 25973 17289 26007 17323
rect 47685 17289 47719 17323
rect 13001 17221 13035 17255
rect 15301 17221 15335 17255
rect 23673 17221 23707 17255
rect 28549 17221 28583 17255
rect 29285 17221 29319 17255
rect 45385 17221 45419 17255
rect 47041 17221 47075 17255
rect 12725 17153 12759 17187
rect 15209 17153 15243 17187
rect 15853 17153 15887 17187
rect 17325 17153 17359 17187
rect 18153 17153 18187 17187
rect 23489 17153 23523 17187
rect 23857 17153 23891 17187
rect 24501 17153 24535 17187
rect 25145 17153 25179 17187
rect 25881 17153 25915 17187
rect 28457 17153 28491 17187
rect 29101 17153 29135 17187
rect 47593 17153 47627 17187
rect 14749 17085 14783 17119
rect 17417 17085 17451 17119
rect 18429 17085 18463 17119
rect 24317 17085 24351 17119
rect 30941 17085 30975 17119
rect 45201 17085 45235 17119
rect 17693 17017 17727 17051
rect 2053 16949 2087 16983
rect 15945 16949 15979 16983
rect 19901 16949 19935 16983
rect 24685 16949 24719 16983
rect 14105 16745 14139 16779
rect 1409 16609 1443 16643
rect 1869 16609 1903 16643
rect 11161 16609 11195 16643
rect 15669 16609 15703 16643
rect 15853 16609 15887 16643
rect 21005 16609 21039 16643
rect 25145 16609 25179 16643
rect 30021 16609 30055 16643
rect 31861 16609 31895 16643
rect 39957 16609 39991 16643
rect 40233 16609 40267 16643
rect 46305 16609 46339 16643
rect 10701 16541 10735 16575
rect 14381 16541 14415 16575
rect 19717 16541 19751 16575
rect 23397 16541 23431 16575
rect 23673 16541 23707 16575
rect 24869 16541 24903 16575
rect 1593 16473 1627 16507
rect 10885 16473 10919 16507
rect 14105 16473 14139 16507
rect 17509 16473 17543 16507
rect 21097 16473 21131 16507
rect 22017 16473 22051 16507
rect 23765 16473 23799 16507
rect 30205 16473 30239 16507
rect 40049 16473 40083 16507
rect 46489 16473 46523 16507
rect 48145 16473 48179 16507
rect 14289 16405 14323 16439
rect 19809 16405 19843 16439
rect 2145 16201 2179 16235
rect 10885 16201 10919 16235
rect 17233 16201 17267 16235
rect 19257 16201 19291 16235
rect 30205 16201 30239 16235
rect 47685 16201 47719 16235
rect 17049 16133 17083 16167
rect 2053 16065 2087 16099
rect 10793 16065 10827 16099
rect 15945 16065 15979 16099
rect 16129 16065 16163 16099
rect 17325 16065 17359 16099
rect 18337 16065 18371 16099
rect 19165 16065 19199 16099
rect 23765 16065 23799 16099
rect 24409 16065 24443 16099
rect 30113 16065 30147 16099
rect 47041 16065 47075 16099
rect 47593 16065 47627 16099
rect 17049 15929 17083 15963
rect 15945 15861 15979 15895
rect 18429 15861 18463 15895
rect 23121 15657 23155 15691
rect 24501 15657 24535 15691
rect 10149 15521 10183 15555
rect 13093 15521 13127 15555
rect 13369 15521 13403 15555
rect 15945 15521 15979 15555
rect 20821 15521 20855 15555
rect 21097 15521 21131 15555
rect 23397 15521 23431 15555
rect 47961 15521 47995 15555
rect 2053 15453 2087 15487
rect 9689 15453 9723 15487
rect 13001 15453 13035 15487
rect 14105 15453 14139 15487
rect 14841 15453 14875 15487
rect 18245 15453 18279 15487
rect 20637 15453 20671 15487
rect 23029 15453 23063 15487
rect 23305 15453 23339 15487
rect 24501 15453 24535 15487
rect 24593 15453 24627 15487
rect 46397 15453 46431 15487
rect 47869 15453 47903 15487
rect 48053 15453 48087 15487
rect 9873 15385 9907 15419
rect 16129 15385 16163 15419
rect 17785 15385 17819 15419
rect 47133 15385 47167 15419
rect 14289 15317 14323 15351
rect 14933 15317 14967 15351
rect 18429 15317 18463 15351
rect 23397 15317 23431 15351
rect 10425 15113 10459 15147
rect 16037 15113 16071 15147
rect 18705 15113 18739 15147
rect 22201 15113 22235 15147
rect 23765 15113 23799 15147
rect 23857 15113 23891 15147
rect 24869 15113 24903 15147
rect 13461 15045 13495 15079
rect 17233 15045 17267 15079
rect 23673 15045 23707 15079
rect 47777 15045 47811 15079
rect 1777 14977 1811 15011
rect 10333 14977 10367 15011
rect 15945 14977 15979 15011
rect 16957 14977 16991 15011
rect 20453 14977 20487 15011
rect 21097 14977 21131 15011
rect 22017 14977 22051 15011
rect 22201 14977 22235 15011
rect 22753 14977 22787 15011
rect 22845 14977 22879 15011
rect 24041 14977 24075 15011
rect 24501 14977 24535 15011
rect 24685 14977 24719 15011
rect 45201 14977 45235 15011
rect 47593 14977 47627 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 13185 14909 13219 14943
rect 15209 14909 15243 14943
rect 45385 14909 45419 14943
rect 45753 14909 45787 14943
rect 23489 14841 23523 14875
rect 20545 14773 20579 14807
rect 21189 14773 21223 14807
rect 23029 14773 23063 14807
rect 47961 14773 47995 14807
rect 2237 14569 2271 14603
rect 16221 14569 16255 14603
rect 16405 14569 16439 14603
rect 17049 14569 17083 14603
rect 24501 14569 24535 14603
rect 45661 14569 45695 14603
rect 21833 14433 21867 14467
rect 23305 14433 23339 14467
rect 25145 14433 25179 14467
rect 46673 14433 46707 14467
rect 47225 14433 47259 14467
rect 2145 14365 2179 14399
rect 14105 14365 14139 14399
rect 14933 14365 14967 14399
rect 15209 14365 15243 14399
rect 15393 14365 15427 14399
rect 19349 14365 19383 14399
rect 20269 14365 20303 14399
rect 23029 14365 23063 14399
rect 24409 14365 24443 14399
rect 24593 14365 24627 14399
rect 25053 14365 25087 14399
rect 25237 14365 25271 14399
rect 45569 14365 45603 14399
rect 46489 14365 46523 14399
rect 47777 14365 47811 14399
rect 47961 14365 47995 14399
rect 14197 14297 14231 14331
rect 16037 14297 16071 14331
rect 16865 14297 16899 14331
rect 20453 14297 20487 14331
rect 14749 14229 14783 14263
rect 16247 14229 16281 14263
rect 17065 14229 17099 14263
rect 17233 14229 17267 14263
rect 19441 14229 19475 14263
rect 23857 14229 23891 14263
rect 47869 14229 47903 14263
rect 23765 14025 23799 14059
rect 24409 14025 24443 14059
rect 46397 14025 46431 14059
rect 14013 13957 14047 13991
rect 47685 13957 47719 13991
rect 13185 13889 13219 13923
rect 15945 13889 15979 13923
rect 16773 13889 16807 13923
rect 16957 13889 16991 13923
rect 17601 13889 17635 13923
rect 18429 13889 18463 13923
rect 23673 13889 23707 13923
rect 23857 13889 23891 13923
rect 24317 13889 24351 13923
rect 47041 13889 47075 13923
rect 47593 13889 47627 13923
rect 13277 13821 13311 13855
rect 13737 13821 13771 13855
rect 15485 13821 15519 13855
rect 16865 13821 16899 13855
rect 17509 13821 17543 13855
rect 18705 13821 18739 13855
rect 46765 13821 46799 13855
rect 46857 13821 46891 13855
rect 17969 13753 18003 13787
rect 16037 13685 16071 13719
rect 20177 13685 20211 13719
rect 19441 13481 19475 13515
rect 46673 13481 46707 13515
rect 15301 13345 15335 13379
rect 16129 13345 16163 13379
rect 20545 13345 20579 13379
rect 20729 13345 20763 13379
rect 45845 13345 45879 13379
rect 15117 13277 15151 13311
rect 17601 13277 17635 13311
rect 18429 13277 18463 13311
rect 19441 13277 19475 13311
rect 46029 13277 46063 13311
rect 46673 13277 46707 13311
rect 46857 13277 46891 13311
rect 47685 13277 47719 13311
rect 22385 13209 22419 13243
rect 46213 13209 46247 13243
rect 17601 13141 17635 13175
rect 18521 13141 18555 13175
rect 23489 12869 23523 12903
rect 24225 12869 24259 12903
rect 45293 12869 45327 12903
rect 46213 12869 46247 12903
rect 46857 12869 46891 12903
rect 1409 12801 1443 12835
rect 17141 12801 17175 12835
rect 23397 12801 23431 12835
rect 24041 12801 24075 12835
rect 45201 12801 45235 12835
rect 45385 12801 45419 12835
rect 46029 12801 46063 12835
rect 46305 12801 46339 12835
rect 46765 12801 46799 12835
rect 46949 12801 46983 12835
rect 17417 12733 17451 12767
rect 25881 12733 25915 12767
rect 1593 12597 1627 12631
rect 18889 12597 18923 12631
rect 45845 12597 45879 12631
rect 45385 12393 45419 12427
rect 17049 12325 17083 12359
rect 16773 12257 16807 12291
rect 45753 12257 45787 12291
rect 46305 12257 46339 12291
rect 46489 12257 46523 12291
rect 48145 12257 48179 12291
rect 16681 12189 16715 12223
rect 45569 12189 45603 12223
rect 45845 12189 45879 12223
rect 15117 11713 15151 11747
rect 45753 11713 45787 11747
rect 46213 11713 46247 11747
rect 46397 11577 46431 11611
rect 15209 11509 15243 11543
rect 47777 11509 47811 11543
rect 45845 11305 45879 11339
rect 45661 11237 45695 11271
rect 15025 11169 15059 11203
rect 15209 11169 15243 11203
rect 15485 11169 15519 11203
rect 22201 11169 22235 11203
rect 45385 11169 45419 11203
rect 46305 11169 46339 11203
rect 21741 11101 21775 11135
rect 21925 11033 21959 11067
rect 46489 11033 46523 11067
rect 48145 11033 48179 11067
rect 21925 10761 21959 10795
rect 45385 10761 45419 10795
rect 46121 10693 46155 10727
rect 21833 10625 21867 10659
rect 45293 10625 45327 10659
rect 45477 10625 45511 10659
rect 46029 10557 46063 10591
rect 46305 10557 46339 10591
rect 47777 10421 47811 10455
rect 45661 10217 45695 10251
rect 46305 10081 46339 10115
rect 48145 10081 48179 10115
rect 45569 10013 45603 10047
rect 45753 10013 45787 10047
rect 46489 9945 46523 9979
rect 46857 9673 46891 9707
rect 47685 9605 47719 9639
rect 47041 9537 47075 9571
rect 47593 9537 47627 9571
rect 16313 8993 16347 9027
rect 16773 8993 16807 9027
rect 15669 8925 15703 8959
rect 47317 8925 47351 8959
rect 47593 8925 47627 8959
rect 15761 8857 15795 8891
rect 16497 8857 16531 8891
rect 47777 8517 47811 8551
rect 47961 8313 47995 8347
rect 46305 7905 46339 7939
rect 46489 7905 46523 7939
rect 47685 7905 47719 7939
rect 48145 7361 48179 7395
rect 47961 7157 47995 7191
rect 47133 6817 47167 6851
rect 48145 6817 48179 6851
rect 7573 6749 7607 6783
rect 47225 6681 47259 6715
rect 7665 6613 7699 6647
rect 6929 6341 6963 6375
rect 6745 6205 6779 6239
rect 7205 6205 7239 6239
rect 6929 5865 6963 5899
rect 47317 5729 47351 5763
rect 22201 5661 22235 5695
rect 47593 5661 47627 5695
rect 22293 5525 22327 5559
rect 18889 5185 18923 5219
rect 19901 5185 19935 5219
rect 21833 5185 21867 5219
rect 22477 5185 22511 5219
rect 23489 5185 23523 5219
rect 47041 5185 47075 5219
rect 47869 5185 47903 5219
rect 18981 4981 19015 5015
rect 19993 4981 20027 5015
rect 21925 4981 21959 5015
rect 22569 4981 22603 5015
rect 23305 4981 23339 5015
rect 46857 4981 46891 5015
rect 48053 4981 48087 5015
rect 20821 4777 20855 4811
rect 22753 4777 22787 4811
rect 25237 4641 25271 4675
rect 25421 4641 25455 4675
rect 47133 4641 47167 4675
rect 48145 4641 48179 4675
rect 10609 4573 10643 4607
rect 18521 4573 18555 4607
rect 19441 4573 19475 4607
rect 20085 4573 20119 4607
rect 20729 4573 20763 4607
rect 21373 4573 21407 4607
rect 22017 4573 22051 4607
rect 22661 4573 22695 4607
rect 23305 4573 23339 4607
rect 44097 4573 44131 4607
rect 45937 4573 45971 4607
rect 46397 4573 46431 4607
rect 20177 4505 20211 4539
rect 27077 4505 27111 4539
rect 47225 4505 47259 4539
rect 18613 4437 18647 4471
rect 19533 4437 19567 4471
rect 21465 4437 21499 4471
rect 22109 4437 22143 4471
rect 23397 4437 23431 4471
rect 43913 4437 43947 4471
rect 45753 4437 45787 4471
rect 46489 4437 46523 4471
rect 18153 4233 18187 4267
rect 19533 4233 19567 4267
rect 40601 4233 40635 4267
rect 43729 4165 43763 4199
rect 46581 4165 46615 4199
rect 47777 4165 47811 4199
rect 2053 4097 2087 4131
rect 8769 4097 8803 4131
rect 10149 4097 10183 4131
rect 10425 4097 10459 4131
rect 17417 4097 17451 4131
rect 18061 4097 18095 4131
rect 18797 4097 18831 4131
rect 18889 4097 18923 4131
rect 19441 4097 19475 4131
rect 20637 4097 20671 4131
rect 21833 4097 21867 4131
rect 21925 4097 21959 4131
rect 22477 4097 22511 4131
rect 23213 4097 23247 4131
rect 23857 4097 23891 4131
rect 24685 4097 24719 4131
rect 39865 4097 39899 4131
rect 40509 4097 40543 4131
rect 41153 4097 41187 4131
rect 42901 4097 42935 4131
rect 43545 4097 43579 4131
rect 17509 4029 17543 4063
rect 41337 4029 41371 4063
rect 45109 4029 45143 4063
rect 47961 3961 47995 3995
rect 2145 3893 2179 3927
rect 2881 3893 2915 3927
rect 8861 3893 8895 3927
rect 9597 3893 9631 3927
rect 10517 3893 10551 3927
rect 20729 3893 20763 3927
rect 22569 3893 22603 3927
rect 23305 3893 23339 3927
rect 23949 3893 23983 3927
rect 24777 3893 24811 3927
rect 25513 3893 25547 3927
rect 39957 3893 39991 3927
rect 41521 3893 41555 3927
rect 42993 3893 43027 3927
rect 46029 3893 46063 3927
rect 46673 3893 46707 3927
rect 9689 3689 9723 3723
rect 17693 3689 17727 3723
rect 19441 3689 19475 3723
rect 24869 3689 24903 3723
rect 39221 3689 39255 3723
rect 23305 3621 23339 3655
rect 10333 3553 10367 3587
rect 10517 3553 10551 3587
rect 10977 3553 11011 3587
rect 20177 3553 20211 3587
rect 20453 3553 20487 3587
rect 25421 3553 25455 3587
rect 29561 3553 29595 3587
rect 31401 3553 31435 3587
rect 40049 3553 40083 3587
rect 41521 3553 41555 3587
rect 46305 3553 46339 3587
rect 46489 3553 46523 3587
rect 1409 3485 1443 3519
rect 2145 3485 2179 3519
rect 2973 3485 3007 3519
rect 6653 3485 6687 3519
rect 7481 3485 7515 3519
rect 8217 3485 8251 3519
rect 13553 3485 13587 3519
rect 14105 3485 14139 3519
rect 15301 3485 15335 3519
rect 17601 3485 17635 3519
rect 18245 3485 18279 3519
rect 19349 3485 19383 3519
rect 19993 3485 20027 3519
rect 22753 3485 22787 3519
rect 23213 3485 23247 3519
rect 33057 3485 33091 3519
rect 33885 3485 33919 3519
rect 35909 3485 35943 3519
rect 37749 3485 37783 3519
rect 39129 3485 39163 3519
rect 40325 3485 40359 3519
rect 44005 3485 44039 3519
rect 45201 3485 45235 3519
rect 45661 3485 45695 3519
rect 9413 3417 9447 3451
rect 15485 3417 15519 3451
rect 17141 3417 17175 3451
rect 24777 3417 24811 3451
rect 25605 3417 25639 3451
rect 27261 3417 27295 3451
rect 29745 3417 29779 3451
rect 36093 3417 36127 3451
rect 41705 3417 41739 3451
rect 43361 3417 43395 3451
rect 48145 3417 48179 3451
rect 1593 3349 1627 3383
rect 2237 3349 2271 3383
rect 6745 3349 6779 3383
rect 14197 3349 14231 3383
rect 18337 3349 18371 3383
rect 33149 3349 33183 3383
rect 45753 3349 45787 3383
rect 18245 3145 18279 3179
rect 18889 3145 18923 3179
rect 20821 3145 20855 3179
rect 36185 3145 36219 3179
rect 39129 3145 39163 3179
rect 47869 3145 47903 3179
rect 1961 3077 1995 3111
rect 8125 3077 8159 3111
rect 13737 3077 13771 3111
rect 22753 3077 22787 3111
rect 24961 3077 24995 3111
rect 25053 3077 25087 3111
rect 25973 3077 26007 3111
rect 27629 3077 27663 3111
rect 33149 3077 33183 3111
rect 42901 3077 42935 3111
rect 44557 3077 44591 3111
rect 45385 3077 45419 3111
rect 1777 3009 1811 3043
rect 7941 3009 7975 3043
rect 10241 3009 10275 3043
rect 13553 3009 13587 3043
rect 17325 3009 17359 3043
rect 18153 3009 18187 3043
rect 18797 3009 18831 3043
rect 19441 3009 19475 3043
rect 20269 3009 20303 3043
rect 20729 3009 20763 3043
rect 21925 3009 21959 3043
rect 22569 3009 22603 3043
rect 27445 3009 27479 3043
rect 32965 3009 32999 3043
rect 36369 3009 36403 3043
rect 38485 3009 38519 3043
rect 39589 3009 39623 3043
rect 42717 3009 42751 3043
rect 45201 3009 45235 3043
rect 47777 3009 47811 3043
rect 2237 2941 2271 2975
rect 8401 2941 8435 2975
rect 14197 2941 14231 2975
rect 17233 2941 17267 2975
rect 17693 2941 17727 2975
rect 23029 2941 23063 2975
rect 33517 2941 33551 2975
rect 38669 2941 38703 2975
rect 39773 2941 39807 2975
rect 40049 2941 40083 2975
rect 47041 2941 47075 2975
rect 22109 2873 22143 2907
rect 10333 2805 10367 2839
rect 19533 2805 19567 2839
rect 15577 2601 15611 2635
rect 17969 2601 18003 2635
rect 18613 2601 18647 2635
rect 20913 2601 20947 2635
rect 22017 2601 22051 2635
rect 28641 2601 28675 2635
rect 29745 2601 29779 2635
rect 39221 2601 39255 2635
rect 40417 2601 40451 2635
rect 17325 2533 17359 2567
rect 20177 2533 20211 2567
rect 44373 2533 44407 2567
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2881 2465 2915 2499
rect 5273 2465 5307 2499
rect 6745 2465 6779 2499
rect 7113 2465 7147 2499
rect 9137 2465 9171 2499
rect 9321 2465 9355 2499
rect 10517 2465 10551 2499
rect 24593 2465 24627 2499
rect 24777 2465 24811 2499
rect 25145 2465 25179 2499
rect 35817 2465 35851 2499
rect 41337 2465 41371 2499
rect 42717 2465 42751 2499
rect 45201 2465 45235 2499
rect 45385 2465 45419 2499
rect 45845 2465 45879 2499
rect 3801 2397 3835 2431
rect 4997 2397 5031 2431
rect 6561 2397 6595 2431
rect 15761 2397 15795 2431
rect 17877 2397 17911 2431
rect 18521 2397 18555 2431
rect 20085 2397 20119 2431
rect 22109 2397 22143 2431
rect 22845 2397 22879 2431
rect 26985 2397 27019 2431
rect 27261 2397 27295 2431
rect 29929 2397 29963 2431
rect 35541 2397 35575 2431
rect 38117 2397 38151 2431
rect 39129 2397 39163 2431
rect 41061 2397 41095 2431
rect 42441 2397 42475 2431
rect 44189 2397 44223 2431
rect 17141 2329 17175 2363
rect 20821 2329 20855 2363
rect 28549 2329 28583 2363
rect 40325 2329 40359 2363
rect 47777 2329 47811 2363
rect 3985 2261 4019 2295
rect 38301 2261 38335 2295
rect 47869 2261 47903 2295
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 28445 47243 28503 47249
rect 28445 47209 28457 47243
rect 28491 47240 28503 47243
rect 29270 47240 29276 47252
rect 28491 47212 29276 47240
rect 28491 47209 28503 47212
rect 28445 47203 28503 47209
rect 29270 47200 29276 47212
rect 29328 47200 29334 47252
rect 19429 47175 19487 47181
rect 19429 47141 19441 47175
rect 19475 47172 19487 47175
rect 19978 47172 19984 47184
rect 19475 47144 19984 47172
rect 19475 47141 19487 47144
rect 19429 47135 19487 47141
rect 19978 47132 19984 47144
rect 20036 47132 20042 47184
rect 47949 47175 48007 47181
rect 47949 47172 47961 47175
rect 26206 47144 47961 47172
rect 12250 47064 12256 47116
rect 12308 47104 12314 47116
rect 12345 47107 12403 47113
rect 12345 47104 12357 47107
rect 12308 47076 12357 47104
rect 12308 47064 12314 47076
rect 12345 47073 12357 47076
rect 12391 47073 12403 47107
rect 12345 47067 12403 47073
rect 13814 47064 13820 47116
rect 13872 47104 13878 47116
rect 14093 47107 14151 47113
rect 14093 47104 14105 47107
rect 13872 47076 14105 47104
rect 13872 47064 13878 47076
rect 14093 47073 14105 47076
rect 14139 47073 14151 47107
rect 20070 47104 20076 47116
rect 20031 47076 20076 47104
rect 14093 47067 14151 47073
rect 20070 47064 20076 47076
rect 20128 47064 20134 47116
rect 20530 47064 20536 47116
rect 20588 47104 20594 47116
rect 26206 47104 26234 47144
rect 47949 47141 47961 47144
rect 47995 47141 48007 47175
rect 47949 47135 48007 47141
rect 30742 47104 30748 47116
rect 20588 47076 26234 47104
rect 30703 47076 30748 47104
rect 20588 47064 20594 47076
rect 30742 47064 30748 47076
rect 30800 47064 30806 47116
rect 44453 47107 44511 47113
rect 44453 47073 44465 47107
rect 44499 47104 44511 47107
rect 45094 47104 45100 47116
rect 44499 47076 45100 47104
rect 44499 47073 44511 47076
rect 44453 47067 44511 47073
rect 45094 47064 45100 47076
rect 45152 47064 45158 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 1946 47036 1952 47048
rect 1907 47008 1952 47036
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 2590 46996 2596 47048
rect 2648 47036 2654 47048
rect 2685 47039 2743 47045
rect 2685 47036 2697 47039
rect 2648 47008 2697 47036
rect 2648 46996 2654 47008
rect 2685 47005 2697 47008
rect 2731 47005 2743 47039
rect 2685 46999 2743 47005
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4798 47036 4804 47048
rect 4759 47008 4804 47036
rect 3789 46999 3847 47005
rect 4798 46996 4804 47008
rect 4856 46996 4862 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6825 47039 6883 47045
rect 6825 47036 6837 47039
rect 5868 47008 6837 47036
rect 5868 46996 5874 47008
rect 6825 47005 6837 47008
rect 6871 47005 6883 47039
rect 6825 46999 6883 47005
rect 7098 46996 7104 47048
rect 7156 47036 7162 47048
rect 7745 47039 7803 47045
rect 7745 47036 7757 47039
rect 7156 47008 7757 47036
rect 7156 46996 7162 47008
rect 7745 47005 7757 47008
rect 7791 47005 7803 47039
rect 7745 46999 7803 47005
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 9088 47008 9413 47036
rect 9088 46996 9094 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 12618 47036 12624 47048
rect 12579 47008 12624 47036
rect 9401 46999 9459 47005
rect 12618 46996 12624 47008
rect 12676 46996 12682 47048
rect 14369 47039 14427 47045
rect 14369 47005 14381 47039
rect 14415 47036 14427 47039
rect 14458 47036 14464 47048
rect 14415 47008 14464 47036
rect 14415 47005 14427 47008
rect 14369 46999 14427 47005
rect 14458 46996 14464 47008
rect 14516 46996 14522 47048
rect 16482 46996 16488 47048
rect 16540 47036 16546 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16540 47008 16681 47036
rect 16540 46996 16546 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16669 46999 16727 47005
rect 16945 47039 17003 47045
rect 16945 47005 16957 47039
rect 16991 47005 17003 47039
rect 16945 46999 17003 47005
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 5074 46928 5080 46980
rect 5132 46968 5138 46980
rect 5169 46971 5227 46977
rect 5169 46968 5181 46971
rect 5132 46940 5181 46968
rect 5132 46928 5138 46940
rect 5169 46937 5181 46940
rect 5215 46937 5227 46971
rect 5169 46931 5227 46937
rect 7834 46928 7840 46980
rect 7892 46968 7898 46980
rect 7929 46971 7987 46977
rect 7929 46968 7941 46971
rect 7892 46940 7941 46968
rect 7892 46928 7898 46940
rect 7929 46937 7941 46940
rect 7975 46937 7987 46971
rect 7929 46931 7987 46937
rect 9490 46928 9496 46980
rect 9548 46968 9554 46980
rect 9585 46971 9643 46977
rect 9585 46968 9597 46971
rect 9548 46940 9597 46968
rect 9548 46928 9554 46940
rect 9585 46937 9597 46940
rect 9631 46937 9643 46971
rect 16960 46968 16988 46999
rect 18690 46996 18696 47048
rect 18748 47036 18754 47048
rect 19245 47039 19303 47045
rect 19245 47036 19257 47039
rect 18748 47008 19257 47036
rect 18748 46996 18754 47008
rect 19245 47005 19257 47008
rect 19291 47005 19303 47039
rect 20346 47036 20352 47048
rect 20307 47008 20352 47036
rect 19245 46999 19303 47005
rect 20346 46996 20352 47008
rect 20404 46996 20410 47048
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28629 47039 28687 47045
rect 28629 47036 28641 47039
rect 28408 47008 28641 47036
rect 28408 46996 28414 47008
rect 28629 47005 28641 47008
rect 28675 47005 28687 47039
rect 28629 46999 28687 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 30098 46996 30104 47048
rect 30156 47036 30162 47048
rect 31021 47039 31079 47045
rect 31021 47036 31033 47039
rect 30156 47008 31033 47036
rect 30156 46996 30162 47008
rect 31021 47005 31033 47008
rect 31067 47005 31079 47039
rect 31021 46999 31079 47005
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38381 47039 38439 47045
rect 38381 47036 38393 47039
rect 38160 47008 38393 47036
rect 38160 46996 38166 47008
rect 38381 47005 38393 47008
rect 38427 47005 38439 47039
rect 42610 47036 42616 47048
rect 42571 47008 42616 47036
rect 38381 46999 38439 47005
rect 42610 46996 42616 47008
rect 42668 46996 42674 47048
rect 45186 47036 45192 47048
rect 45147 47008 45192 47036
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47765 47039 47823 47045
rect 47765 47036 47777 47039
rect 47728 47008 47777 47036
rect 47728 46996 47734 47008
rect 47765 47005 47777 47008
rect 47811 47005 47823 47039
rect 47765 46999 47823 47005
rect 20162 46968 20168 46980
rect 16960 46940 20168 46968
rect 9585 46931 9643 46937
rect 20162 46928 20168 46940
rect 20220 46928 20226 46980
rect 40313 46971 40371 46977
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 40313 46931 40371 46937
rect 2130 46900 2136 46912
rect 2091 46872 2136 46900
rect 2130 46860 2136 46872
rect 2188 46860 2194 46912
rect 2866 46900 2872 46912
rect 2827 46872 2872 46900
rect 2866 46860 2872 46872
rect 2924 46860 2930 46912
rect 6914 46860 6920 46912
rect 6972 46900 6978 46912
rect 29914 46900 29920 46912
rect 6972 46872 7017 46900
rect 29875 46872 29920 46900
rect 6972 46860 6978 46872
rect 29914 46860 29920 46872
rect 29972 46860 29978 46912
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 40402 46928 40408 46980
rect 40460 46968 40466 46980
rect 40497 46971 40555 46977
rect 40497 46968 40509 46971
rect 40460 46940 40509 46968
rect 40460 46928 40466 46940
rect 40497 46937 40509 46940
rect 40543 46937 40555 46971
rect 40497 46931 40555 46937
rect 42797 46971 42855 46977
rect 42797 46937 42809 46971
rect 42843 46968 42855 46971
rect 43254 46968 43260 46980
rect 42843 46940 43260 46968
rect 42843 46937 42855 46940
rect 42797 46931 42855 46937
rect 43254 46928 43260 46940
rect 43312 46928 43318 46980
rect 45373 46971 45431 46977
rect 45373 46937 45385 46971
rect 45419 46968 45431 46971
rect 45462 46968 45468 46980
rect 45419 46940 45468 46968
rect 45419 46937 45431 46940
rect 45373 46931 45431 46937
rect 45462 46928 45468 46940
rect 45520 46928 45526 46980
rect 39356 46872 40356 46900
rect 39356 46860 39362 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 2866 46588 2872 46640
rect 2924 46628 2930 46640
rect 29457 46631 29515 46637
rect 29457 46628 29469 46631
rect 2924 46600 29469 46628
rect 2924 46588 2930 46600
rect 29457 46597 29469 46600
rect 29503 46597 29515 46631
rect 29457 46591 29515 46597
rect 1394 46560 1400 46572
rect 1355 46532 1400 46560
rect 1394 46520 1400 46532
rect 1452 46520 1458 46572
rect 11606 46520 11612 46572
rect 11664 46560 11670 46572
rect 11701 46563 11759 46569
rect 11701 46560 11713 46563
rect 11664 46532 11713 46560
rect 11664 46520 11670 46532
rect 11701 46529 11713 46532
rect 11747 46529 11759 46563
rect 29270 46560 29276 46572
rect 29231 46532 29276 46560
rect 11701 46523 11759 46529
rect 29270 46520 29276 46532
rect 29328 46520 29334 46572
rect 38102 46560 38108 46572
rect 38063 46532 38108 46560
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 47854 46560 47860 46572
rect 47815 46532 47860 46560
rect 47854 46520 47860 46532
rect 47912 46520 47918 46572
rect 3970 46492 3976 46504
rect 3931 46464 3976 46492
rect 3970 46452 3976 46464
rect 4028 46452 4034 46504
rect 4157 46495 4215 46501
rect 4157 46461 4169 46495
rect 4203 46492 4215 46495
rect 4982 46492 4988 46504
rect 4203 46464 4988 46492
rect 4203 46461 4215 46464
rect 4157 46455 4215 46461
rect 4982 46452 4988 46464
rect 5040 46452 5046 46504
rect 5077 46495 5135 46501
rect 5077 46461 5089 46495
rect 5123 46461 5135 46495
rect 5077 46455 5135 46461
rect 11977 46495 12035 46501
rect 11977 46461 11989 46495
rect 12023 46461 12035 46495
rect 11977 46455 12035 46461
rect 13173 46495 13231 46501
rect 13173 46461 13185 46495
rect 13219 46492 13231 46495
rect 13633 46495 13691 46501
rect 13633 46492 13645 46495
rect 13219 46464 13645 46492
rect 13219 46461 13231 46464
rect 13173 46455 13231 46461
rect 13633 46461 13645 46464
rect 13679 46461 13691 46495
rect 13633 46455 13691 46461
rect 13817 46495 13875 46501
rect 13817 46461 13829 46495
rect 13863 46492 13875 46495
rect 14182 46492 14188 46504
rect 13863 46464 14188 46492
rect 13863 46461 13875 46464
rect 13817 46455 13875 46461
rect 3878 46384 3884 46436
rect 3936 46424 3942 46436
rect 5092 46424 5120 46455
rect 3936 46396 5120 46424
rect 3936 46384 3942 46396
rect 1581 46359 1639 46365
rect 1581 46325 1593 46359
rect 1627 46356 1639 46359
rect 1670 46356 1676 46368
rect 1627 46328 1676 46356
rect 1627 46325 1639 46328
rect 1581 46319 1639 46325
rect 1670 46316 1676 46328
rect 1728 46316 1734 46368
rect 2314 46356 2320 46368
rect 2275 46328 2320 46356
rect 2314 46316 2320 46328
rect 2372 46316 2378 46368
rect 10594 46316 10600 46368
rect 10652 46356 10658 46368
rect 10781 46359 10839 46365
rect 10781 46356 10793 46359
rect 10652 46328 10793 46356
rect 10652 46316 10658 46328
rect 10781 46325 10793 46328
rect 10827 46325 10839 46359
rect 11992 46356 12020 46455
rect 14182 46452 14188 46464
rect 14240 46452 14246 46504
rect 14274 46452 14280 46504
rect 14332 46492 14338 46504
rect 19429 46495 19487 46501
rect 14332 46464 14377 46492
rect 14332 46452 14338 46464
rect 19429 46461 19441 46495
rect 19475 46461 19487 46495
rect 19610 46492 19616 46504
rect 19571 46464 19616 46492
rect 19429 46455 19487 46461
rect 19444 46424 19472 46455
rect 19610 46452 19616 46464
rect 19668 46452 19674 46504
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 26145 46495 26203 46501
rect 26145 46461 26157 46495
rect 26191 46492 26203 46495
rect 26973 46495 27031 46501
rect 26973 46492 26985 46495
rect 26191 46464 26985 46492
rect 26191 46461 26203 46464
rect 26145 46455 26203 46461
rect 26973 46461 26985 46464
rect 27019 46461 27031 46495
rect 26973 46455 27031 46461
rect 27157 46495 27215 46501
rect 27157 46461 27169 46495
rect 27203 46492 27215 46495
rect 27614 46492 27620 46504
rect 27203 46464 27620 46492
rect 27203 46461 27215 46464
rect 27157 46455 27215 46461
rect 27614 46452 27620 46464
rect 27672 46452 27678 46504
rect 27709 46495 27767 46501
rect 27709 46461 27721 46495
rect 27755 46461 27767 46495
rect 27709 46455 27767 46461
rect 31113 46495 31171 46501
rect 31113 46461 31125 46495
rect 31159 46492 31171 46495
rect 37734 46492 37740 46504
rect 31159 46464 37740 46492
rect 31159 46461 31171 46464
rect 31113 46455 31171 46461
rect 20070 46424 20076 46436
rect 19444 46396 20076 46424
rect 20070 46384 20076 46396
rect 20128 46384 20134 46436
rect 25774 46384 25780 46436
rect 25832 46424 25838 46436
rect 27724 46424 27752 46455
rect 37734 46452 37740 46464
rect 37792 46452 37798 46504
rect 38289 46495 38347 46501
rect 38289 46461 38301 46495
rect 38335 46492 38347 46495
rect 38378 46492 38384 46504
rect 38335 46464 38384 46492
rect 38335 46461 38347 46464
rect 38289 46455 38347 46461
rect 38378 46452 38384 46464
rect 38436 46452 38442 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 41877 46495 41935 46501
rect 41877 46461 41889 46495
rect 41923 46492 41935 46495
rect 42429 46495 42487 46501
rect 42429 46492 42441 46495
rect 41923 46464 42441 46492
rect 41923 46461 41935 46464
rect 41877 46455 41935 46461
rect 42429 46461 42441 46464
rect 42475 46461 42487 46495
rect 42610 46492 42616 46504
rect 42571 46464 42616 46492
rect 42429 46455 42487 46461
rect 42610 46452 42616 46464
rect 42668 46452 42674 46504
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46461 42947 46495
rect 45186 46492 45192 46504
rect 45147 46464 45192 46492
rect 42889 46455 42947 46461
rect 25832 46396 27752 46424
rect 25832 46384 25838 46396
rect 42518 46384 42524 46436
rect 42576 46424 42582 46436
rect 42904 46424 42932 46455
rect 45186 46452 45192 46464
rect 45244 46452 45250 46504
rect 45370 46492 45376 46504
rect 45331 46464 45376 46492
rect 45370 46452 45376 46464
rect 45428 46452 45434 46504
rect 46842 46492 46848 46504
rect 46803 46464 46848 46492
rect 46842 46452 46848 46464
rect 46900 46452 46906 46504
rect 42576 46396 42932 46424
rect 42576 46384 42582 46396
rect 17218 46356 17224 46368
rect 11992 46328 17224 46356
rect 10781 46319 10839 46325
rect 17218 46316 17224 46328
rect 17276 46316 17282 46368
rect 25222 46316 25228 46368
rect 25280 46356 25286 46368
rect 25501 46359 25559 46365
rect 25501 46356 25513 46359
rect 25280 46328 25513 46356
rect 25280 46316 25286 46328
rect 25501 46325 25513 46328
rect 25547 46325 25559 46359
rect 25501 46319 25559 46325
rect 31662 46316 31668 46368
rect 31720 46356 31726 46368
rect 32309 46359 32367 46365
rect 32309 46356 32321 46359
rect 31720 46328 32321 46356
rect 31720 46316 31726 46328
rect 32309 46325 32321 46328
rect 32355 46325 32367 46359
rect 32309 46319 32367 46325
rect 34514 46316 34520 46368
rect 34572 46356 34578 46368
rect 39942 46356 39948 46368
rect 34572 46328 39948 46356
rect 34572 46316 34578 46328
rect 39942 46316 39948 46328
rect 40000 46316 40006 46368
rect 41233 46359 41291 46365
rect 41233 46325 41245 46359
rect 41279 46356 41291 46359
rect 41322 46356 41328 46368
rect 41279 46328 41328 46356
rect 41279 46325 41291 46328
rect 41233 46319 41291 46325
rect 41322 46316 41328 46328
rect 41380 46316 41386 46368
rect 44910 46316 44916 46368
rect 44968 46356 44974 46368
rect 48041 46359 48099 46365
rect 48041 46356 48053 46359
rect 44968 46328 48053 46356
rect 44968 46316 44974 46328
rect 48041 46325 48053 46328
rect 48087 46325 48099 46359
rect 48041 46319 48099 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 3970 46112 3976 46164
rect 4028 46152 4034 46164
rect 4341 46155 4399 46161
rect 4341 46152 4353 46155
rect 4028 46124 4353 46152
rect 4028 46112 4034 46124
rect 4341 46121 4353 46124
rect 4387 46121 4399 46155
rect 4982 46152 4988 46164
rect 4943 46124 4988 46152
rect 4341 46115 4399 46121
rect 4982 46112 4988 46124
rect 5040 46112 5046 46164
rect 14182 46152 14188 46164
rect 14143 46124 14188 46152
rect 14182 46112 14188 46124
rect 14240 46112 14246 46164
rect 19337 46155 19395 46161
rect 19337 46121 19349 46155
rect 19383 46152 19395 46155
rect 19610 46152 19616 46164
rect 19383 46124 19616 46152
rect 19383 46121 19395 46124
rect 19337 46115 19395 46121
rect 19610 46112 19616 46124
rect 19668 46112 19674 46164
rect 20070 46152 20076 46164
rect 20031 46124 20076 46152
rect 20070 46112 20076 46124
rect 20128 46112 20134 46164
rect 27614 46152 27620 46164
rect 27575 46124 27620 46152
rect 27614 46112 27620 46124
rect 27672 46112 27678 46164
rect 38378 46152 38384 46164
rect 38339 46124 38384 46152
rect 38378 46112 38384 46124
rect 38436 46112 38442 46164
rect 38286 46044 38292 46096
rect 38344 46084 38350 46096
rect 44174 46084 44180 46096
rect 38344 46056 44180 46084
rect 38344 46044 38350 46056
rect 44174 46044 44180 46056
rect 44232 46044 44238 46096
rect 1397 46019 1455 46025
rect 1397 45985 1409 46019
rect 1443 46016 1455 46019
rect 2314 46016 2320 46028
rect 1443 45988 2320 46016
rect 1443 45985 1455 45988
rect 1397 45979 1455 45985
rect 2314 45976 2320 45988
rect 2372 45976 2378 46028
rect 2774 46016 2780 46028
rect 2735 45988 2780 46016
rect 2774 45976 2780 45988
rect 2832 45976 2838 46028
rect 10594 46016 10600 46028
rect 10555 45988 10600 46016
rect 10594 45976 10600 45988
rect 10652 45976 10658 46028
rect 10962 45976 10968 46028
rect 11020 46016 11026 46028
rect 11057 46019 11115 46025
rect 11057 46016 11069 46019
rect 11020 45988 11069 46016
rect 11020 45976 11026 45988
rect 11057 45985 11069 45988
rect 11103 45985 11115 46019
rect 11057 45979 11115 45985
rect 21266 45976 21272 46028
rect 21324 46016 21330 46028
rect 21361 46019 21419 46025
rect 21361 46016 21373 46019
rect 21324 45988 21373 46016
rect 21324 45976 21330 45988
rect 21361 45985 21373 45988
rect 21407 45985 21419 46019
rect 25222 46016 25228 46028
rect 25183 45988 25228 46016
rect 21361 45979 21419 45985
rect 25222 45976 25228 45988
rect 25280 45976 25286 46028
rect 25406 45976 25412 46028
rect 25464 46016 25470 46028
rect 25685 46019 25743 46025
rect 25685 46016 25697 46019
rect 25464 45988 25697 46016
rect 25464 45976 25470 45988
rect 25685 45985 25697 45988
rect 25731 45985 25743 46019
rect 25685 45979 25743 45985
rect 27062 45976 27068 46028
rect 27120 46016 27126 46028
rect 27614 46016 27620 46028
rect 27120 45988 27620 46016
rect 27120 45976 27126 45988
rect 27614 45976 27620 45988
rect 27672 45976 27678 46028
rect 31662 46016 31668 46028
rect 31623 45988 31668 46016
rect 31662 45976 31668 45988
rect 31720 45976 31726 46028
rect 32214 46016 32220 46028
rect 32175 45988 32220 46016
rect 32214 45976 32220 45988
rect 32272 45976 32278 46028
rect 41322 46016 41328 46028
rect 41283 45988 41328 46016
rect 41322 45976 41328 45988
rect 41380 45976 41386 46028
rect 41874 46016 41880 46028
rect 41835 45988 41880 46016
rect 41874 45976 41880 45988
rect 41932 45976 41938 46028
rect 47026 46016 47032 46028
rect 46987 45988 47032 46016
rect 47026 45976 47032 45988
rect 47084 45976 47090 46028
rect 4890 45948 4896 45960
rect 4851 45920 4896 45948
rect 4890 45908 4896 45920
rect 4948 45908 4954 45960
rect 12894 45908 12900 45960
rect 12952 45948 12958 45960
rect 13081 45951 13139 45957
rect 13081 45948 13093 45951
rect 12952 45920 13093 45948
rect 12952 45908 12958 45920
rect 13081 45917 13093 45920
rect 13127 45917 13139 45951
rect 14090 45948 14096 45960
rect 14003 45920 14096 45948
rect 13081 45911 13139 45917
rect 14090 45908 14096 45920
rect 14148 45948 14154 45960
rect 18966 45948 18972 45960
rect 14148 45920 18972 45948
rect 14148 45908 14154 45920
rect 18966 45908 18972 45920
rect 19024 45948 19030 45960
rect 19245 45951 19303 45957
rect 19245 45948 19257 45951
rect 19024 45920 19257 45948
rect 19024 45908 19030 45920
rect 19245 45917 19257 45920
rect 19291 45917 19303 45951
rect 20898 45948 20904 45960
rect 20859 45920 20904 45948
rect 19245 45911 19303 45917
rect 20898 45908 20904 45920
rect 20956 45908 20962 45960
rect 27525 45951 27583 45957
rect 27525 45917 27537 45951
rect 27571 45917 27583 45951
rect 38286 45948 38292 45960
rect 38247 45920 38292 45948
rect 27525 45911 27583 45917
rect 1581 45883 1639 45889
rect 1581 45849 1593 45883
rect 1627 45880 1639 45883
rect 2222 45880 2228 45892
rect 1627 45852 2228 45880
rect 1627 45849 1639 45852
rect 1581 45843 1639 45849
rect 2222 45840 2228 45852
rect 2280 45840 2286 45892
rect 10778 45880 10784 45892
rect 10739 45852 10784 45880
rect 10778 45840 10784 45852
rect 10836 45840 10842 45892
rect 13449 45883 13507 45889
rect 13449 45849 13461 45883
rect 13495 45880 13507 45883
rect 21082 45880 21088 45892
rect 13495 45852 16574 45880
rect 21043 45852 21088 45880
rect 13495 45849 13507 45852
rect 13449 45843 13507 45849
rect 16546 45812 16574 45852
rect 21082 45840 21088 45852
rect 21140 45840 21146 45892
rect 25406 45880 25412 45892
rect 25367 45852 25412 45880
rect 25406 45840 25412 45852
rect 25464 45840 25470 45892
rect 20990 45812 20996 45824
rect 16546 45784 20996 45812
rect 20990 45772 20996 45784
rect 21048 45772 21054 45824
rect 27540 45812 27568 45911
rect 38286 45908 38292 45920
rect 38344 45908 38350 45960
rect 43806 45908 43812 45960
rect 43864 45948 43870 45960
rect 43901 45951 43959 45957
rect 43901 45948 43913 45951
rect 43864 45920 43913 45948
rect 43864 45908 43870 45920
rect 43901 45917 43913 45920
rect 43947 45917 43959 45951
rect 43901 45911 43959 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45948 45707 45951
rect 45738 45948 45744 45960
rect 45695 45920 45744 45948
rect 45695 45917 45707 45920
rect 45649 45911 45707 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 46290 45948 46296 45960
rect 46251 45920 46296 45948
rect 46290 45908 46296 45920
rect 46348 45908 46354 45960
rect 31849 45883 31907 45889
rect 31849 45849 31861 45883
rect 31895 45880 31907 45883
rect 32214 45880 32220 45892
rect 31895 45852 32220 45880
rect 31895 45849 31907 45852
rect 31849 45843 31907 45849
rect 32214 45840 32220 45852
rect 32272 45840 32278 45892
rect 41506 45880 41512 45892
rect 41467 45852 41512 45880
rect 41506 45840 41512 45852
rect 41564 45840 41570 45892
rect 46474 45880 46480 45892
rect 46435 45852 46480 45880
rect 46474 45840 46480 45852
rect 46532 45840 46538 45892
rect 41690 45812 41696 45824
rect 27540 45784 41696 45812
rect 41690 45772 41696 45784
rect 41748 45772 41754 45824
rect 43990 45772 43996 45824
rect 44048 45812 44054 45824
rect 44085 45815 44143 45821
rect 44085 45812 44097 45815
rect 44048 45784 44097 45812
rect 44048 45772 44054 45784
rect 44085 45781 44097 45784
rect 44131 45781 44143 45815
rect 45738 45812 45744 45824
rect 45699 45784 45744 45812
rect 44085 45775 44143 45781
rect 45738 45772 45744 45784
rect 45796 45772 45802 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 2222 45608 2228 45620
rect 2183 45580 2228 45608
rect 2222 45568 2228 45580
rect 2280 45568 2286 45620
rect 10778 45608 10784 45620
rect 10739 45580 10784 45608
rect 10778 45568 10784 45580
rect 10836 45568 10842 45620
rect 32214 45608 32220 45620
rect 32175 45580 32220 45608
rect 32214 45568 32220 45580
rect 32272 45568 32278 45620
rect 41785 45611 41843 45617
rect 41785 45577 41797 45611
rect 41831 45608 41843 45611
rect 42610 45608 42616 45620
rect 41831 45580 42616 45608
rect 41831 45577 41843 45580
rect 41785 45571 41843 45577
rect 42610 45568 42616 45580
rect 42668 45568 42674 45620
rect 45925 45611 45983 45617
rect 45925 45577 45937 45611
rect 45971 45608 45983 45611
rect 46474 45608 46480 45620
rect 45971 45580 46480 45608
rect 45971 45577 45983 45580
rect 45925 45571 45983 45577
rect 46474 45568 46480 45580
rect 46532 45568 46538 45620
rect 41141 45543 41199 45549
rect 41141 45509 41153 45543
rect 41187 45540 41199 45543
rect 41506 45540 41512 45552
rect 41187 45512 41512 45540
rect 41187 45509 41199 45512
rect 41141 45503 41199 45509
rect 41506 45500 41512 45512
rect 41564 45500 41570 45552
rect 42628 45512 45968 45540
rect 2133 45475 2191 45481
rect 2133 45441 2145 45475
rect 2179 45472 2191 45475
rect 2406 45472 2412 45484
rect 2179 45444 2412 45472
rect 2179 45441 2191 45444
rect 2133 45435 2191 45441
rect 2406 45432 2412 45444
rect 2464 45472 2470 45484
rect 10689 45475 10747 45481
rect 10689 45472 10701 45475
rect 2464 45444 10701 45472
rect 2464 45432 2470 45444
rect 10689 45441 10701 45444
rect 10735 45441 10747 45475
rect 10689 45435 10747 45441
rect 20898 45432 20904 45484
rect 20956 45472 20962 45484
rect 21085 45475 21143 45481
rect 21085 45472 21097 45475
rect 20956 45444 21097 45472
rect 20956 45432 20962 45444
rect 21085 45441 21097 45444
rect 21131 45441 21143 45475
rect 32122 45472 32128 45484
rect 21085 45435 21143 45441
rect 26206 45444 32128 45472
rect 25774 45364 25780 45416
rect 25832 45404 25838 45416
rect 26206 45404 26234 45444
rect 32122 45432 32128 45444
rect 32180 45432 32186 45484
rect 41046 45432 41052 45484
rect 41104 45472 41110 45484
rect 41690 45472 41696 45484
rect 41104 45444 41149 45472
rect 41603 45444 41696 45472
rect 41104 45432 41110 45444
rect 41690 45432 41696 45444
rect 41748 45472 41754 45484
rect 42628 45472 42656 45512
rect 41748 45444 42656 45472
rect 45281 45475 45339 45481
rect 41748 45432 41754 45444
rect 45281 45441 45293 45475
rect 45327 45441 45339 45475
rect 45830 45472 45836 45484
rect 45791 45444 45836 45472
rect 45281 45435 45339 45441
rect 42426 45404 42432 45416
rect 25832 45376 26234 45404
rect 35866 45376 42432 45404
rect 25832 45364 25838 45376
rect 4890 45296 4896 45348
rect 4948 45336 4954 45348
rect 35866 45336 35894 45376
rect 42426 45364 42432 45376
rect 42484 45364 42490 45416
rect 42610 45404 42616 45416
rect 42571 45376 42616 45404
rect 42610 45364 42616 45376
rect 42668 45364 42674 45416
rect 42794 45404 42800 45416
rect 42755 45376 42800 45404
rect 42794 45364 42800 45376
rect 42852 45364 42858 45416
rect 43162 45404 43168 45416
rect 43123 45376 43168 45404
rect 43162 45364 43168 45376
rect 43220 45364 43226 45416
rect 45296 45404 45324 45435
rect 45830 45432 45836 45444
rect 45888 45432 45894 45484
rect 45940 45472 45968 45512
rect 46382 45500 46388 45552
rect 46440 45540 46446 45552
rect 46569 45543 46627 45549
rect 46569 45540 46581 45543
rect 46440 45512 46581 45540
rect 46440 45500 46446 45512
rect 46569 45509 46581 45512
rect 46615 45509 46627 45543
rect 46569 45503 46627 45509
rect 46474 45472 46480 45484
rect 45940 45444 46480 45472
rect 46474 45432 46480 45444
rect 46532 45432 46538 45484
rect 47302 45432 47308 45484
rect 47360 45472 47366 45484
rect 47581 45475 47639 45481
rect 47581 45472 47593 45475
rect 47360 45444 47593 45472
rect 47360 45432 47366 45444
rect 47581 45441 47593 45444
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 46934 45404 46940 45416
rect 45296 45376 46940 45404
rect 46934 45364 46940 45376
rect 46992 45364 46998 45416
rect 4948 45308 35894 45336
rect 4948 45296 4954 45308
rect 41046 45296 41052 45348
rect 41104 45336 41110 45348
rect 46750 45336 46756 45348
rect 41104 45308 46756 45336
rect 41104 45296 41110 45308
rect 46750 45296 46756 45308
rect 46808 45296 46814 45348
rect 45094 45268 45100 45280
rect 45055 45240 45100 45268
rect 45094 45228 45100 45240
rect 45152 45228 45158 45280
rect 45922 45228 45928 45280
rect 45980 45268 45986 45280
rect 46661 45271 46719 45277
rect 46661 45268 46673 45271
rect 45980 45240 46673 45268
rect 45980 45228 45986 45240
rect 46661 45237 46673 45240
rect 46707 45237 46719 45271
rect 47670 45268 47676 45280
rect 47631 45240 47676 45268
rect 46661 45231 46719 45237
rect 47670 45228 47676 45240
rect 47728 45228 47734 45280
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 21082 45024 21088 45076
rect 21140 45064 21146 45076
rect 21177 45067 21235 45073
rect 21177 45064 21189 45067
rect 21140 45036 21189 45064
rect 21140 45024 21146 45036
rect 21177 45033 21189 45036
rect 21223 45033 21235 45067
rect 21177 45027 21235 45033
rect 42613 45067 42671 45073
rect 42613 45033 42625 45067
rect 42659 45064 42671 45067
rect 42794 45064 42800 45076
rect 42659 45036 42800 45064
rect 42659 45033 42671 45036
rect 42613 45027 42671 45033
rect 42794 45024 42800 45036
rect 42852 45024 42858 45076
rect 43254 45064 43260 45076
rect 43215 45036 43260 45064
rect 43254 45024 43260 45036
rect 43312 45024 43318 45076
rect 44453 45067 44511 45073
rect 44453 45033 44465 45067
rect 44499 45064 44511 45067
rect 45186 45064 45192 45076
rect 44499 45036 45192 45064
rect 44499 45033 44511 45036
rect 44453 45027 44511 45033
rect 45186 45024 45192 45036
rect 45244 45024 45250 45076
rect 45830 45024 45836 45076
rect 45888 45064 45894 45076
rect 47394 45064 47400 45076
rect 45888 45036 47400 45064
rect 45888 45024 45894 45036
rect 47394 45024 47400 45036
rect 47452 45024 47458 45076
rect 25406 44956 25412 45008
rect 25464 44996 25470 45008
rect 45094 44996 45100 45008
rect 25464 44968 45100 44996
rect 25464 44956 25470 44968
rect 45094 44956 45100 44968
rect 45152 44956 45158 45008
rect 42426 44888 42432 44940
rect 42484 44928 42490 44940
rect 45848 44928 45876 45024
rect 42484 44900 45876 44928
rect 46477 44931 46535 44937
rect 42484 44888 42490 44900
rect 46477 44897 46489 44931
rect 46523 44928 46535 44931
rect 47670 44928 47676 44940
rect 46523 44900 47676 44928
rect 46523 44897 46535 44900
rect 46477 44891 46535 44897
rect 47670 44888 47676 44900
rect 47728 44888 47734 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 21085 44863 21143 44869
rect 21085 44829 21097 44863
rect 21131 44860 21143 44863
rect 21818 44860 21824 44872
rect 21131 44832 21824 44860
rect 21131 44829 21143 44832
rect 21085 44823 21143 44829
rect 21818 44820 21824 44832
rect 21876 44820 21882 44872
rect 24765 44863 24823 44869
rect 24765 44829 24777 44863
rect 24811 44860 24823 44863
rect 25774 44860 25780 44872
rect 24811 44832 25780 44860
rect 24811 44829 24823 44832
rect 24765 44823 24823 44829
rect 25774 44820 25780 44832
rect 25832 44820 25838 44872
rect 42521 44863 42579 44869
rect 42521 44829 42533 44863
rect 42567 44829 42579 44863
rect 43162 44860 43168 44872
rect 43123 44832 43168 44860
rect 42521 44823 42579 44829
rect 24670 44684 24676 44736
rect 24728 44724 24734 44736
rect 24857 44727 24915 44733
rect 24857 44724 24869 44727
rect 24728 44696 24869 44724
rect 24728 44684 24734 44696
rect 24857 44693 24869 44696
rect 24903 44693 24915 44727
rect 42536 44724 42564 44823
rect 43162 44820 43168 44832
rect 43220 44820 43226 44872
rect 44450 44820 44456 44872
rect 44508 44860 44514 44872
rect 45465 44863 45523 44869
rect 45465 44860 45477 44863
rect 44508 44832 45477 44860
rect 44508 44820 44514 44832
rect 45465 44829 45477 44832
rect 45511 44829 45523 44863
rect 45465 44823 45523 44829
rect 46293 44863 46351 44869
rect 46293 44829 46305 44863
rect 46339 44829 46351 44863
rect 46293 44823 46351 44829
rect 45649 44795 45707 44801
rect 45649 44761 45661 44795
rect 45695 44792 45707 44795
rect 46014 44792 46020 44804
rect 45695 44764 46020 44792
rect 45695 44761 45707 44764
rect 45649 44755 45707 44761
rect 46014 44752 46020 44764
rect 46072 44752 46078 44804
rect 46308 44792 46336 44823
rect 47026 44792 47032 44804
rect 46308 44764 47032 44792
rect 47026 44752 47032 44764
rect 47084 44752 47090 44804
rect 47578 44724 47584 44736
rect 42536 44696 47584 44724
rect 24857 44687 24915 44693
rect 47578 44684 47584 44696
rect 47636 44684 47642 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 45281 44523 45339 44529
rect 45281 44489 45293 44523
rect 45327 44520 45339 44523
rect 45370 44520 45376 44532
rect 45327 44492 45376 44520
rect 45327 44489 45339 44492
rect 45281 44483 45339 44489
rect 45370 44480 45376 44492
rect 45428 44480 45434 44532
rect 45462 44480 45468 44532
rect 45520 44520 45526 44532
rect 46937 44523 46995 44529
rect 46937 44520 46949 44523
rect 45520 44492 46949 44520
rect 45520 44480 45526 44492
rect 46937 44489 46949 44492
rect 46983 44489 46995 44523
rect 46937 44483 46995 44489
rect 24670 44452 24676 44464
rect 24631 44424 24676 44452
rect 24670 44412 24676 44424
rect 24728 44412 24734 44464
rect 21818 44344 21824 44396
rect 21876 44384 21882 44396
rect 23753 44387 23811 44393
rect 23753 44384 23765 44387
rect 21876 44356 23765 44384
rect 21876 44344 21882 44356
rect 23753 44353 23765 44356
rect 23799 44353 23811 44387
rect 23753 44347 23811 44353
rect 42610 44344 42616 44396
rect 42668 44384 42674 44396
rect 42889 44387 42947 44393
rect 42889 44384 42901 44387
rect 42668 44356 42901 44384
rect 42668 44344 42674 44356
rect 42889 44353 42901 44356
rect 42935 44353 42947 44387
rect 42889 44347 42947 44353
rect 44174 44344 44180 44396
rect 44232 44384 44238 44396
rect 45189 44387 45247 44393
rect 45189 44384 45201 44387
rect 44232 44356 45201 44384
rect 44232 44344 44238 44356
rect 45189 44353 45201 44356
rect 45235 44353 45247 44387
rect 45189 44347 45247 44353
rect 46290 44344 46296 44396
rect 46348 44384 46354 44396
rect 46385 44387 46443 44393
rect 46385 44384 46397 44387
rect 46348 44356 46397 44384
rect 46348 44344 46354 44356
rect 46385 44353 46397 44356
rect 46431 44353 46443 44387
rect 46385 44347 46443 44353
rect 46845 44387 46903 44393
rect 46845 44353 46857 44387
rect 46891 44384 46903 44387
rect 47302 44384 47308 44396
rect 46891 44356 47308 44384
rect 46891 44353 46903 44356
rect 46845 44347 46903 44353
rect 47302 44344 47308 44356
rect 47360 44384 47366 44396
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 47360 44356 47593 44384
rect 47360 44344 47366 44356
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 24486 44316 24492 44328
rect 24447 44288 24492 44316
rect 24486 44276 24492 44288
rect 24544 44276 24550 44328
rect 24949 44319 25007 44325
rect 24949 44285 24961 44319
rect 24995 44285 25007 44319
rect 24949 44279 25007 44285
rect 2958 44208 2964 44260
rect 3016 44248 3022 44260
rect 24964 44248 24992 44279
rect 42702 44276 42708 44328
rect 42760 44316 42766 44328
rect 44085 44319 44143 44325
rect 44085 44316 44097 44319
rect 42760 44288 44097 44316
rect 42760 44276 42766 44288
rect 44085 44285 44097 44288
rect 44131 44285 44143 44319
rect 44085 44279 44143 44285
rect 3016 44220 24992 44248
rect 3016 44208 3022 44220
rect 23845 44183 23903 44189
rect 23845 44149 23857 44183
rect 23891 44180 23903 44183
rect 24578 44180 24584 44192
rect 23891 44152 24584 44180
rect 23891 44149 23903 44152
rect 23845 44143 23903 44149
rect 24578 44140 24584 44152
rect 24636 44140 24642 44192
rect 47670 44180 47676 44192
rect 47631 44152 47676 44180
rect 47670 44140 47676 44152
rect 47728 44140 47734 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 24578 43840 24584 43852
rect 24539 43812 24584 43840
rect 24578 43800 24584 43812
rect 24636 43800 24642 43852
rect 26237 43843 26295 43849
rect 26237 43809 26249 43843
rect 26283 43840 26295 43843
rect 34514 43840 34520 43852
rect 26283 43812 34520 43840
rect 26283 43809 26295 43812
rect 26237 43803 26295 43809
rect 34514 43800 34520 43812
rect 34572 43800 34578 43852
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 47670 43840 47676 43852
rect 46523 43812 47676 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 47670 43800 47676 43812
rect 47728 43800 47734 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 23474 43732 23480 43784
rect 23532 43772 23538 43784
rect 23661 43775 23719 43781
rect 23661 43772 23673 43775
rect 23532 43744 23673 43772
rect 23532 43732 23538 43744
rect 23661 43741 23673 43744
rect 23707 43741 23719 43775
rect 23661 43735 23719 43741
rect 23753 43775 23811 43781
rect 23753 43741 23765 43775
rect 23799 43772 23811 43775
rect 24397 43775 24455 43781
rect 24397 43772 24409 43775
rect 23799 43744 24409 43772
rect 23799 43741 23811 43744
rect 23753 43735 23811 43741
rect 24397 43741 24409 43744
rect 24443 43741 24455 43775
rect 24397 43735 24455 43741
rect 45833 43775 45891 43781
rect 45833 43741 45845 43775
rect 45879 43772 45891 43775
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 45879 43744 46305 43772
rect 45879 43741 45891 43744
rect 45833 43735 45891 43741
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1854 43296 1860 43308
rect 1815 43268 1860 43296
rect 1854 43256 1860 43268
rect 1912 43256 1918 43308
rect 45278 43256 45284 43308
rect 45336 43296 45342 43308
rect 46385 43299 46443 43305
rect 46385 43296 46397 43299
rect 45336 43268 46397 43296
rect 45336 43256 45342 43268
rect 46385 43265 46397 43268
rect 46431 43265 46443 43299
rect 47026 43296 47032 43308
rect 46987 43268 47032 43296
rect 46385 43259 46443 43265
rect 47026 43256 47032 43268
rect 47084 43256 47090 43308
rect 1946 43092 1952 43104
rect 1907 43064 1952 43092
rect 1946 43052 1952 43064
rect 2004 43052 2010 43104
rect 47762 43092 47768 43104
rect 47723 43064 47768 43092
rect 47762 43052 47768 43064
rect 47820 43052 47826 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46293 42755 46351 42761
rect 46293 42721 46305 42755
rect 46339 42752 46351 42755
rect 47762 42752 47768 42764
rect 46339 42724 47768 42752
rect 46339 42721 46351 42724
rect 46293 42715 46351 42721
rect 47762 42712 47768 42724
rect 47820 42712 47826 42764
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 47670 42616 47676 42628
rect 46523 42588 47676 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 47670 42576 47676 42588
rect 47728 42576 47734 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 47670 42344 47676 42356
rect 47631 42316 47676 42344
rect 47670 42304 47676 42316
rect 47728 42304 47734 42356
rect 47118 42168 47124 42220
rect 47176 42208 47182 42220
rect 47578 42208 47584 42220
rect 47176 42180 47584 42208
rect 47176 42168 47182 42180
rect 47578 42168 47584 42180
rect 47636 42168 47642 42220
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 27614 41664 27620 41676
rect 27575 41636 27620 41664
rect 27614 41624 27620 41636
rect 27672 41624 27678 41676
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41664 46351 41667
rect 47762 41664 47768 41676
rect 46339 41636 47768 41664
rect 46339 41633 46351 41636
rect 46293 41627 46351 41633
rect 47762 41624 47768 41636
rect 47820 41624 47826 41676
rect 25774 41596 25780 41608
rect 25735 41568 25780 41596
rect 25774 41556 25780 41568
rect 25832 41556 25838 41608
rect 26418 41596 26424 41608
rect 26379 41568 26424 41596
rect 26418 41556 26424 41568
rect 26476 41556 26482 41608
rect 48130 41596 48136 41608
rect 48091 41568 48136 41596
rect 48130 41556 48136 41568
rect 48188 41556 48194 41608
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 25869 41531 25927 41537
rect 25869 41497 25881 41531
rect 25915 41528 25927 41531
rect 26605 41531 26663 41537
rect 26605 41528 26617 41531
rect 25915 41500 26617 41528
rect 25915 41497 25927 41500
rect 25869 41491 25927 41497
rect 26605 41497 26617 41500
rect 26651 41497 26663 41531
rect 26605 41491 26663 41497
rect 46477 41531 46535 41537
rect 46477 41497 46489 41531
rect 46523 41528 46535 41531
rect 46934 41528 46940 41540
rect 46523 41500 46940 41528
rect 46523 41497 46535 41500
rect 46477 41491 46535 41497
rect 46934 41488 46940 41500
rect 46992 41488 46998 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2133 41259 2191 41265
rect 2133 41256 2145 41259
rect 1636 41228 2145 41256
rect 1636 41216 1642 41228
rect 2133 41225 2145 41228
rect 2179 41225 2191 41259
rect 46934 41256 46940 41268
rect 46895 41228 46940 41256
rect 2133 41219 2191 41225
rect 46934 41216 46940 41228
rect 46992 41216 46998 41268
rect 2041 41123 2099 41129
rect 2041 41089 2053 41123
rect 2087 41120 2099 41123
rect 14090 41120 14096 41132
rect 2087 41092 14096 41120
rect 2087 41089 2099 41092
rect 2041 41083 2099 41089
rect 14090 41080 14096 41092
rect 14148 41080 14154 41132
rect 46566 41080 46572 41132
rect 46624 41120 46630 41132
rect 46845 41123 46903 41129
rect 46845 41120 46857 41123
rect 46624 41092 46857 41120
rect 46624 41080 46630 41092
rect 46845 41089 46857 41092
rect 46891 41089 46903 41123
rect 47762 41120 47768 41132
rect 47723 41092 47768 41120
rect 46845 41083 46903 41089
rect 47762 41080 47768 41092
rect 47820 41080 47826 41132
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 26418 40604 26424 40656
rect 26476 40644 26482 40656
rect 46293 40647 46351 40653
rect 46293 40644 46305 40647
rect 26476 40616 46305 40644
rect 26476 40604 26482 40616
rect 46293 40613 46305 40616
rect 46339 40613 46351 40647
rect 46293 40607 46351 40613
rect 25593 40579 25651 40585
rect 25593 40545 25605 40579
rect 25639 40576 25651 40579
rect 26436 40576 26464 40604
rect 25639 40548 26464 40576
rect 25639 40545 25651 40548
rect 25593 40539 25651 40545
rect 1394 40508 1400 40520
rect 1355 40480 1400 40508
rect 1394 40468 1400 40480
rect 1452 40468 1458 40520
rect 1673 40511 1731 40517
rect 1673 40477 1685 40511
rect 1719 40477 1731 40511
rect 1673 40471 1731 40477
rect 45925 40511 45983 40517
rect 45925 40477 45937 40511
rect 45971 40477 45983 40511
rect 46106 40508 46112 40520
rect 46067 40480 46112 40508
rect 45925 40471 45983 40477
rect 1688 40372 1716 40471
rect 2130 40400 2136 40452
rect 2188 40440 2194 40452
rect 25777 40443 25835 40449
rect 25777 40440 25789 40443
rect 2188 40412 25789 40440
rect 2188 40400 2194 40412
rect 25777 40409 25789 40412
rect 25823 40409 25835 40443
rect 27430 40440 27436 40452
rect 27391 40412 27436 40440
rect 25777 40403 25835 40409
rect 27430 40400 27436 40412
rect 27488 40400 27494 40452
rect 45940 40440 45968 40471
rect 46106 40468 46112 40480
rect 46164 40468 46170 40520
rect 47670 40508 47676 40520
rect 47631 40480 47676 40508
rect 47670 40468 47676 40480
rect 47728 40468 47734 40520
rect 46198 40440 46204 40452
rect 45940 40412 46204 40440
rect 46198 40400 46204 40412
rect 46256 40400 46262 40452
rect 10962 40372 10968 40384
rect 1688 40344 10968 40372
rect 10962 40332 10968 40344
rect 11020 40332 11026 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 47949 40171 48007 40177
rect 47949 40168 47961 40171
rect 45526 40140 47961 40168
rect 45526 40100 45554 40140
rect 47949 40137 47961 40140
rect 47995 40137 48007 40171
rect 47949 40131 48007 40137
rect 44836 40072 45554 40100
rect 44836 40041 44864 40072
rect 48038 40060 48044 40112
rect 48096 40060 48102 40112
rect 44821 40035 44879 40041
rect 44821 40001 44833 40035
rect 44867 40001 44879 40035
rect 44821 39995 44879 40001
rect 45465 40035 45523 40041
rect 45465 40001 45477 40035
rect 45511 40032 45523 40035
rect 46106 40032 46112 40044
rect 45511 40004 46112 40032
rect 45511 40001 45523 40004
rect 45465 39995 45523 40001
rect 46106 39992 46112 40004
rect 46164 39992 46170 40044
rect 46750 40032 46756 40044
rect 46711 40004 46756 40032
rect 46750 39992 46756 40004
rect 46808 39992 46814 40044
rect 48056 40032 48084 40060
rect 48133 40035 48191 40041
rect 48133 40032 48145 40035
rect 48056 40004 48145 40032
rect 48133 40001 48145 40004
rect 48179 40001 48191 40035
rect 48133 39995 48191 40001
rect 44726 39964 44732 39976
rect 44687 39936 44732 39964
rect 44726 39924 44732 39936
rect 44784 39924 44790 39976
rect 46474 39788 46480 39840
rect 46532 39828 46538 39840
rect 46845 39831 46903 39837
rect 46845 39828 46857 39831
rect 46532 39800 46857 39828
rect 46532 39788 46538 39800
rect 46845 39797 46857 39800
rect 46891 39797 46903 39831
rect 46845 39791 46903 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 47670 39556 47676 39568
rect 46308 39528 47676 39556
rect 46308 39497 46336 39528
rect 47670 39516 47676 39528
rect 47728 39516 47734 39568
rect 46293 39491 46351 39497
rect 46293 39457 46305 39491
rect 46339 39457 46351 39491
rect 46474 39488 46480 39500
rect 46435 39460 46480 39488
rect 46293 39451 46351 39457
rect 46474 39448 46480 39460
rect 46532 39448 46538 39500
rect 48133 39491 48191 39497
rect 48133 39457 48145 39491
rect 48179 39488 48191 39491
rect 48222 39488 48228 39500
rect 48179 39460 48228 39488
rect 48179 39457 48191 39460
rect 48133 39451 48191 39457
rect 48222 39448 48228 39460
rect 48280 39448 48286 39500
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 20165 39083 20223 39089
rect 20165 39049 20177 39083
rect 20211 39049 20223 39083
rect 20530 39080 20536 39092
rect 20165 39043 20223 39049
rect 20272 39052 20536 39080
rect 19521 38947 19579 38953
rect 19521 38913 19533 38947
rect 19567 38944 19579 38947
rect 20180 38944 20208 39043
rect 19567 38916 20208 38944
rect 19567 38913 19579 38916
rect 19521 38907 19579 38913
rect 19889 38879 19947 38885
rect 19889 38845 19901 38879
rect 19935 38876 19947 38879
rect 20272 38876 20300 39052
rect 20530 39040 20536 39052
rect 20588 39040 20594 39092
rect 24581 39083 24639 39089
rect 24581 39049 24593 39083
rect 24627 39049 24639 39083
rect 24581 39043 24639 39049
rect 23937 38947 23995 38953
rect 23937 38913 23949 38947
rect 23983 38944 23995 38947
rect 24596 38944 24624 39043
rect 24949 38947 25007 38953
rect 24949 38944 24961 38947
rect 23983 38916 24624 38944
rect 24872 38916 24961 38944
rect 23983 38913 23995 38916
rect 23937 38907 23995 38913
rect 20622 38876 20628 38888
rect 19935 38848 20300 38876
rect 20583 38848 20628 38876
rect 19935 38845 19947 38848
rect 19889 38839 19947 38845
rect 20622 38836 20628 38848
rect 20680 38836 20686 38888
rect 20809 38879 20867 38885
rect 20809 38845 20821 38879
rect 20855 38845 20867 38879
rect 20809 38839 20867 38845
rect 24305 38879 24363 38885
rect 24305 38845 24317 38879
rect 24351 38876 24363 38879
rect 24872 38876 24900 38916
rect 24949 38913 24961 38916
rect 24995 38944 25007 38947
rect 45738 38944 45744 38956
rect 24995 38916 45744 38944
rect 24995 38913 25007 38916
rect 24949 38907 25007 38913
rect 45738 38904 45744 38916
rect 45796 38904 45802 38956
rect 46845 38947 46903 38953
rect 46845 38913 46857 38947
rect 46891 38944 46903 38947
rect 47026 38944 47032 38956
rect 46891 38916 47032 38944
rect 46891 38913 46903 38916
rect 46845 38907 46903 38913
rect 47026 38904 47032 38916
rect 47084 38944 47090 38956
rect 47302 38944 47308 38956
rect 47084 38916 47308 38944
rect 47084 38904 47090 38916
rect 47302 38904 47308 38916
rect 47360 38904 47366 38956
rect 47762 38944 47768 38956
rect 47723 38916 47768 38944
rect 47762 38904 47768 38916
rect 47820 38904 47826 38956
rect 25038 38876 25044 38888
rect 24351 38848 24900 38876
rect 24999 38848 25044 38876
rect 24351 38845 24363 38848
rect 24305 38839 24363 38845
rect 20824 38808 20852 38839
rect 25038 38836 25044 38848
rect 25096 38836 25102 38888
rect 25133 38879 25191 38885
rect 25133 38845 25145 38879
rect 25179 38845 25191 38879
rect 25133 38839 25191 38845
rect 22002 38808 22008 38820
rect 20824 38780 22008 38808
rect 22002 38768 22008 38780
rect 22060 38808 22066 38820
rect 25148 38808 25176 38839
rect 22060 38780 25176 38808
rect 22060 38768 22066 38780
rect 45646 38768 45652 38820
rect 45704 38808 45710 38820
rect 47949 38811 48007 38817
rect 47949 38808 47961 38811
rect 45704 38780 47961 38808
rect 45704 38768 45710 38780
rect 47949 38777 47961 38780
rect 47995 38777 48007 38811
rect 47949 38771 48007 38777
rect 19337 38743 19395 38749
rect 19337 38709 19349 38743
rect 19383 38740 19395 38743
rect 19518 38740 19524 38752
rect 19383 38712 19524 38740
rect 19383 38709 19395 38712
rect 19337 38703 19395 38709
rect 19518 38700 19524 38712
rect 19576 38700 19582 38752
rect 23750 38740 23756 38752
rect 23711 38712 23756 38740
rect 23750 38700 23756 38712
rect 23808 38700 23814 38752
rect 46934 38740 46940 38752
rect 46895 38712 46940 38740
rect 46934 38700 46940 38712
rect 46992 38700 46998 38752
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 24949 38539 25007 38545
rect 24949 38505 24961 38539
rect 24995 38536 25007 38539
rect 25038 38536 25044 38548
rect 24995 38508 25044 38536
rect 24995 38505 25007 38508
rect 24949 38499 25007 38505
rect 25038 38496 25044 38508
rect 25096 38496 25102 38548
rect 17773 38403 17831 38409
rect 17773 38369 17785 38403
rect 17819 38400 17831 38403
rect 18322 38400 18328 38412
rect 17819 38372 18328 38400
rect 17819 38369 17831 38372
rect 17773 38363 17831 38369
rect 18322 38360 18328 38372
rect 18380 38360 18386 38412
rect 19245 38403 19303 38409
rect 19245 38369 19257 38403
rect 19291 38400 19303 38403
rect 21266 38400 21272 38412
rect 19291 38372 21272 38400
rect 19291 38369 19303 38372
rect 19245 38363 19303 38369
rect 21266 38360 21272 38372
rect 21324 38360 21330 38412
rect 23934 38360 23940 38412
rect 23992 38400 23998 38412
rect 24489 38403 24547 38409
rect 24489 38400 24501 38403
rect 23992 38372 24501 38400
rect 23992 38360 23998 38372
rect 24489 38369 24501 38372
rect 24535 38369 24547 38403
rect 24489 38363 24547 38369
rect 46477 38403 46535 38409
rect 46477 38369 46489 38403
rect 46523 38400 46535 38403
rect 46934 38400 46940 38412
rect 46523 38372 46940 38400
rect 46523 38369 46535 38372
rect 46477 38363 46535 38369
rect 46934 38360 46940 38372
rect 46992 38360 46998 38412
rect 48130 38400 48136 38412
rect 48091 38372 48136 38400
rect 48130 38360 48136 38372
rect 48188 38360 48194 38412
rect 23198 38332 23204 38344
rect 23159 38304 23204 38332
rect 23198 38292 23204 38304
rect 23256 38292 23262 38344
rect 24581 38335 24639 38341
rect 24581 38301 24593 38335
rect 24627 38301 24639 38335
rect 24581 38295 24639 38301
rect 19518 38264 19524 38276
rect 19479 38236 19524 38264
rect 19518 38224 19524 38236
rect 19576 38224 19582 38276
rect 20254 38224 20260 38276
rect 20312 38224 20318 38276
rect 24596 38264 24624 38295
rect 45830 38292 45836 38344
rect 45888 38332 45894 38344
rect 46293 38335 46351 38341
rect 46293 38332 46305 38335
rect 45888 38304 46305 38332
rect 45888 38292 45894 38304
rect 46293 38301 46305 38304
rect 46339 38301 46351 38335
rect 46293 38295 46351 38301
rect 24670 38264 24676 38276
rect 24596 38236 24676 38264
rect 24670 38224 24676 38236
rect 24728 38224 24734 38276
rect 16850 38156 16856 38208
rect 16908 38196 16914 38208
rect 17129 38199 17187 38205
rect 17129 38196 17141 38199
rect 16908 38168 17141 38196
rect 16908 38156 16914 38168
rect 17129 38165 17141 38168
rect 17175 38165 17187 38199
rect 17494 38196 17500 38208
rect 17455 38168 17500 38196
rect 17129 38159 17187 38165
rect 17494 38156 17500 38168
rect 17552 38156 17558 38208
rect 17586 38156 17592 38208
rect 17644 38196 17650 38208
rect 17644 38168 17689 38196
rect 17644 38156 17650 38168
rect 19242 38156 19248 38208
rect 19300 38196 19306 38208
rect 20993 38199 21051 38205
rect 20993 38196 21005 38199
rect 19300 38168 21005 38196
rect 19300 38156 19306 38168
rect 20993 38165 21005 38168
rect 21039 38165 21051 38199
rect 23290 38196 23296 38208
rect 23251 38168 23296 38196
rect 20993 38159 21051 38165
rect 23290 38156 23296 38168
rect 23348 38156 23354 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 17586 37992 17592 38004
rect 17547 37964 17592 37992
rect 17586 37952 17592 37964
rect 17644 37952 17650 38004
rect 20254 37992 20260 38004
rect 20215 37964 20260 37992
rect 20254 37952 20260 37964
rect 20312 37952 20318 38004
rect 21177 37995 21235 38001
rect 21177 37961 21189 37995
rect 21223 37992 21235 37995
rect 22370 37992 22376 38004
rect 21223 37964 22376 37992
rect 21223 37961 21235 37964
rect 21177 37955 21235 37961
rect 22370 37952 22376 37964
rect 22428 37992 22434 38004
rect 23198 37992 23204 38004
rect 22428 37964 23204 37992
rect 22428 37952 22434 37964
rect 23198 37952 23204 37964
rect 23256 37952 23262 38004
rect 17218 37884 17224 37936
rect 17276 37924 17282 37936
rect 17957 37927 18015 37933
rect 17957 37924 17969 37927
rect 17276 37896 17969 37924
rect 17276 37884 17282 37896
rect 17957 37893 17969 37896
rect 18003 37893 18015 37927
rect 17957 37887 18015 37893
rect 18248 37896 21864 37924
rect 15286 37816 15292 37868
rect 15344 37856 15350 37868
rect 15933 37859 15991 37865
rect 15933 37856 15945 37859
rect 15344 37828 15945 37856
rect 15344 37816 15350 37828
rect 15933 37825 15945 37828
rect 15979 37825 15991 37859
rect 16850 37856 16856 37868
rect 16811 37828 16856 37856
rect 15933 37819 15991 37825
rect 16850 37816 16856 37828
rect 16908 37816 16914 37868
rect 18046 37788 18052 37800
rect 18007 37760 18052 37788
rect 18046 37748 18052 37760
rect 18104 37748 18110 37800
rect 18248 37797 18276 37896
rect 18690 37816 18696 37868
rect 18748 37856 18754 37868
rect 19242 37856 19248 37868
rect 18748 37828 19248 37856
rect 18748 37816 18754 37828
rect 19242 37816 19248 37828
rect 19300 37856 19306 37868
rect 19337 37859 19395 37865
rect 19337 37856 19349 37859
rect 19300 37828 19349 37856
rect 19300 37816 19306 37828
rect 19337 37825 19349 37828
rect 19383 37825 19395 37859
rect 19337 37819 19395 37825
rect 20165 37859 20223 37865
rect 20165 37825 20177 37859
rect 20211 37856 20223 37859
rect 20530 37856 20536 37868
rect 20211 37828 20536 37856
rect 20211 37825 20223 37828
rect 20165 37819 20223 37825
rect 20530 37816 20536 37828
rect 20588 37816 20594 37868
rect 20990 37856 20996 37868
rect 20903 37828 20996 37856
rect 20990 37816 20996 37828
rect 21048 37856 21054 37868
rect 21542 37856 21548 37868
rect 21048 37828 21548 37856
rect 21048 37816 21054 37828
rect 21542 37816 21548 37828
rect 21600 37816 21606 37868
rect 21836 37865 21864 37896
rect 23290 37884 23296 37936
rect 23348 37924 23354 37936
rect 23348 37896 23690 37924
rect 23348 37884 23354 37896
rect 21821 37859 21879 37865
rect 21821 37825 21833 37859
rect 21867 37856 21879 37859
rect 22278 37856 22284 37868
rect 21867 37828 22284 37856
rect 21867 37825 21879 37828
rect 21821 37819 21879 37825
rect 22278 37816 22284 37828
rect 22336 37816 22342 37868
rect 47578 37856 47584 37868
rect 47539 37828 47584 37856
rect 47578 37816 47584 37828
rect 47636 37816 47642 37868
rect 18233 37791 18291 37797
rect 18233 37757 18245 37791
rect 18279 37757 18291 37791
rect 18233 37751 18291 37757
rect 19429 37791 19487 37797
rect 19429 37757 19441 37791
rect 19475 37757 19487 37791
rect 19429 37751 19487 37757
rect 19705 37791 19763 37797
rect 19705 37757 19717 37791
rect 19751 37788 19763 37791
rect 20622 37788 20628 37800
rect 19751 37760 20628 37788
rect 19751 37757 19763 37760
rect 19705 37751 19763 37757
rect 15838 37680 15844 37732
rect 15896 37720 15902 37732
rect 16669 37723 16727 37729
rect 16669 37720 16681 37723
rect 15896 37692 16681 37720
rect 15896 37680 15902 37692
rect 16669 37689 16681 37692
rect 16715 37689 16727 37723
rect 16669 37683 16727 37689
rect 19334 37680 19340 37732
rect 19392 37720 19398 37732
rect 19444 37720 19472 37751
rect 20622 37748 20628 37760
rect 20680 37748 20686 37800
rect 21266 37748 21272 37800
rect 21324 37788 21330 37800
rect 22925 37791 22983 37797
rect 22925 37788 22937 37791
rect 21324 37760 22937 37788
rect 21324 37748 21330 37760
rect 22925 37757 22937 37760
rect 22971 37757 22983 37791
rect 22925 37751 22983 37757
rect 23201 37791 23259 37797
rect 23201 37757 23213 37791
rect 23247 37788 23259 37791
rect 23750 37788 23756 37800
rect 23247 37760 23756 37788
rect 23247 37757 23259 37760
rect 23201 37751 23259 37757
rect 23750 37748 23756 37760
rect 23808 37748 23814 37800
rect 19392 37692 19472 37720
rect 19392 37680 19398 37692
rect 16025 37655 16083 37661
rect 16025 37621 16037 37655
rect 16071 37652 16083 37655
rect 16574 37652 16580 37664
rect 16071 37624 16580 37652
rect 16071 37621 16083 37624
rect 16025 37615 16083 37621
rect 16574 37612 16580 37624
rect 16632 37612 16638 37664
rect 21358 37612 21364 37664
rect 21416 37652 21422 37664
rect 22002 37652 22008 37664
rect 21416 37624 22008 37652
rect 21416 37612 21422 37624
rect 22002 37612 22008 37624
rect 22060 37612 22066 37664
rect 24670 37652 24676 37664
rect 24631 37624 24676 37652
rect 24670 37612 24676 37624
rect 24728 37612 24734 37664
rect 47026 37652 47032 37664
rect 46987 37624 47032 37652
rect 47026 37612 47032 37624
rect 47084 37612 47090 37664
rect 47670 37652 47676 37664
rect 47631 37624 47676 37652
rect 47670 37612 47676 37624
rect 47728 37612 47734 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 17313 37451 17371 37457
rect 17313 37417 17325 37451
rect 17359 37448 17371 37451
rect 17494 37448 17500 37460
rect 17359 37420 17500 37448
rect 17359 37417 17371 37420
rect 17313 37411 17371 37417
rect 17494 37408 17500 37420
rect 17552 37408 17558 37460
rect 18046 37408 18052 37460
rect 18104 37448 18110 37460
rect 18233 37451 18291 37457
rect 18233 37448 18245 37451
rect 18104 37420 18245 37448
rect 18104 37408 18110 37420
rect 18233 37417 18245 37420
rect 18279 37417 18291 37451
rect 18233 37411 18291 37417
rect 15838 37312 15844 37324
rect 15799 37284 15844 37312
rect 15838 37272 15844 37284
rect 15896 37272 15902 37324
rect 18046 37312 18052 37324
rect 18007 37284 18052 37312
rect 18046 37272 18052 37284
rect 18104 37272 18110 37324
rect 20349 37315 20407 37321
rect 20349 37281 20361 37315
rect 20395 37312 20407 37315
rect 21545 37315 21603 37321
rect 21545 37312 21557 37315
rect 20395 37284 21557 37312
rect 20395 37281 20407 37284
rect 20349 37275 20407 37281
rect 21545 37281 21557 37284
rect 21591 37281 21603 37315
rect 48130 37312 48136 37324
rect 48091 37284 48136 37312
rect 21545 37275 21603 37281
rect 48130 37272 48136 37284
rect 48188 37272 48194 37324
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 2041 37247 2099 37253
rect 2041 37244 2053 37247
rect 1820 37216 2053 37244
rect 1820 37204 1826 37216
rect 2041 37213 2053 37216
rect 2087 37213 2099 37247
rect 2041 37207 2099 37213
rect 14182 37204 14188 37256
rect 14240 37244 14246 37256
rect 15565 37247 15623 37253
rect 15565 37244 15577 37247
rect 14240 37216 15577 37244
rect 14240 37204 14246 37216
rect 15565 37213 15577 37216
rect 15611 37213 15623 37247
rect 15565 37207 15623 37213
rect 17494 37204 17500 37256
rect 17552 37244 17558 37256
rect 17957 37247 18015 37253
rect 17957 37244 17969 37247
rect 17552 37216 17969 37244
rect 17552 37204 17558 37216
rect 17957 37213 17969 37216
rect 18003 37213 18015 37247
rect 20530 37244 20536 37256
rect 20491 37216 20536 37244
rect 17957 37207 18015 37213
rect 20530 37204 20536 37216
rect 20588 37204 20594 37256
rect 20717 37247 20775 37253
rect 20717 37213 20729 37247
rect 20763 37213 20775 37247
rect 20717 37207 20775 37213
rect 20809 37247 20867 37253
rect 20809 37213 20821 37247
rect 20855 37244 20867 37247
rect 20898 37244 20904 37256
rect 20855 37216 20904 37244
rect 20855 37213 20867 37216
rect 20809 37207 20867 37213
rect 16574 37136 16580 37188
rect 16632 37136 16638 37188
rect 20732 37176 20760 37207
rect 20898 37204 20904 37216
rect 20956 37204 20962 37256
rect 21266 37244 21272 37256
rect 21227 37216 21272 37244
rect 21266 37204 21272 37216
rect 21324 37204 21330 37256
rect 22646 37204 22652 37256
rect 22704 37204 22710 37256
rect 25501 37247 25559 37253
rect 25501 37213 25513 37247
rect 25547 37213 25559 37247
rect 25501 37207 25559 37213
rect 20456 37148 20760 37176
rect 12618 37068 12624 37120
rect 12676 37108 12682 37120
rect 20456 37108 20484 37148
rect 12676 37080 20484 37108
rect 12676 37068 12682 37080
rect 20530 37068 20536 37120
rect 20588 37108 20594 37120
rect 22922 37108 22928 37120
rect 20588 37080 22928 37108
rect 20588 37068 20594 37080
rect 22922 37068 22928 37080
rect 22980 37068 22986 37120
rect 23017 37111 23075 37117
rect 23017 37077 23029 37111
rect 23063 37108 23075 37111
rect 23106 37108 23112 37120
rect 23063 37080 23112 37108
rect 23063 37077 23075 37080
rect 23017 37071 23075 37077
rect 23106 37068 23112 37080
rect 23164 37068 23170 37120
rect 25516 37108 25544 37207
rect 28442 37204 28448 37256
rect 28500 37244 28506 37256
rect 28537 37247 28595 37253
rect 28537 37244 28549 37247
rect 28500 37216 28549 37244
rect 28500 37204 28506 37216
rect 28537 37213 28549 37216
rect 28583 37213 28595 37247
rect 28537 37207 28595 37213
rect 46293 37247 46351 37253
rect 46293 37213 46305 37247
rect 46339 37213 46351 37247
rect 46293 37207 46351 37213
rect 25774 37176 25780 37188
rect 25735 37148 25780 37176
rect 25774 37136 25780 37148
rect 25832 37136 25838 37188
rect 27062 37176 27068 37188
rect 27002 37148 27068 37176
rect 27062 37136 27068 37148
rect 27120 37136 27126 37188
rect 27890 37176 27896 37188
rect 27172 37148 27896 37176
rect 27172 37108 27200 37148
rect 27890 37136 27896 37148
rect 27948 37136 27954 37188
rect 25516 37080 27200 37108
rect 27246 37068 27252 37120
rect 27304 37108 27310 37120
rect 28626 37108 28632 37120
rect 27304 37080 27349 37108
rect 28587 37080 28632 37108
rect 27304 37068 27310 37080
rect 28626 37068 28632 37080
rect 28684 37068 28690 37120
rect 46308 37108 46336 37207
rect 46477 37179 46535 37185
rect 46477 37145 46489 37179
rect 46523 37176 46535 37179
rect 47670 37176 47676 37188
rect 46523 37148 47676 37176
rect 46523 37145 46535 37148
rect 46477 37139 46535 37145
rect 47670 37136 47676 37148
rect 47728 37136 47734 37188
rect 47026 37108 47032 37120
rect 46308 37080 47032 37108
rect 47026 37068 47032 37080
rect 47084 37068 47090 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 9490 36864 9496 36916
rect 9548 36904 9554 36916
rect 22005 36907 22063 36913
rect 9548 36876 18736 36904
rect 9548 36864 9554 36876
rect 15194 36796 15200 36848
rect 15252 36796 15258 36848
rect 18325 36839 18383 36845
rect 18325 36836 18337 36839
rect 17420 36808 18337 36836
rect 1762 36768 1768 36780
rect 1723 36740 1768 36768
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 17420 36777 17448 36808
rect 18325 36805 18337 36808
rect 18371 36805 18383 36839
rect 18325 36799 18383 36805
rect 17405 36771 17463 36777
rect 17405 36737 17417 36771
rect 17451 36737 17463 36771
rect 17405 36731 17463 36737
rect 1949 36703 2007 36709
rect 1949 36669 1961 36703
rect 1995 36700 2007 36703
rect 2222 36700 2228 36712
rect 1995 36672 2228 36700
rect 1995 36669 2007 36672
rect 1949 36663 2007 36669
rect 2222 36660 2228 36672
rect 2280 36660 2286 36712
rect 2774 36700 2780 36712
rect 2735 36672 2780 36700
rect 2774 36660 2780 36672
rect 2832 36660 2838 36712
rect 14182 36660 14188 36712
rect 14240 36700 14246 36712
rect 14369 36703 14427 36709
rect 14369 36700 14381 36703
rect 14240 36672 14381 36700
rect 14240 36660 14246 36672
rect 14369 36669 14381 36672
rect 14415 36669 14427 36703
rect 14369 36663 14427 36669
rect 14645 36703 14703 36709
rect 14645 36669 14657 36703
rect 14691 36700 14703 36703
rect 16482 36700 16488 36712
rect 14691 36672 16488 36700
rect 14691 36669 14703 36672
rect 14645 36663 14703 36669
rect 16482 36660 16488 36672
rect 16540 36660 16546 36712
rect 16022 36592 16028 36644
rect 16080 36632 16086 36644
rect 16117 36635 16175 36641
rect 16117 36632 16129 36635
rect 16080 36604 16129 36632
rect 16080 36592 16086 36604
rect 16117 36601 16129 36604
rect 16163 36632 16175 36635
rect 17420 36632 17448 36731
rect 17494 36728 17500 36780
rect 17552 36768 17558 36780
rect 17681 36771 17739 36777
rect 17681 36768 17693 36771
rect 17552 36740 17693 36768
rect 17552 36728 17558 36740
rect 17681 36737 17693 36740
rect 17727 36768 17739 36771
rect 18141 36771 18199 36777
rect 18141 36768 18153 36771
rect 17727 36740 18153 36768
rect 17727 36737 17739 36740
rect 17681 36731 17739 36737
rect 18141 36737 18153 36740
rect 18187 36737 18199 36771
rect 18141 36731 18199 36737
rect 17589 36703 17647 36709
rect 17589 36669 17601 36703
rect 17635 36700 17647 36703
rect 18046 36700 18052 36712
rect 17635 36672 18052 36700
rect 17635 36669 17647 36672
rect 17589 36663 17647 36669
rect 18046 36660 18052 36672
rect 18104 36700 18110 36712
rect 18598 36700 18604 36712
rect 18104 36672 18604 36700
rect 18104 36660 18110 36672
rect 18598 36660 18604 36672
rect 18656 36660 18662 36712
rect 18708 36700 18736 36876
rect 22005 36873 22017 36907
rect 22051 36873 22063 36907
rect 22646 36904 22652 36916
rect 22607 36876 22652 36904
rect 22005 36867 22063 36873
rect 21542 36728 21548 36780
rect 21600 36768 21606 36780
rect 21821 36771 21879 36777
rect 21821 36768 21833 36771
rect 21600 36740 21833 36768
rect 21600 36728 21606 36740
rect 21821 36737 21833 36740
rect 21867 36737 21879 36771
rect 22020 36768 22048 36867
rect 22646 36864 22652 36876
rect 22704 36864 22710 36916
rect 22922 36864 22928 36916
rect 22980 36904 22986 36916
rect 23293 36907 23351 36913
rect 23293 36904 23305 36907
rect 22980 36876 23305 36904
rect 22980 36864 22986 36876
rect 23293 36873 23305 36876
rect 23339 36873 23351 36907
rect 23293 36867 23351 36873
rect 23382 36864 23388 36916
rect 23440 36904 23446 36916
rect 25314 36904 25320 36916
rect 23440 36876 25320 36904
rect 23440 36864 23446 36876
rect 25314 36864 25320 36876
rect 25372 36864 25378 36916
rect 25774 36904 25780 36916
rect 25735 36876 25780 36904
rect 25774 36864 25780 36876
rect 25832 36864 25838 36916
rect 27062 36904 27068 36916
rect 27023 36876 27068 36904
rect 27062 36864 27068 36876
rect 27120 36864 27126 36916
rect 25682 36836 25688 36848
rect 22572 36808 25688 36836
rect 22572 36777 22600 36808
rect 25682 36796 25688 36808
rect 25740 36836 25746 36848
rect 28442 36836 28448 36848
rect 25740 36808 28448 36836
rect 25740 36796 25746 36808
rect 22557 36771 22615 36777
rect 22557 36768 22569 36771
rect 22020 36740 22569 36768
rect 21821 36731 21879 36737
rect 22557 36737 22569 36740
rect 22603 36737 22615 36771
rect 22557 36731 22615 36737
rect 23106 36728 23112 36780
rect 23164 36768 23170 36780
rect 23845 36771 23903 36777
rect 23845 36768 23857 36771
rect 23164 36740 23857 36768
rect 23164 36728 23170 36740
rect 23845 36737 23857 36740
rect 23891 36737 23903 36771
rect 23845 36731 23903 36737
rect 24029 36771 24087 36777
rect 24029 36737 24041 36771
rect 24075 36737 24087 36771
rect 24029 36731 24087 36737
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36768 24823 36771
rect 24854 36768 24860 36780
rect 24811 36740 24860 36768
rect 24811 36737 24823 36740
rect 24765 36731 24823 36737
rect 23569 36703 23627 36709
rect 18708 36672 22094 36700
rect 16163 36604 17448 36632
rect 22066 36632 22094 36672
rect 23569 36669 23581 36703
rect 23615 36700 23627 36703
rect 23658 36700 23664 36712
rect 23615 36672 23664 36700
rect 23615 36669 23627 36672
rect 23569 36663 23627 36669
rect 23658 36660 23664 36672
rect 23716 36660 23722 36712
rect 23753 36703 23811 36709
rect 23753 36669 23765 36703
rect 23799 36700 23811 36703
rect 23934 36700 23940 36712
rect 23799 36672 23940 36700
rect 23799 36669 23811 36672
rect 23753 36663 23811 36669
rect 23934 36660 23940 36672
rect 23992 36660 23998 36712
rect 24044 36700 24072 36731
rect 24854 36728 24860 36740
rect 24912 36728 24918 36780
rect 24946 36728 24952 36780
rect 25004 36768 25010 36780
rect 25961 36771 26019 36777
rect 25004 36740 25049 36768
rect 25004 36728 25010 36740
rect 25961 36737 25973 36771
rect 26007 36768 26019 36771
rect 26142 36768 26148 36780
rect 26007 36740 26148 36768
rect 26007 36737 26019 36740
rect 25961 36731 26019 36737
rect 26142 36728 26148 36740
rect 26200 36728 26206 36780
rect 26988 36777 27016 36808
rect 28442 36796 28448 36808
rect 28500 36796 28506 36848
rect 28626 36796 28632 36848
rect 28684 36796 28690 36848
rect 26973 36771 27031 36777
rect 26973 36737 26985 36771
rect 27019 36737 27031 36771
rect 27890 36768 27896 36780
rect 27851 36740 27896 36768
rect 26973 36731 27031 36737
rect 27890 36728 27896 36740
rect 27948 36728 27954 36780
rect 25133 36703 25191 36709
rect 25133 36700 25145 36703
rect 24044 36672 25145 36700
rect 25133 36669 25145 36672
rect 25179 36700 25191 36703
rect 26050 36700 26056 36712
rect 25179 36672 26056 36700
rect 25179 36669 25191 36672
rect 25133 36663 25191 36669
rect 26050 36660 26056 36672
rect 26108 36660 26114 36712
rect 26237 36703 26295 36709
rect 26237 36669 26249 36703
rect 26283 36669 26295 36703
rect 28166 36700 28172 36712
rect 28127 36672 28172 36700
rect 26237 36663 26295 36669
rect 25038 36632 25044 36644
rect 22066 36604 25044 36632
rect 16163 36601 16175 36604
rect 16117 36595 16175 36601
rect 25038 36592 25044 36604
rect 25096 36592 25102 36644
rect 26252 36632 26280 36663
rect 28166 36660 28172 36672
rect 28224 36660 28230 36712
rect 27706 36632 27712 36644
rect 25884 36604 27712 36632
rect 17221 36567 17279 36573
rect 17221 36533 17233 36567
rect 17267 36564 17279 36567
rect 17402 36564 17408 36576
rect 17267 36536 17408 36564
rect 17267 36533 17279 36536
rect 17221 36527 17279 36533
rect 17402 36524 17408 36536
rect 17460 36524 17466 36576
rect 18414 36524 18420 36576
rect 18472 36564 18478 36576
rect 18509 36567 18567 36573
rect 18509 36564 18521 36567
rect 18472 36536 18521 36564
rect 18472 36524 18478 36536
rect 18509 36533 18521 36536
rect 18555 36533 18567 36567
rect 18509 36527 18567 36533
rect 18598 36524 18604 36576
rect 18656 36564 18662 36576
rect 23382 36564 23388 36576
rect 18656 36536 23388 36564
rect 18656 36524 18662 36536
rect 23382 36524 23388 36536
rect 23440 36524 23446 36576
rect 23566 36524 23572 36576
rect 23624 36564 23630 36576
rect 23661 36567 23719 36573
rect 23661 36564 23673 36567
rect 23624 36536 23673 36564
rect 23624 36524 23630 36536
rect 23661 36533 23673 36536
rect 23707 36533 23719 36567
rect 23661 36527 23719 36533
rect 23934 36524 23940 36576
rect 23992 36564 23998 36576
rect 25884 36564 25912 36604
rect 27706 36592 27712 36604
rect 27764 36592 27770 36644
rect 23992 36536 25912 36564
rect 23992 36524 23998 36536
rect 25958 36524 25964 36576
rect 26016 36564 26022 36576
rect 26145 36567 26203 36573
rect 26145 36564 26157 36567
rect 26016 36536 26157 36564
rect 26016 36524 26022 36536
rect 26145 36533 26157 36536
rect 26191 36533 26203 36567
rect 26145 36527 26203 36533
rect 27982 36524 27988 36576
rect 28040 36564 28046 36576
rect 28810 36564 28816 36576
rect 28040 36536 28816 36564
rect 28040 36524 28046 36536
rect 28810 36524 28816 36536
rect 28868 36564 28874 36576
rect 29641 36567 29699 36573
rect 29641 36564 29653 36567
rect 28868 36536 29653 36564
rect 28868 36524 28874 36536
rect 29641 36533 29653 36536
rect 29687 36533 29699 36567
rect 29641 36527 29699 36533
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 2222 36360 2228 36372
rect 2183 36332 2228 36360
rect 2222 36320 2228 36332
rect 2280 36320 2286 36372
rect 15194 36360 15200 36372
rect 15155 36332 15200 36360
rect 15194 36320 15200 36332
rect 15252 36320 15258 36372
rect 15562 36320 15568 36372
rect 15620 36360 15626 36372
rect 16482 36360 16488 36372
rect 15620 36332 16344 36360
rect 16443 36332 16488 36360
rect 15620 36320 15626 36332
rect 10962 36252 10968 36304
rect 11020 36292 11026 36304
rect 16316 36292 16344 36332
rect 16482 36320 16488 36332
rect 16540 36320 16546 36372
rect 17497 36363 17555 36369
rect 17497 36329 17509 36363
rect 17543 36360 17555 36363
rect 23293 36363 23351 36369
rect 17543 36332 22692 36360
rect 17543 36329 17555 36332
rect 17497 36323 17555 36329
rect 18601 36295 18659 36301
rect 18601 36292 18613 36295
rect 11020 36264 16160 36292
rect 16316 36264 18613 36292
rect 11020 36252 11026 36264
rect 15562 36184 15568 36236
rect 15620 36224 15626 36236
rect 16022 36224 16028 36236
rect 15620 36196 15884 36224
rect 15983 36196 16028 36224
rect 15620 36184 15626 36196
rect 2133 36159 2191 36165
rect 2133 36125 2145 36159
rect 2179 36156 2191 36159
rect 2222 36156 2228 36168
rect 2179 36128 2228 36156
rect 2179 36125 2191 36128
rect 2133 36119 2191 36125
rect 2222 36116 2228 36128
rect 2280 36116 2286 36168
rect 15105 36159 15163 36165
rect 15105 36125 15117 36159
rect 15151 36156 15163 36159
rect 15286 36156 15292 36168
rect 15151 36128 15292 36156
rect 15151 36125 15163 36128
rect 15105 36119 15163 36125
rect 15286 36116 15292 36128
rect 15344 36116 15350 36168
rect 15749 36159 15807 36165
rect 15749 36125 15761 36159
rect 15795 36125 15807 36159
rect 15856 36154 15884 36196
rect 16022 36184 16028 36196
rect 16080 36184 16086 36236
rect 16132 36233 16160 36264
rect 18601 36261 18613 36264
rect 18647 36292 18659 36295
rect 22554 36292 22560 36304
rect 18647 36264 22560 36292
rect 18647 36261 18659 36264
rect 18601 36255 18659 36261
rect 22554 36252 22560 36264
rect 22612 36252 22618 36304
rect 22664 36292 22692 36332
rect 23293 36329 23305 36363
rect 23339 36360 23351 36363
rect 23658 36360 23664 36372
rect 23339 36332 23664 36360
rect 23339 36329 23351 36332
rect 23293 36323 23351 36329
rect 23658 36320 23664 36332
rect 23716 36320 23722 36372
rect 25317 36363 25375 36369
rect 25317 36329 25329 36363
rect 25363 36360 25375 36363
rect 25774 36360 25780 36372
rect 25363 36332 25780 36360
rect 25363 36329 25375 36332
rect 25317 36323 25375 36329
rect 25774 36320 25780 36332
rect 25832 36320 25838 36372
rect 25958 36360 25964 36372
rect 25919 36332 25964 36360
rect 25958 36320 25964 36332
rect 26016 36320 26022 36372
rect 28166 36320 28172 36372
rect 28224 36360 28230 36372
rect 28445 36363 28503 36369
rect 28445 36360 28457 36363
rect 28224 36332 28457 36360
rect 28224 36320 28230 36332
rect 28445 36329 28457 36332
rect 28491 36329 28503 36363
rect 28445 36323 28503 36329
rect 23566 36292 23572 36304
rect 22664 36264 23572 36292
rect 23566 36252 23572 36264
rect 23624 36252 23630 36304
rect 27798 36252 27804 36304
rect 27856 36292 27862 36304
rect 29178 36292 29184 36304
rect 27856 36264 29184 36292
rect 27856 36252 27862 36264
rect 29178 36252 29184 36264
rect 29236 36252 29242 36304
rect 16117 36227 16175 36233
rect 16117 36193 16129 36227
rect 16163 36193 16175 36227
rect 16117 36187 16175 36193
rect 16482 36184 16488 36236
rect 16540 36224 16546 36236
rect 17402 36224 17408 36236
rect 16540 36196 17264 36224
rect 17363 36196 17408 36224
rect 16540 36184 16546 36196
rect 15921 36157 15979 36163
rect 15921 36154 15933 36157
rect 15856 36126 15933 36154
rect 15749 36119 15807 36125
rect 15921 36123 15933 36126
rect 15967 36123 15979 36157
rect 15764 36088 15792 36119
rect 15921 36117 15979 36123
rect 16206 36116 16212 36168
rect 16264 36156 16270 36168
rect 16301 36159 16359 36165
rect 16301 36156 16313 36159
rect 16264 36128 16313 36156
rect 16264 36116 16270 36128
rect 16301 36125 16313 36128
rect 16347 36125 16359 36159
rect 16301 36119 16359 36125
rect 17034 36116 17040 36168
rect 17092 36156 17098 36168
rect 17129 36159 17187 36165
rect 17129 36156 17141 36159
rect 17092 36128 17141 36156
rect 17092 36116 17098 36128
rect 17129 36125 17141 36128
rect 17175 36125 17187 36159
rect 17236 36156 17264 36196
rect 17402 36184 17408 36196
rect 17460 36184 17466 36236
rect 23106 36224 23112 36236
rect 18248 36196 19288 36224
rect 23067 36196 23112 36224
rect 18248 36156 18276 36196
rect 17236 36128 18276 36156
rect 17129 36119 17187 36125
rect 18322 36116 18328 36168
rect 18380 36156 18386 36168
rect 18417 36159 18475 36165
rect 18417 36156 18429 36159
rect 18380 36128 18429 36156
rect 18380 36116 18386 36128
rect 18417 36125 18429 36128
rect 18463 36156 18475 36159
rect 19058 36156 19064 36168
rect 18463 36128 19064 36156
rect 18463 36125 18475 36128
rect 18417 36119 18475 36125
rect 19058 36116 19064 36128
rect 19116 36116 19122 36168
rect 19260 36165 19288 36196
rect 23106 36184 23112 36196
rect 23164 36224 23170 36236
rect 23164 36196 24624 36224
rect 23164 36184 23170 36196
rect 19245 36159 19303 36165
rect 19245 36125 19257 36159
rect 19291 36125 19303 36159
rect 19245 36119 19303 36125
rect 20073 36159 20131 36165
rect 20073 36125 20085 36159
rect 20119 36125 20131 36159
rect 20254 36156 20260 36168
rect 20215 36128 20260 36156
rect 20073 36119 20131 36125
rect 19337 36091 19395 36097
rect 15764 36060 16620 36088
rect 15286 35980 15292 36032
rect 15344 36020 15350 36032
rect 16482 36020 16488 36032
rect 15344 35992 16488 36020
rect 15344 35980 15350 35992
rect 16482 35980 16488 35992
rect 16540 35980 16546 36032
rect 16592 36020 16620 36060
rect 19337 36057 19349 36091
rect 19383 36088 19395 36091
rect 19978 36088 19984 36100
rect 19383 36060 19984 36088
rect 19383 36057 19395 36060
rect 19337 36051 19395 36057
rect 19978 36048 19984 36060
rect 20036 36048 20042 36100
rect 20088 36088 20116 36119
rect 20254 36116 20260 36128
rect 20312 36116 20318 36168
rect 20349 36159 20407 36165
rect 20349 36125 20361 36159
rect 20395 36156 20407 36159
rect 23566 36156 23572 36168
rect 20395 36128 21956 36156
rect 23527 36128 23572 36156
rect 20395 36125 20407 36128
rect 20349 36119 20407 36125
rect 21928 36100 21956 36128
rect 23566 36116 23572 36128
rect 23624 36116 23630 36168
rect 24596 36165 24624 36196
rect 25038 36184 25044 36236
rect 25096 36224 25102 36236
rect 28077 36227 28135 36233
rect 28077 36224 28089 36227
rect 25096 36196 28089 36224
rect 25096 36184 25102 36196
rect 28077 36193 28089 36196
rect 28123 36193 28135 36227
rect 28077 36187 28135 36193
rect 24581 36159 24639 36165
rect 24581 36125 24593 36159
rect 24627 36125 24639 36159
rect 24581 36119 24639 36125
rect 24854 36116 24860 36168
rect 24912 36156 24918 36168
rect 25225 36159 25283 36165
rect 25225 36156 25237 36159
rect 24912 36128 25237 36156
rect 24912 36116 24918 36128
rect 25225 36125 25237 36128
rect 25271 36125 25283 36159
rect 25409 36159 25467 36165
rect 25409 36156 25421 36159
rect 25225 36119 25283 36125
rect 25332 36128 25421 36156
rect 20530 36088 20536 36100
rect 20088 36060 20536 36088
rect 20530 36048 20536 36060
rect 20588 36048 20594 36100
rect 21910 36048 21916 36100
rect 21968 36088 21974 36100
rect 24397 36091 24455 36097
rect 21968 36060 22094 36088
rect 21968 36048 21974 36060
rect 17681 36023 17739 36029
rect 17681 36020 17693 36023
rect 16592 35992 17693 36020
rect 17681 35989 17693 35992
rect 17727 35989 17739 36023
rect 17681 35983 17739 35989
rect 19426 35980 19432 36032
rect 19484 36020 19490 36032
rect 19889 36023 19947 36029
rect 19889 36020 19901 36023
rect 19484 35992 19901 36020
rect 19484 35980 19490 35992
rect 19889 35989 19901 35992
rect 19935 35989 19947 36023
rect 22066 36020 22094 36060
rect 24397 36057 24409 36091
rect 24443 36088 24455 36091
rect 24946 36088 24952 36100
rect 24443 36060 24952 36088
rect 24443 36057 24455 36060
rect 24397 36051 24455 36057
rect 24946 36048 24952 36060
rect 25004 36088 25010 36100
rect 25332 36088 25360 36128
rect 25409 36125 25421 36128
rect 25455 36156 25467 36159
rect 25455 36128 25728 36156
rect 25455 36125 25467 36128
rect 25409 36119 25467 36125
rect 25004 36060 25360 36088
rect 25004 36048 25010 36060
rect 23382 36020 23388 36032
rect 22066 35992 23388 36020
rect 19889 35983 19947 35989
rect 23382 35980 23388 35992
rect 23440 35980 23446 36032
rect 23477 36023 23535 36029
rect 23477 35989 23489 36023
rect 23523 36020 23535 36023
rect 23750 36020 23756 36032
rect 23523 35992 23756 36020
rect 23523 35989 23535 35992
rect 23477 35983 23535 35989
rect 23750 35980 23756 35992
rect 23808 35980 23814 36032
rect 24762 36020 24768 36032
rect 24723 35992 24768 36020
rect 24762 35980 24768 35992
rect 24820 35980 24826 36032
rect 25700 36020 25728 36128
rect 25866 36116 25872 36168
rect 25924 36156 25930 36168
rect 26050 36156 26056 36168
rect 25924 36128 25969 36156
rect 26011 36128 26056 36156
rect 25924 36116 25930 36128
rect 26050 36116 26056 36128
rect 26108 36116 26114 36168
rect 27709 36159 27767 36165
rect 27709 36125 27721 36159
rect 27755 36125 27767 36159
rect 27709 36119 27767 36125
rect 27724 36088 27752 36119
rect 27798 36116 27804 36168
rect 27856 36156 27862 36168
rect 27893 36159 27951 36165
rect 27893 36156 27905 36159
rect 27856 36128 27905 36156
rect 27856 36116 27862 36128
rect 27893 36125 27905 36128
rect 27939 36125 27951 36159
rect 27893 36119 27951 36125
rect 27982 36116 27988 36168
rect 28040 36156 28046 36168
rect 28261 36159 28319 36165
rect 28040 36128 28085 36156
rect 28040 36116 28046 36128
rect 28261 36125 28273 36159
rect 28307 36125 28319 36159
rect 28261 36119 28319 36125
rect 28166 36088 28172 36100
rect 27724 36060 28172 36088
rect 28166 36048 28172 36060
rect 28224 36048 28230 36100
rect 27246 36020 27252 36032
rect 25700 35992 27252 36020
rect 27246 35980 27252 35992
rect 27304 35980 27310 36032
rect 28074 35980 28080 36032
rect 28132 36020 28138 36032
rect 28276 36020 28304 36119
rect 28442 36116 28448 36168
rect 28500 36156 28506 36168
rect 29549 36159 29607 36165
rect 29549 36156 29561 36159
rect 28500 36128 29561 36156
rect 28500 36116 28506 36128
rect 29549 36125 29561 36128
rect 29595 36125 29607 36159
rect 29549 36119 29607 36125
rect 29638 36020 29644 36032
rect 28132 35992 28304 36020
rect 29599 35992 29644 36020
rect 28132 35980 28138 35992
rect 29638 35980 29644 35992
rect 29696 35980 29702 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 20622 35816 20628 35828
rect 16408 35788 20628 35816
rect 16408 35692 16436 35788
rect 20622 35776 20628 35788
rect 20680 35816 20686 35828
rect 24118 35816 24124 35828
rect 20680 35788 22094 35816
rect 24079 35788 24124 35816
rect 20680 35776 20686 35788
rect 19337 35751 19395 35757
rect 19337 35717 19349 35751
rect 19383 35748 19395 35751
rect 19426 35748 19432 35760
rect 19383 35720 19432 35748
rect 19383 35717 19395 35720
rect 19337 35711 19395 35717
rect 19426 35708 19432 35720
rect 19484 35708 19490 35760
rect 19978 35708 19984 35760
rect 20036 35708 20042 35760
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 15289 35683 15347 35689
rect 15289 35649 15301 35683
rect 15335 35680 15347 35683
rect 16390 35680 16396 35692
rect 15335 35652 16396 35680
rect 15335 35649 15347 35652
rect 15289 35643 15347 35649
rect 16390 35640 16396 35652
rect 16448 35640 16454 35692
rect 22066 35680 22094 35788
rect 24118 35776 24124 35788
rect 24176 35776 24182 35828
rect 24673 35819 24731 35825
rect 24673 35816 24685 35819
rect 24320 35788 24685 35816
rect 23750 35748 23756 35760
rect 23711 35720 23756 35748
rect 23750 35708 23756 35720
rect 23808 35708 23814 35760
rect 23969 35751 24027 35757
rect 23969 35717 23981 35751
rect 24015 35748 24027 35751
rect 24320 35748 24348 35788
rect 24673 35785 24685 35788
rect 24719 35785 24731 35819
rect 24673 35779 24731 35785
rect 26436 35788 31248 35816
rect 26436 35760 26464 35788
rect 26418 35748 26424 35760
rect 24015 35720 24348 35748
rect 24504 35720 26424 35748
rect 24015 35717 24027 35720
rect 23969 35711 24027 35717
rect 24504 35680 24532 35720
rect 26418 35708 26424 35720
rect 26476 35708 26482 35760
rect 27890 35748 27896 35760
rect 27632 35720 27896 35748
rect 22066 35652 24532 35680
rect 24581 35683 24639 35689
rect 24581 35649 24593 35683
rect 24627 35649 24639 35683
rect 24762 35680 24768 35692
rect 24723 35652 24768 35680
rect 24581 35643 24639 35649
rect 14182 35572 14188 35624
rect 14240 35612 14246 35624
rect 19061 35615 19119 35621
rect 19061 35612 19073 35615
rect 14240 35584 19073 35612
rect 14240 35572 14246 35584
rect 19061 35581 19073 35584
rect 19107 35612 19119 35615
rect 20714 35612 20720 35624
rect 19107 35584 20720 35612
rect 19107 35581 19119 35584
rect 19061 35575 19119 35581
rect 20714 35572 20720 35584
rect 20772 35612 20778 35624
rect 21266 35612 21272 35624
rect 20772 35584 21272 35612
rect 20772 35572 20778 35584
rect 21266 35572 21272 35584
rect 21324 35572 21330 35624
rect 24596 35612 24624 35643
rect 24762 35640 24768 35652
rect 24820 35640 24826 35692
rect 25682 35640 25688 35692
rect 25740 35680 25746 35692
rect 27632 35689 27660 35720
rect 27890 35708 27896 35720
rect 27948 35708 27954 35760
rect 29638 35748 29644 35760
rect 29118 35720 29644 35748
rect 29638 35708 29644 35720
rect 29696 35708 29702 35760
rect 31220 35689 31248 35788
rect 25777 35683 25835 35689
rect 25777 35680 25789 35683
rect 25740 35652 25789 35680
rect 25740 35640 25746 35652
rect 25777 35649 25789 35652
rect 25823 35649 25835 35683
rect 25777 35643 25835 35649
rect 27617 35683 27675 35689
rect 27617 35649 27629 35683
rect 27663 35649 27675 35683
rect 27617 35643 27675 35649
rect 31205 35683 31263 35689
rect 31205 35649 31217 35683
rect 31251 35680 31263 35683
rect 31294 35680 31300 35692
rect 31251 35652 31300 35680
rect 31251 35649 31263 35652
rect 31205 35643 31263 35649
rect 31294 35640 31300 35652
rect 31352 35640 31358 35692
rect 24854 35612 24860 35624
rect 24596 35584 24860 35612
rect 24854 35572 24860 35584
rect 24912 35572 24918 35624
rect 27893 35615 27951 35621
rect 27893 35581 27905 35615
rect 27939 35612 27951 35615
rect 28350 35612 28356 35624
rect 27939 35584 28356 35612
rect 27939 35581 27951 35584
rect 27893 35575 27951 35581
rect 28350 35572 28356 35584
rect 28408 35572 28414 35624
rect 1397 35479 1455 35485
rect 1397 35445 1409 35479
rect 1443 35476 1455 35479
rect 1486 35476 1492 35488
rect 1443 35448 1492 35476
rect 1443 35445 1455 35448
rect 1397 35439 1455 35445
rect 1486 35436 1492 35448
rect 1544 35436 1550 35488
rect 15381 35479 15439 35485
rect 15381 35445 15393 35479
rect 15427 35476 15439 35479
rect 15470 35476 15476 35488
rect 15427 35448 15476 35476
rect 15427 35445 15439 35448
rect 15381 35439 15439 35445
rect 15470 35436 15476 35448
rect 15528 35436 15534 35488
rect 20806 35436 20812 35488
rect 20864 35476 20870 35488
rect 23934 35476 23940 35488
rect 20864 35448 20909 35476
rect 23895 35448 23940 35476
rect 20864 35436 20870 35448
rect 23934 35436 23940 35448
rect 23992 35436 23998 35488
rect 25869 35479 25927 35485
rect 25869 35445 25881 35479
rect 25915 35476 25927 35479
rect 25958 35476 25964 35488
rect 25915 35448 25964 35476
rect 25915 35445 25927 35448
rect 25869 35439 25927 35445
rect 25958 35436 25964 35448
rect 26016 35436 26022 35488
rect 27706 35436 27712 35488
rect 27764 35476 27770 35488
rect 28258 35476 28264 35488
rect 27764 35448 28264 35476
rect 27764 35436 27770 35448
rect 28258 35436 28264 35448
rect 28316 35436 28322 35488
rect 28902 35436 28908 35488
rect 28960 35476 28966 35488
rect 29365 35479 29423 35485
rect 29365 35476 29377 35479
rect 28960 35448 29377 35476
rect 28960 35436 28966 35448
rect 29365 35445 29377 35448
rect 29411 35445 29423 35479
rect 29365 35439 29423 35445
rect 31202 35436 31208 35488
rect 31260 35476 31266 35488
rect 31297 35479 31355 35485
rect 31297 35476 31309 35479
rect 31260 35448 31309 35476
rect 31260 35436 31266 35448
rect 31297 35445 31309 35448
rect 31343 35445 31355 35479
rect 31297 35439 31355 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 18874 35232 18880 35284
rect 18932 35272 18938 35284
rect 20530 35272 20536 35284
rect 18932 35244 20392 35272
rect 20491 35244 20536 35272
rect 18932 35232 18938 35244
rect 19797 35207 19855 35213
rect 19797 35173 19809 35207
rect 19843 35204 19855 35207
rect 20254 35204 20260 35216
rect 19843 35176 20260 35204
rect 19843 35173 19855 35176
rect 19797 35167 19855 35173
rect 20254 35164 20260 35176
rect 20312 35164 20318 35216
rect 20364 35204 20392 35244
rect 20530 35232 20536 35244
rect 20588 35232 20594 35284
rect 20993 35275 21051 35281
rect 20993 35241 21005 35275
rect 21039 35272 21051 35275
rect 21039 35244 26924 35272
rect 21039 35241 21051 35244
rect 20993 35235 21051 35241
rect 20898 35204 20904 35216
rect 20364 35176 20904 35204
rect 20898 35164 20904 35176
rect 20956 35204 20962 35216
rect 21729 35207 21787 35213
rect 21729 35204 21741 35207
rect 20956 35176 21741 35204
rect 20956 35164 20962 35176
rect 21729 35173 21741 35176
rect 21775 35173 21787 35207
rect 26896 35204 26924 35244
rect 27522 35232 27528 35284
rect 27580 35272 27586 35284
rect 27893 35275 27951 35281
rect 27893 35272 27905 35275
rect 27580 35244 27905 35272
rect 27580 35232 27586 35244
rect 27893 35241 27905 35244
rect 27939 35241 27951 35275
rect 27893 35235 27951 35241
rect 28166 35232 28172 35284
rect 28224 35272 28230 35284
rect 28353 35275 28411 35281
rect 28353 35272 28365 35275
rect 28224 35244 28365 35272
rect 28224 35232 28230 35244
rect 28353 35241 28365 35244
rect 28399 35241 28411 35275
rect 28353 35235 28411 35241
rect 26896 35176 30328 35204
rect 21729 35167 21787 35173
rect 17957 35139 18015 35145
rect 17957 35105 17969 35139
rect 18003 35136 18015 35139
rect 18322 35136 18328 35148
rect 18003 35108 18328 35136
rect 18003 35105 18015 35108
rect 17957 35099 18015 35105
rect 18322 35096 18328 35108
rect 18380 35136 18386 35148
rect 19337 35139 19395 35145
rect 19337 35136 19349 35139
rect 18380 35108 19349 35136
rect 18380 35096 18386 35108
rect 19337 35105 19349 35108
rect 19383 35105 19395 35139
rect 20990 35136 20996 35148
rect 19337 35099 19395 35105
rect 20732 35108 20996 35136
rect 14182 35068 14188 35080
rect 14143 35040 14188 35068
rect 14182 35028 14188 35040
rect 14240 35028 14246 35080
rect 20732 35077 20760 35108
rect 20990 35096 20996 35108
rect 21048 35096 21054 35148
rect 24673 35139 24731 35145
rect 24673 35105 24685 35139
rect 24719 35136 24731 35139
rect 27890 35136 27896 35148
rect 24719 35108 27896 35136
rect 24719 35105 24731 35108
rect 24673 35099 24731 35105
rect 27890 35096 27896 35108
rect 27948 35136 27954 35148
rect 30193 35139 30251 35145
rect 30193 35136 30205 35139
rect 27948 35108 30205 35136
rect 27948 35096 27954 35108
rect 30193 35105 30205 35108
rect 30239 35105 30251 35139
rect 30300 35136 30328 35176
rect 43990 35136 43996 35148
rect 30300 35108 43996 35136
rect 30193 35099 30251 35105
rect 43990 35096 43996 35108
rect 44048 35096 44054 35148
rect 17773 35071 17831 35077
rect 17773 35037 17785 35071
rect 17819 35037 17831 35071
rect 17773 35031 17831 35037
rect 18049 35071 18107 35077
rect 18049 35037 18061 35071
rect 18095 35068 18107 35071
rect 19429 35071 19487 35077
rect 19429 35068 19441 35071
rect 18095 35040 19441 35068
rect 18095 35037 18107 35040
rect 18049 35031 18107 35037
rect 19429 35037 19441 35040
rect 19475 35037 19487 35071
rect 19429 35031 19487 35037
rect 20717 35071 20775 35077
rect 20717 35037 20729 35071
rect 20763 35037 20775 35071
rect 20717 35031 20775 35037
rect 14458 35000 14464 35012
rect 14419 34972 14464 35000
rect 14458 34960 14464 34972
rect 14516 34960 14522 35012
rect 15470 34960 15476 35012
rect 15528 34960 15534 35012
rect 17788 35000 17816 35031
rect 18506 35000 18512 35012
rect 15948 34972 18512 35000
rect 15838 34892 15844 34944
rect 15896 34932 15902 34944
rect 15948 34941 15976 34972
rect 18506 34960 18512 34972
rect 18564 34960 18570 35012
rect 19334 34960 19340 35012
rect 19392 35000 19398 35012
rect 19444 35000 19472 35031
rect 20806 35028 20812 35080
rect 20864 35068 20870 35080
rect 21085 35071 21143 35077
rect 20864 35040 20909 35068
rect 20864 35028 20870 35040
rect 21085 35037 21097 35071
rect 21131 35068 21143 35071
rect 21174 35068 21180 35080
rect 21131 35040 21180 35068
rect 21131 35037 21143 35040
rect 21085 35031 21143 35037
rect 21174 35028 21180 35040
rect 21232 35068 21238 35080
rect 21545 35071 21603 35077
rect 21545 35068 21557 35071
rect 21232 35040 21557 35068
rect 21232 35028 21238 35040
rect 21545 35037 21557 35040
rect 21591 35037 21603 35071
rect 22370 35068 22376 35080
rect 22331 35040 22376 35068
rect 21545 35031 21603 35037
rect 20824 35000 20852 35028
rect 19392 34972 20852 35000
rect 21560 35000 21588 35031
rect 22370 35028 22376 35040
rect 22428 35028 22434 35080
rect 27798 35068 27804 35080
rect 27759 35040 27804 35068
rect 27798 35028 27804 35040
rect 27856 35028 27862 35080
rect 28166 35068 28172 35080
rect 28127 35040 28172 35068
rect 28166 35028 28172 35040
rect 28224 35028 28230 35080
rect 48130 35068 48136 35080
rect 48091 35040 48136 35068
rect 48130 35028 48136 35040
rect 48188 35028 48194 35080
rect 22646 35000 22652 35012
rect 21560 34972 22652 35000
rect 19392 34960 19398 34972
rect 22646 34960 22652 34972
rect 22704 34960 22710 35012
rect 24949 35003 25007 35009
rect 24949 34969 24961 35003
rect 24995 35000 25007 35003
rect 25222 35000 25228 35012
rect 24995 34972 25228 35000
rect 24995 34969 25007 34972
rect 24949 34963 25007 34969
rect 25222 34960 25228 34972
rect 25280 34960 25286 35012
rect 25958 34960 25964 35012
rect 26016 34960 26022 35012
rect 26234 34960 26240 35012
rect 26292 35000 26298 35012
rect 27157 35003 27215 35009
rect 27157 35000 27169 35003
rect 26292 34972 27169 35000
rect 26292 34960 26298 34972
rect 27157 34969 27169 34972
rect 27203 35000 27215 35003
rect 29086 35000 29092 35012
rect 27203 34972 29092 35000
rect 27203 34969 27215 34972
rect 27157 34963 27215 34969
rect 29086 34960 29092 34972
rect 29144 34960 29150 35012
rect 30466 35000 30472 35012
rect 30427 34972 30472 35000
rect 30466 34960 30472 34972
rect 30524 34960 30530 35012
rect 31202 34960 31208 35012
rect 31260 34960 31266 35012
rect 15933 34935 15991 34941
rect 15933 34932 15945 34935
rect 15896 34904 15945 34932
rect 15896 34892 15902 34904
rect 15933 34901 15945 34904
rect 15979 34901 15991 34935
rect 15933 34895 15991 34901
rect 17589 34935 17647 34941
rect 17589 34901 17601 34935
rect 17635 34932 17647 34935
rect 17678 34932 17684 34944
rect 17635 34904 17684 34932
rect 17635 34901 17647 34904
rect 17589 34895 17647 34901
rect 17678 34892 17684 34904
rect 17736 34892 17742 34944
rect 22465 34935 22523 34941
rect 22465 34901 22477 34935
rect 22511 34932 22523 34935
rect 22554 34932 22560 34944
rect 22511 34904 22560 34932
rect 22511 34901 22523 34904
rect 22465 34895 22523 34901
rect 22554 34892 22560 34904
rect 22612 34892 22618 34944
rect 25590 34892 25596 34944
rect 25648 34932 25654 34944
rect 26421 34935 26479 34941
rect 26421 34932 26433 34935
rect 25648 34904 26433 34932
rect 25648 34892 25654 34904
rect 26421 34901 26433 34904
rect 26467 34901 26479 34935
rect 27246 34932 27252 34944
rect 27207 34904 27252 34932
rect 26421 34895 26479 34901
rect 27246 34892 27252 34904
rect 27304 34932 27310 34944
rect 28074 34932 28080 34944
rect 27304 34904 28080 34932
rect 27304 34892 27310 34904
rect 28074 34892 28080 34904
rect 28132 34892 28138 34944
rect 28258 34892 28264 34944
rect 28316 34932 28322 34944
rect 30006 34932 30012 34944
rect 28316 34904 30012 34932
rect 28316 34892 28322 34904
rect 30006 34892 30012 34904
rect 30064 34892 30070 34944
rect 30190 34892 30196 34944
rect 30248 34932 30254 34944
rect 31941 34935 31999 34941
rect 31941 34932 31953 34935
rect 30248 34904 31953 34932
rect 30248 34892 30254 34904
rect 31941 34901 31953 34904
rect 31987 34901 31999 34935
rect 31941 34895 31999 34901
rect 47118 34892 47124 34944
rect 47176 34932 47182 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47176 34904 47961 34932
rect 47176 34892 47182 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 14458 34688 14464 34740
rect 14516 34728 14522 34740
rect 16117 34731 16175 34737
rect 16117 34728 16129 34731
rect 14516 34700 16129 34728
rect 14516 34688 14522 34700
rect 16117 34697 16129 34700
rect 16163 34697 16175 34731
rect 16117 34691 16175 34697
rect 18506 34688 18512 34740
rect 18564 34728 18570 34740
rect 18564 34700 19564 34728
rect 18564 34688 18570 34700
rect 15396 34632 16252 34660
rect 15396 34601 15424 34632
rect 15381 34595 15439 34601
rect 15381 34561 15393 34595
rect 15427 34561 15439 34595
rect 15381 34555 15439 34561
rect 15470 34552 15476 34604
rect 15528 34592 15534 34604
rect 15565 34595 15623 34601
rect 15565 34592 15577 34595
rect 15528 34564 15577 34592
rect 15528 34552 15534 34564
rect 15565 34561 15577 34564
rect 15611 34561 15623 34595
rect 15565 34555 15623 34561
rect 15657 34595 15715 34601
rect 15657 34561 15669 34595
rect 15703 34592 15715 34595
rect 15838 34592 15844 34604
rect 15703 34564 15844 34592
rect 15703 34561 15715 34564
rect 15657 34555 15715 34561
rect 15838 34552 15844 34564
rect 15896 34552 15902 34604
rect 15933 34595 15991 34601
rect 15933 34561 15945 34595
rect 15979 34592 15991 34595
rect 16114 34592 16120 34604
rect 15979 34564 16120 34592
rect 15979 34561 15991 34564
rect 15933 34555 15991 34561
rect 16114 34552 16120 34564
rect 16172 34552 16178 34604
rect 15746 34484 15752 34536
rect 15804 34524 15810 34536
rect 16224 34524 16252 34632
rect 17954 34620 17960 34672
rect 18012 34660 18018 34672
rect 18012 34632 19472 34660
rect 18012 34620 18018 34632
rect 17402 34592 17408 34604
rect 17363 34564 17408 34592
rect 17402 34552 17408 34564
rect 17460 34552 17466 34604
rect 17678 34592 17684 34604
rect 17639 34564 17684 34592
rect 17678 34552 17684 34564
rect 17736 34552 17742 34604
rect 18417 34595 18475 34601
rect 18417 34561 18429 34595
rect 18463 34592 18475 34595
rect 18463 34564 18644 34592
rect 18463 34561 18475 34564
rect 18417 34555 18475 34561
rect 18506 34524 18512 34536
rect 15804 34496 15849 34524
rect 16224 34496 18000 34524
rect 18467 34496 18512 34524
rect 15804 34484 15810 34496
rect 17972 34465 18000 34496
rect 18506 34484 18512 34496
rect 18564 34484 18570 34536
rect 18616 34524 18644 34564
rect 18690 34552 18696 34604
rect 18748 34592 18754 34604
rect 19334 34592 19340 34604
rect 18748 34564 18793 34592
rect 19295 34564 19340 34592
rect 18748 34552 18754 34564
rect 19334 34552 19340 34564
rect 19392 34552 19398 34604
rect 19352 34524 19380 34552
rect 18616 34496 19380 34524
rect 19444 34524 19472 34632
rect 19536 34601 19564 34700
rect 20898 34688 20904 34740
rect 20956 34728 20962 34740
rect 23566 34728 23572 34740
rect 20956 34700 23572 34728
rect 20956 34688 20962 34700
rect 23566 34688 23572 34700
rect 23624 34688 23630 34740
rect 24854 34688 24860 34740
rect 24912 34728 24918 34740
rect 25038 34728 25044 34740
rect 24912 34700 25044 34728
rect 24912 34688 24918 34700
rect 25038 34688 25044 34700
rect 25096 34728 25102 34740
rect 25777 34731 25835 34737
rect 25777 34728 25789 34731
rect 25096 34700 25789 34728
rect 25096 34688 25102 34700
rect 25777 34697 25789 34700
rect 25823 34697 25835 34731
rect 25777 34691 25835 34697
rect 26878 34688 26884 34740
rect 26936 34728 26942 34740
rect 29273 34731 29331 34737
rect 29273 34728 29285 34731
rect 26936 34700 29285 34728
rect 26936 34688 26942 34700
rect 29273 34697 29285 34700
rect 29319 34697 29331 34731
rect 29273 34691 29331 34697
rect 30466 34688 30472 34740
rect 30524 34728 30530 34740
rect 30929 34731 30987 34737
rect 30929 34728 30941 34731
rect 30524 34700 30941 34728
rect 30524 34688 30530 34700
rect 30929 34697 30941 34700
rect 30975 34697 30987 34731
rect 30929 34691 30987 34697
rect 22554 34620 22560 34672
rect 22612 34620 22618 34672
rect 24397 34663 24455 34669
rect 24397 34629 24409 34663
rect 24443 34660 24455 34663
rect 24762 34660 24768 34672
rect 24443 34632 24768 34660
rect 24443 34629 24455 34632
rect 24397 34623 24455 34629
rect 24762 34620 24768 34632
rect 24820 34620 24826 34672
rect 25317 34663 25375 34669
rect 25317 34629 25329 34663
rect 25363 34660 25375 34663
rect 26896 34660 26924 34688
rect 27982 34660 27988 34672
rect 25363 34632 26924 34660
rect 27895 34632 27988 34660
rect 25363 34629 25375 34632
rect 25317 34623 25375 34629
rect 19521 34595 19579 34601
rect 19521 34561 19533 34595
rect 19567 34561 19579 34595
rect 19521 34555 19579 34561
rect 20714 34552 20720 34604
rect 20772 34592 20778 34604
rect 21821 34595 21879 34601
rect 21821 34592 21833 34595
rect 20772 34564 21833 34592
rect 20772 34552 20778 34564
rect 21821 34561 21833 34564
rect 21867 34561 21879 34595
rect 24670 34592 24676 34604
rect 24631 34564 24676 34592
rect 21821 34555 21879 34561
rect 24670 34552 24676 34564
rect 24728 34552 24734 34604
rect 25332 34592 25360 34623
rect 25590 34592 25596 34604
rect 25240 34564 25360 34592
rect 25551 34564 25596 34592
rect 19705 34527 19763 34533
rect 19705 34524 19717 34527
rect 19444 34496 19717 34524
rect 19705 34493 19717 34496
rect 19751 34493 19763 34527
rect 19705 34487 19763 34493
rect 22094 34484 22100 34536
rect 22152 34524 22158 34536
rect 24581 34527 24639 34533
rect 22152 34496 22197 34524
rect 22152 34484 22158 34496
rect 24581 34493 24593 34527
rect 24627 34524 24639 34527
rect 25240 34524 25268 34564
rect 25590 34552 25596 34564
rect 25648 34552 25654 34604
rect 27614 34592 27620 34604
rect 27575 34564 27620 34592
rect 27614 34552 27620 34564
rect 27672 34552 27678 34604
rect 27706 34552 27712 34604
rect 27764 34592 27770 34604
rect 27908 34601 27936 34632
rect 27982 34620 27988 34632
rect 28040 34660 28046 34672
rect 28902 34660 28908 34672
rect 28040 34632 28908 34660
rect 28040 34620 28046 34632
rect 28902 34620 28908 34632
rect 28960 34660 28966 34672
rect 28960 34632 29132 34660
rect 28960 34620 28966 34632
rect 27801 34595 27859 34601
rect 27801 34592 27813 34595
rect 27764 34564 27813 34592
rect 27764 34552 27770 34564
rect 27801 34561 27813 34564
rect 27847 34561 27859 34595
rect 27801 34555 27859 34561
rect 27893 34595 27951 34601
rect 27893 34561 27905 34595
rect 27939 34561 27951 34595
rect 27893 34555 27951 34561
rect 28074 34552 28080 34604
rect 28132 34592 28138 34604
rect 28169 34595 28227 34601
rect 28169 34592 28181 34595
rect 28132 34564 28181 34592
rect 28132 34552 28138 34564
rect 28169 34561 28181 34564
rect 28215 34561 28227 34595
rect 28350 34592 28356 34604
rect 28311 34564 28356 34592
rect 28169 34555 28227 34561
rect 28350 34552 28356 34564
rect 28408 34552 28414 34604
rect 29104 34601 29132 34632
rect 30006 34620 30012 34672
rect 30064 34660 30070 34672
rect 30064 34632 31432 34660
rect 30064 34620 30070 34632
rect 28813 34595 28871 34601
rect 28813 34561 28825 34595
rect 28859 34561 28871 34595
rect 28813 34555 28871 34561
rect 29089 34595 29147 34601
rect 29089 34561 29101 34595
rect 29135 34561 29147 34595
rect 29089 34555 29147 34561
rect 30101 34595 30159 34601
rect 30101 34561 30113 34595
rect 30147 34592 30159 34595
rect 30190 34592 30196 34604
rect 30147 34564 30196 34592
rect 30147 34561 30159 34564
rect 30101 34555 30159 34561
rect 25406 34524 25412 34536
rect 24627 34496 25268 34524
rect 25367 34496 25412 34524
rect 24627 34493 24639 34496
rect 24581 34487 24639 34493
rect 25406 34484 25412 34496
rect 25464 34484 25470 34536
rect 27985 34527 28043 34533
rect 27985 34493 27997 34527
rect 28031 34524 28043 34527
rect 28718 34524 28724 34536
rect 28031 34496 28724 34524
rect 28031 34493 28043 34496
rect 27985 34487 28043 34493
rect 28718 34484 28724 34496
rect 28776 34484 28782 34536
rect 17957 34459 18015 34465
rect 17957 34425 17969 34459
rect 18003 34425 18015 34459
rect 17957 34419 18015 34425
rect 18046 34416 18052 34468
rect 18104 34456 18110 34468
rect 18877 34459 18935 34465
rect 18877 34456 18889 34459
rect 18104 34428 18889 34456
rect 18104 34416 18110 34428
rect 18877 34425 18889 34428
rect 18923 34425 18935 34459
rect 18877 34419 18935 34425
rect 19058 34416 19064 34468
rect 19116 34456 19122 34468
rect 20990 34456 20996 34468
rect 19116 34428 20996 34456
rect 19116 34416 19122 34428
rect 20990 34416 20996 34428
rect 21048 34416 21054 34468
rect 25590 34456 25596 34468
rect 24688 34428 25596 34456
rect 17773 34391 17831 34397
rect 17773 34357 17785 34391
rect 17819 34388 17831 34391
rect 17862 34388 17868 34400
rect 17819 34360 17868 34388
rect 17819 34357 17831 34360
rect 17773 34351 17831 34357
rect 17862 34348 17868 34360
rect 17920 34348 17926 34400
rect 18138 34348 18144 34400
rect 18196 34388 18202 34400
rect 18417 34391 18475 34397
rect 18417 34388 18429 34391
rect 18196 34360 18429 34388
rect 18196 34348 18202 34360
rect 18417 34357 18429 34360
rect 18463 34357 18475 34391
rect 23566 34388 23572 34400
rect 23527 34360 23572 34388
rect 18417 34351 18475 34357
rect 23566 34348 23572 34360
rect 23624 34348 23630 34400
rect 24688 34397 24716 34428
rect 25590 34416 25596 34428
rect 25648 34416 25654 34468
rect 28828 34456 28856 34555
rect 30190 34552 30196 34564
rect 30248 34552 30254 34604
rect 31110 34592 31116 34604
rect 31071 34564 31116 34592
rect 31110 34552 31116 34564
rect 31168 34552 31174 34604
rect 31404 34601 31432 34632
rect 31389 34595 31447 34601
rect 31389 34561 31401 34595
rect 31435 34561 31447 34595
rect 48130 34592 48136 34604
rect 48091 34564 48136 34592
rect 31389 34555 31447 34561
rect 48130 34552 48136 34564
rect 48188 34552 48194 34604
rect 28994 34524 29000 34536
rect 28955 34496 29000 34524
rect 28994 34484 29000 34496
rect 29052 34484 29058 34536
rect 30006 34524 30012 34536
rect 29967 34496 30012 34524
rect 30006 34484 30012 34496
rect 30064 34484 30070 34536
rect 29362 34456 29368 34468
rect 28828 34428 29368 34456
rect 29362 34416 29368 34428
rect 29420 34416 29426 34468
rect 30469 34459 30527 34465
rect 30469 34425 30481 34459
rect 30515 34456 30527 34459
rect 31297 34459 31355 34465
rect 31297 34456 31309 34459
rect 30515 34428 31309 34456
rect 30515 34425 30527 34428
rect 30469 34419 30527 34425
rect 31297 34425 31309 34428
rect 31343 34425 31355 34459
rect 31297 34419 31355 34425
rect 24673 34391 24731 34397
rect 24673 34357 24685 34391
rect 24719 34357 24731 34391
rect 24854 34388 24860 34400
rect 24815 34360 24860 34388
rect 24673 34351 24731 34357
rect 24854 34348 24860 34360
rect 24912 34348 24918 34400
rect 25314 34388 25320 34400
rect 25275 34360 25320 34388
rect 25314 34348 25320 34360
rect 25372 34348 25378 34400
rect 28810 34388 28816 34400
rect 28771 34360 28816 34388
rect 28810 34348 28816 34360
rect 28868 34348 28874 34400
rect 47210 34348 47216 34400
rect 47268 34388 47274 34400
rect 47949 34391 48007 34397
rect 47949 34388 47961 34391
rect 47268 34360 47961 34388
rect 47268 34348 47274 34360
rect 47949 34357 47961 34360
rect 47995 34357 48007 34391
rect 47949 34351 48007 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 17313 34187 17371 34193
rect 17313 34153 17325 34187
rect 17359 34153 17371 34187
rect 17313 34147 17371 34153
rect 17328 34116 17356 34147
rect 17402 34144 17408 34196
rect 17460 34184 17466 34196
rect 17589 34187 17647 34193
rect 17589 34184 17601 34187
rect 17460 34156 17601 34184
rect 17460 34144 17466 34156
rect 17589 34153 17601 34156
rect 17635 34153 17647 34187
rect 18230 34184 18236 34196
rect 18191 34156 18236 34184
rect 17589 34147 17647 34153
rect 18230 34144 18236 34156
rect 18288 34144 18294 34196
rect 22005 34187 22063 34193
rect 22005 34153 22017 34187
rect 22051 34184 22063 34187
rect 22094 34184 22100 34196
rect 22051 34156 22100 34184
rect 22051 34153 22063 34156
rect 22005 34147 22063 34153
rect 22094 34144 22100 34156
rect 22152 34144 22158 34196
rect 22646 34184 22652 34196
rect 22607 34156 22652 34184
rect 22646 34144 22652 34156
rect 22704 34144 22710 34196
rect 23753 34187 23811 34193
rect 23753 34153 23765 34187
rect 23799 34184 23811 34187
rect 24854 34184 24860 34196
rect 23799 34156 24860 34184
rect 23799 34153 23811 34156
rect 23753 34147 23811 34153
rect 24854 34144 24860 34156
rect 24912 34144 24918 34196
rect 25222 34144 25228 34196
rect 25280 34184 25286 34196
rect 26145 34187 26203 34193
rect 26145 34184 26157 34187
rect 25280 34156 26157 34184
rect 25280 34144 25286 34156
rect 26145 34153 26157 34156
rect 26191 34153 26203 34187
rect 26145 34147 26203 34153
rect 27525 34187 27583 34193
rect 27525 34153 27537 34187
rect 27571 34184 27583 34187
rect 27614 34184 27620 34196
rect 27571 34156 27620 34184
rect 27571 34153 27583 34156
rect 27525 34147 27583 34153
rect 27614 34144 27620 34156
rect 27672 34144 27678 34196
rect 28166 34144 28172 34196
rect 28224 34184 28230 34196
rect 28537 34187 28595 34193
rect 28537 34184 28549 34187
rect 28224 34156 28549 34184
rect 28224 34144 28230 34156
rect 28537 34153 28549 34156
rect 28583 34153 28595 34187
rect 28537 34147 28595 34153
rect 30285 34187 30343 34193
rect 30285 34153 30297 34187
rect 30331 34184 30343 34187
rect 31110 34184 31116 34196
rect 30331 34156 31116 34184
rect 30331 34153 30343 34156
rect 30285 34147 30343 34153
rect 31110 34144 31116 34156
rect 31168 34144 31174 34196
rect 18248 34116 18276 34144
rect 24949 34119 25007 34125
rect 17328 34088 18276 34116
rect 19352 34088 21864 34116
rect 16206 34008 16212 34060
rect 16264 34048 16270 34060
rect 17313 34051 17371 34057
rect 16264 34020 16988 34048
rect 16264 34008 16270 34020
rect 1302 33940 1308 33992
rect 1360 33980 1366 33992
rect 1581 33983 1639 33989
rect 1581 33980 1593 33983
rect 1360 33952 1593 33980
rect 1360 33940 1366 33952
rect 1581 33949 1593 33952
rect 1627 33949 1639 33983
rect 14182 33980 14188 33992
rect 14143 33952 14188 33980
rect 1581 33943 1639 33949
rect 14182 33940 14188 33952
rect 14240 33940 14246 33992
rect 16390 33980 16396 33992
rect 16351 33952 16396 33980
rect 16390 33940 16396 33952
rect 16448 33940 16454 33992
rect 14458 33912 14464 33924
rect 14419 33884 14464 33912
rect 14458 33872 14464 33884
rect 14516 33872 14522 33924
rect 16485 33915 16543 33921
rect 16485 33912 16497 33915
rect 15686 33884 16497 33912
rect 16485 33881 16497 33884
rect 16531 33881 16543 33915
rect 16485 33875 16543 33881
rect 1397 33847 1455 33853
rect 1397 33813 1409 33847
rect 1443 33844 1455 33847
rect 1578 33844 1584 33856
rect 1443 33816 1584 33844
rect 1443 33813 1455 33816
rect 1397 33807 1455 33813
rect 1578 33804 1584 33816
rect 1636 33804 1642 33856
rect 15933 33847 15991 33853
rect 15933 33813 15945 33847
rect 15979 33844 15991 33847
rect 16390 33844 16396 33856
rect 15979 33816 16396 33844
rect 15979 33813 15991 33816
rect 15933 33807 15991 33813
rect 16390 33804 16396 33816
rect 16448 33804 16454 33856
rect 16960 33844 16988 34020
rect 17313 34017 17325 34051
rect 17359 34048 17371 34051
rect 17954 34048 17960 34060
rect 17359 34020 17960 34048
rect 17359 34017 17371 34020
rect 17313 34011 17371 34017
rect 17954 34008 17960 34020
rect 18012 34008 18018 34060
rect 18233 34051 18291 34057
rect 18233 34017 18245 34051
rect 18279 34048 18291 34051
rect 18414 34048 18420 34060
rect 18279 34020 18420 34048
rect 18279 34017 18291 34020
rect 18233 34011 18291 34017
rect 18414 34008 18420 34020
rect 18472 34048 18478 34060
rect 18966 34048 18972 34060
rect 18472 34020 18972 34048
rect 18472 34008 18478 34020
rect 18966 34008 18972 34020
rect 19024 34008 19030 34060
rect 17034 33940 17040 33992
rect 17092 33980 17098 33992
rect 17129 33983 17187 33989
rect 17129 33980 17141 33983
rect 17092 33952 17141 33980
rect 17092 33940 17098 33952
rect 17129 33949 17141 33952
rect 17175 33949 17187 33983
rect 17129 33943 17187 33949
rect 17218 33940 17224 33992
rect 17276 33980 17282 33992
rect 17405 33983 17463 33989
rect 17405 33980 17417 33983
rect 17276 33952 17417 33980
rect 17276 33940 17282 33952
rect 17405 33949 17417 33952
rect 17451 33949 17463 33983
rect 18046 33980 18052 33992
rect 18007 33952 18052 33980
rect 17405 33943 17463 33949
rect 17420 33912 17448 33943
rect 18046 33940 18052 33952
rect 18104 33940 18110 33992
rect 18325 33983 18383 33989
rect 18325 33949 18337 33983
rect 18371 33949 18383 33983
rect 18325 33943 18383 33949
rect 18340 33912 18368 33943
rect 19058 33940 19064 33992
rect 19116 33980 19122 33992
rect 19245 33983 19303 33989
rect 19245 33980 19257 33983
rect 19116 33952 19257 33980
rect 19116 33940 19122 33952
rect 19245 33949 19257 33952
rect 19291 33949 19303 33983
rect 19245 33943 19303 33949
rect 19352 33912 19380 34088
rect 20162 34008 20168 34060
rect 20220 34048 20226 34060
rect 21637 34051 21695 34057
rect 21637 34048 21649 34051
rect 20220 34020 21649 34048
rect 20220 34008 20226 34020
rect 21637 34017 21649 34020
rect 21683 34017 21695 34051
rect 21637 34011 21695 34017
rect 21836 34048 21864 34088
rect 22066 34088 24900 34116
rect 22066 34048 22094 34088
rect 21836 34020 22094 34048
rect 24872 34048 24900 34088
rect 24949 34085 24961 34119
rect 24995 34116 25007 34119
rect 25038 34116 25044 34128
rect 24995 34088 25044 34116
rect 24995 34085 25007 34088
rect 24949 34079 25007 34085
rect 25038 34076 25044 34088
rect 25096 34076 25102 34128
rect 27246 34116 27252 34128
rect 25516 34088 27252 34116
rect 25516 34048 25544 34088
rect 27246 34076 27252 34088
rect 27304 34076 27310 34128
rect 27982 34076 27988 34128
rect 28040 34076 28046 34128
rect 29086 34076 29092 34128
rect 29144 34116 29150 34128
rect 29144 34088 30696 34116
rect 29144 34076 29150 34088
rect 24872 34020 25544 34048
rect 21266 33980 21272 33992
rect 21227 33952 21272 33980
rect 21266 33940 21272 33952
rect 21324 33940 21330 33992
rect 21450 33980 21456 33992
rect 21376 33952 21456 33980
rect 20254 33912 20260 33924
rect 17420 33884 18368 33912
rect 18432 33884 19380 33912
rect 19444 33884 20260 33912
rect 18432 33844 18460 33884
rect 16960 33816 18460 33844
rect 18509 33847 18567 33853
rect 18509 33813 18521 33847
rect 18555 33844 18567 33847
rect 19334 33844 19340 33856
rect 18555 33816 19340 33844
rect 18555 33813 18567 33816
rect 18509 33807 18567 33813
rect 19334 33804 19340 33816
rect 19392 33804 19398 33856
rect 19444 33853 19472 33884
rect 20254 33872 20260 33884
rect 20312 33912 20318 33924
rect 21376 33912 21404 33952
rect 21450 33940 21456 33952
rect 21508 33940 21514 33992
rect 21836 33989 21864 34020
rect 25590 34008 25596 34060
rect 25648 34048 25654 34060
rect 25869 34051 25927 34057
rect 25869 34048 25881 34051
rect 25648 34020 25881 34048
rect 25648 34008 25654 34020
rect 25869 34017 25881 34020
rect 25915 34017 25927 34051
rect 27522 34048 27528 34060
rect 25869 34011 25927 34017
rect 26160 34020 27528 34048
rect 21545 33983 21603 33989
rect 21545 33949 21557 33983
rect 21591 33949 21603 33983
rect 21545 33943 21603 33949
rect 21821 33983 21879 33989
rect 21821 33949 21833 33983
rect 21867 33949 21879 33983
rect 21821 33943 21879 33949
rect 20312 33884 21404 33912
rect 21560 33912 21588 33943
rect 22278 33940 22284 33992
rect 22336 33980 22342 33992
rect 22557 33983 22615 33989
rect 22557 33980 22569 33983
rect 22336 33952 22569 33980
rect 22336 33940 22342 33952
rect 22557 33949 22569 33952
rect 22603 33980 22615 33983
rect 22738 33980 22744 33992
rect 22603 33952 22744 33980
rect 22603 33949 22615 33952
rect 22557 33943 22615 33949
rect 22738 33940 22744 33952
rect 22796 33940 22802 33992
rect 23566 33940 23572 33992
rect 23624 33980 23630 33992
rect 23845 33983 23903 33989
rect 23624 33952 23717 33980
rect 23624 33940 23630 33952
rect 23845 33949 23857 33983
rect 23891 33980 23903 33983
rect 24394 33980 24400 33992
rect 23891 33952 24400 33980
rect 23891 33949 23903 33952
rect 23845 33943 23903 33949
rect 24394 33940 24400 33952
rect 24452 33940 24458 33992
rect 24578 33983 24636 33989
rect 24578 33949 24590 33983
rect 24624 33980 24636 33983
rect 24762 33980 24768 33992
rect 24624 33952 24768 33980
rect 24624 33949 24636 33952
rect 24578 33943 24636 33949
rect 24762 33940 24768 33952
rect 24820 33940 24826 33992
rect 25038 33980 25044 33992
rect 24951 33952 25044 33980
rect 25038 33940 25044 33952
rect 25096 33980 25102 33992
rect 25096 33952 25636 33980
rect 25096 33940 25102 33952
rect 23584 33912 23612 33940
rect 25501 33915 25559 33921
rect 25501 33912 25513 33915
rect 21560 33884 23612 33912
rect 24412 33884 25513 33912
rect 20312 33872 20318 33884
rect 19429 33847 19487 33853
rect 19429 33813 19441 33847
rect 19475 33813 19487 33847
rect 19429 33807 19487 33813
rect 20990 33804 20996 33856
rect 21048 33844 21054 33856
rect 22462 33844 22468 33856
rect 21048 33816 22468 33844
rect 21048 33804 21054 33816
rect 22462 33804 22468 33816
rect 22520 33804 22526 33856
rect 22554 33804 22560 33856
rect 22612 33844 22618 33856
rect 24412 33853 24440 33884
rect 25501 33881 25513 33884
rect 25547 33881 25559 33915
rect 25608 33912 25636 33952
rect 25958 33940 25964 33992
rect 26016 33980 26022 33992
rect 26016 33952 26061 33980
rect 26016 33940 26022 33952
rect 26160 33912 26188 34020
rect 27522 34008 27528 34020
rect 27580 34008 27586 34060
rect 28000 34048 28028 34076
rect 27816 34020 28028 34048
rect 28905 34051 28963 34057
rect 26878 33980 26884 33992
rect 26839 33952 26884 33980
rect 26878 33940 26884 33952
rect 26936 33940 26942 33992
rect 26970 33940 26976 33992
rect 27028 33980 27034 33992
rect 27065 33983 27123 33989
rect 27065 33980 27077 33983
rect 27028 33952 27077 33980
rect 27028 33940 27034 33952
rect 27065 33949 27077 33952
rect 27111 33949 27123 33983
rect 27065 33943 27123 33949
rect 27614 33940 27620 33992
rect 27672 33980 27678 33992
rect 27816 33989 27844 34020
rect 28905 34017 28917 34051
rect 28951 34048 28963 34051
rect 29270 34048 29276 34060
rect 28951 34020 29276 34048
rect 28951 34017 28963 34020
rect 28905 34011 28963 34017
rect 29270 34008 29276 34020
rect 29328 34048 29334 34060
rect 30006 34048 30012 34060
rect 29328 34020 30012 34048
rect 29328 34008 29334 34020
rect 30006 34008 30012 34020
rect 30064 34008 30070 34060
rect 30190 34008 30196 34060
rect 30248 34048 30254 34060
rect 30248 34020 30604 34048
rect 30248 34008 30254 34020
rect 27709 33983 27767 33989
rect 27709 33980 27721 33983
rect 27672 33952 27721 33980
rect 27672 33940 27678 33952
rect 27709 33949 27721 33952
rect 27755 33949 27767 33983
rect 27709 33943 27767 33949
rect 27801 33983 27859 33989
rect 27801 33949 27813 33983
rect 27847 33949 27859 33983
rect 27801 33943 27859 33949
rect 27985 33983 28043 33989
rect 27985 33949 27997 33983
rect 28031 33949 28043 33983
rect 27985 33943 28043 33949
rect 28077 33983 28135 33989
rect 28077 33949 28089 33983
rect 28123 33980 28135 33983
rect 28258 33980 28264 33992
rect 28123 33952 28264 33980
rect 28123 33949 28135 33952
rect 28077 33943 28135 33949
rect 28000 33912 28028 33943
rect 28258 33940 28264 33952
rect 28316 33940 28322 33992
rect 28721 33983 28779 33989
rect 28721 33949 28733 33983
rect 28767 33980 28779 33983
rect 28810 33980 28816 33992
rect 28767 33952 28816 33980
rect 28767 33949 28779 33952
rect 28721 33943 28779 33949
rect 28810 33940 28816 33952
rect 28868 33940 28874 33992
rect 28994 33940 29000 33992
rect 29052 33980 29058 33992
rect 30208 33980 30236 34008
rect 30576 33989 30604 34020
rect 29052 33952 30236 33980
rect 30469 33983 30527 33989
rect 29052 33940 29058 33952
rect 30469 33949 30481 33983
rect 30515 33949 30527 33983
rect 30469 33943 30527 33949
rect 30561 33983 30619 33989
rect 30561 33949 30573 33983
rect 30607 33949 30619 33983
rect 30668 33980 30696 34088
rect 45554 34076 45560 34128
rect 45612 34116 45618 34128
rect 45612 34088 47440 34116
rect 45612 34076 45618 34088
rect 30745 34051 30803 34057
rect 30745 34017 30757 34051
rect 30791 34048 30803 34051
rect 44174 34048 44180 34060
rect 30791 34020 44180 34048
rect 30791 34017 30803 34020
rect 30745 34011 30803 34017
rect 44174 34008 44180 34020
rect 44232 34008 44238 34060
rect 47118 34048 47124 34060
rect 47079 34020 47124 34048
rect 47118 34008 47124 34020
rect 47176 34008 47182 34060
rect 47412 34057 47440 34088
rect 47397 34051 47455 34057
rect 47397 34017 47409 34051
rect 47443 34017 47455 34051
rect 47397 34011 47455 34017
rect 30837 33983 30895 33989
rect 30837 33980 30849 33983
rect 30668 33952 30849 33980
rect 30561 33943 30619 33949
rect 30837 33949 30849 33952
rect 30883 33949 30895 33983
rect 30837 33943 30895 33949
rect 25608 33884 26188 33912
rect 27080 33884 28028 33912
rect 25501 33875 25559 33881
rect 27080 33856 27108 33884
rect 23385 33847 23443 33853
rect 23385 33844 23397 33847
rect 22612 33816 23397 33844
rect 22612 33804 22618 33816
rect 23385 33813 23397 33816
rect 23431 33813 23443 33847
rect 23385 33807 23443 33813
rect 24397 33847 24455 33853
rect 24397 33813 24409 33847
rect 24443 33813 24455 33847
rect 24397 33807 24455 33813
rect 24581 33847 24639 33853
rect 24581 33813 24593 33847
rect 24627 33844 24639 33847
rect 24670 33844 24676 33856
rect 24627 33816 24676 33844
rect 24627 33813 24639 33816
rect 24581 33807 24639 33813
rect 24670 33804 24676 33816
rect 24728 33844 24734 33856
rect 25317 33847 25375 33853
rect 25317 33844 25329 33847
rect 24728 33816 25329 33844
rect 24728 33804 24734 33816
rect 25317 33813 25329 33816
rect 25363 33813 25375 33847
rect 25317 33807 25375 33813
rect 26973 33847 27031 33853
rect 26973 33813 26985 33847
rect 27019 33844 27031 33847
rect 27062 33844 27068 33856
rect 27019 33816 27068 33844
rect 27019 33813 27031 33816
rect 26973 33807 27031 33813
rect 27062 33804 27068 33816
rect 27120 33804 27126 33856
rect 27246 33804 27252 33856
rect 27304 33844 27310 33856
rect 30484 33844 30512 33943
rect 47210 33872 47216 33924
rect 47268 33912 47274 33924
rect 47268 33884 47313 33912
rect 47268 33872 47274 33884
rect 27304 33816 30512 33844
rect 27304 33804 27310 33816
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 14458 33600 14464 33652
rect 14516 33640 14522 33652
rect 15657 33643 15715 33649
rect 15657 33640 15669 33643
rect 14516 33612 15669 33640
rect 14516 33600 14522 33612
rect 15657 33609 15669 33612
rect 15703 33609 15715 33643
rect 15657 33603 15715 33609
rect 16390 33600 16396 33652
rect 16448 33640 16454 33652
rect 17681 33643 17739 33649
rect 17681 33640 17693 33643
rect 16448 33612 17693 33640
rect 16448 33600 16454 33612
rect 17681 33609 17693 33612
rect 17727 33640 17739 33643
rect 18138 33640 18144 33652
rect 17727 33612 18144 33640
rect 17727 33609 17739 33612
rect 17681 33603 17739 33609
rect 18138 33600 18144 33612
rect 18196 33600 18202 33652
rect 18969 33643 19027 33649
rect 18969 33640 18981 33643
rect 18524 33612 18981 33640
rect 16942 33572 16948 33584
rect 15856 33544 16948 33572
rect 15856 33513 15884 33544
rect 16942 33532 16948 33544
rect 17000 33532 17006 33584
rect 17402 33532 17408 33584
rect 17460 33572 17466 33584
rect 17460 33544 17816 33572
rect 17460 33532 17466 33544
rect 17788 33516 17816 33544
rect 15841 33507 15899 33513
rect 15841 33473 15853 33507
rect 15887 33473 15899 33507
rect 15841 33467 15899 33473
rect 16025 33507 16083 33513
rect 16025 33473 16037 33507
rect 16071 33473 16083 33507
rect 16025 33467 16083 33473
rect 16117 33507 16175 33513
rect 16117 33473 16129 33507
rect 16163 33504 16175 33507
rect 17313 33507 17371 33513
rect 17313 33504 17325 33507
rect 16163 33476 17325 33504
rect 16163 33473 16175 33476
rect 16117 33467 16175 33473
rect 17313 33473 17325 33476
rect 17359 33473 17371 33507
rect 17313 33467 17371 33473
rect 17497 33507 17555 33513
rect 17497 33473 17509 33507
rect 17543 33473 17555 33507
rect 17497 33467 17555 33473
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 1673 33439 1731 33445
rect 1673 33405 1685 33439
rect 1719 33436 1731 33439
rect 2498 33436 2504 33448
rect 1719 33408 2504 33436
rect 1719 33405 1731 33408
rect 1673 33399 1731 33405
rect 2498 33396 2504 33408
rect 2556 33396 2562 33448
rect 16040 33368 16068 33467
rect 17512 33436 17540 33467
rect 17770 33464 17776 33516
rect 17828 33504 17834 33516
rect 17828 33476 17921 33504
rect 17828 33464 17834 33476
rect 18524 33436 18552 33612
rect 18969 33609 18981 33612
rect 19015 33640 19027 33643
rect 19426 33640 19432 33652
rect 19015 33612 19432 33640
rect 19015 33609 19027 33612
rect 18969 33603 19027 33609
rect 19426 33600 19432 33612
rect 19484 33600 19490 33652
rect 19889 33643 19947 33649
rect 19889 33609 19901 33643
rect 19935 33640 19947 33643
rect 20714 33640 20720 33652
rect 19935 33612 20720 33640
rect 19935 33609 19947 33612
rect 19889 33603 19947 33609
rect 20714 33600 20720 33612
rect 20772 33600 20778 33652
rect 21266 33600 21272 33652
rect 21324 33640 21330 33652
rect 22373 33643 22431 33649
rect 22373 33640 22385 33643
rect 21324 33612 22385 33640
rect 21324 33600 21330 33612
rect 22373 33609 22385 33612
rect 22419 33609 22431 33643
rect 22373 33603 22431 33609
rect 22462 33600 22468 33652
rect 22520 33640 22526 33652
rect 22520 33612 25820 33640
rect 22520 33600 22526 33612
rect 18601 33575 18659 33581
rect 18601 33541 18613 33575
rect 18647 33541 18659 33575
rect 18601 33535 18659 33541
rect 18616 33504 18644 33535
rect 18690 33532 18696 33584
rect 18748 33572 18754 33584
rect 18801 33575 18859 33581
rect 18801 33572 18813 33575
rect 18748 33544 18813 33572
rect 18748 33532 18754 33544
rect 18801 33541 18813 33544
rect 18847 33541 18859 33575
rect 18801 33535 18859 33541
rect 19334 33532 19340 33584
rect 19392 33572 19398 33584
rect 23845 33575 23903 33581
rect 19392 33544 22094 33572
rect 19392 33532 19398 33544
rect 19702 33504 19708 33516
rect 18616 33476 19708 33504
rect 19702 33464 19708 33476
rect 19760 33464 19766 33516
rect 19797 33507 19855 33513
rect 19797 33473 19809 33507
rect 19843 33504 19855 33507
rect 19978 33504 19984 33516
rect 19843 33476 19984 33504
rect 19843 33473 19855 33476
rect 19797 33467 19855 33473
rect 19978 33464 19984 33476
rect 20036 33464 20042 33516
rect 20530 33464 20536 33516
rect 20588 33504 20594 33516
rect 20717 33507 20775 33513
rect 20717 33504 20729 33507
rect 20588 33476 20729 33504
rect 20588 33464 20594 33476
rect 20717 33473 20729 33476
rect 20763 33504 20775 33507
rect 21821 33507 21879 33513
rect 21821 33504 21833 33507
rect 20763 33476 21833 33504
rect 20763 33473 20775 33476
rect 20717 33467 20775 33473
rect 21821 33473 21833 33476
rect 21867 33473 21879 33507
rect 22066 33504 22094 33544
rect 23845 33541 23857 33575
rect 23891 33572 23903 33575
rect 24946 33572 24952 33584
rect 23891 33544 24952 33572
rect 23891 33541 23903 33544
rect 23845 33535 23903 33541
rect 24946 33532 24952 33544
rect 25004 33532 25010 33584
rect 25041 33575 25099 33581
rect 25041 33541 25053 33575
rect 25087 33572 25099 33575
rect 25314 33572 25320 33584
rect 25087 33544 25320 33572
rect 25087 33541 25099 33544
rect 25041 33535 25099 33541
rect 25314 33532 25320 33544
rect 25372 33532 25378 33584
rect 25792 33581 25820 33612
rect 25958 33600 25964 33652
rect 26016 33640 26022 33652
rect 27249 33643 27307 33649
rect 27249 33640 27261 33643
rect 26016 33612 27261 33640
rect 26016 33600 26022 33612
rect 27249 33609 27261 33612
rect 27295 33609 27307 33643
rect 27249 33603 27307 33609
rect 27614 33600 27620 33652
rect 27672 33640 27678 33652
rect 27798 33640 27804 33652
rect 27672 33612 27804 33640
rect 27672 33600 27678 33612
rect 27798 33600 27804 33612
rect 27856 33640 27862 33652
rect 28721 33643 28779 33649
rect 28721 33640 28733 33643
rect 27856 33612 28733 33640
rect 27856 33600 27862 33612
rect 28721 33609 28733 33612
rect 28767 33609 28779 33643
rect 28721 33603 28779 33609
rect 29549 33643 29607 33649
rect 29549 33609 29561 33643
rect 29595 33640 29607 33643
rect 30006 33640 30012 33652
rect 29595 33612 30012 33640
rect 29595 33609 29607 33612
rect 29549 33603 29607 33609
rect 30006 33600 30012 33612
rect 30064 33600 30070 33652
rect 25777 33575 25835 33581
rect 25777 33541 25789 33575
rect 25823 33541 25835 33575
rect 29270 33572 29276 33584
rect 25777 33535 25835 33541
rect 28368 33544 29276 33572
rect 22066 33476 23520 33504
rect 21821 33467 21879 33473
rect 18874 33436 18880 33448
rect 17512 33408 18552 33436
rect 18616 33408 18880 33436
rect 18616 33368 18644 33408
rect 18874 33396 18880 33408
rect 18932 33396 18938 33448
rect 20441 33439 20499 33445
rect 20441 33405 20453 33439
rect 20487 33405 20499 33439
rect 20441 33399 20499 33405
rect 22097 33439 22155 33445
rect 22097 33405 22109 33439
rect 22143 33436 22155 33439
rect 23382 33436 23388 33448
rect 22143 33408 23388 33436
rect 22143 33405 22155 33408
rect 22097 33399 22155 33405
rect 16040 33340 18644 33368
rect 20456 33368 20484 33399
rect 23382 33396 23388 33408
rect 23440 33396 23446 33448
rect 23492 33436 23520 33476
rect 23566 33464 23572 33516
rect 23624 33504 23630 33516
rect 24121 33507 24179 33513
rect 24121 33504 24133 33507
rect 23624 33476 24133 33504
rect 23624 33464 23630 33476
rect 24121 33473 24133 33476
rect 24167 33473 24179 33507
rect 24121 33467 24179 33473
rect 24857 33507 24915 33513
rect 24857 33473 24869 33507
rect 24903 33473 24915 33507
rect 24857 33467 24915 33473
rect 23937 33439 23995 33445
rect 23937 33436 23949 33439
rect 23492 33408 23949 33436
rect 23937 33405 23949 33408
rect 23983 33436 23995 33439
rect 24872 33436 24900 33467
rect 25590 33464 25596 33516
rect 25648 33504 25654 33516
rect 26973 33507 27031 33513
rect 26973 33504 26985 33507
rect 25648 33476 26985 33504
rect 25648 33464 25654 33476
rect 26973 33473 26985 33476
rect 27019 33473 27031 33507
rect 26973 33467 27031 33473
rect 27062 33464 27068 33516
rect 27120 33504 27126 33516
rect 28368 33513 28396 33544
rect 29270 33532 29276 33544
rect 29328 33532 29334 33584
rect 29362 33532 29368 33584
rect 29420 33572 29426 33584
rect 29420 33544 30236 33572
rect 29420 33532 29426 33544
rect 28353 33507 28411 33513
rect 27120 33476 27165 33504
rect 27120 33464 27126 33476
rect 28353 33473 28365 33507
rect 28399 33473 28411 33507
rect 28353 33467 28411 33473
rect 28537 33507 28595 33513
rect 28537 33473 28549 33507
rect 28583 33504 28595 33507
rect 28810 33504 28816 33516
rect 28583 33476 28816 33504
rect 28583 33473 28595 33476
rect 28537 33467 28595 33473
rect 28810 33464 28816 33476
rect 28868 33464 28874 33516
rect 30208 33513 30236 33544
rect 29181 33507 29239 33513
rect 29181 33504 29193 33507
rect 28920 33476 29193 33504
rect 25406 33436 25412 33448
rect 23983 33408 25412 33436
rect 23983 33405 23995 33408
rect 23937 33399 23995 33405
rect 25406 33396 25412 33408
rect 25464 33396 25470 33448
rect 25961 33439 26019 33445
rect 25961 33405 25973 33439
rect 26007 33436 26019 33439
rect 26878 33436 26884 33448
rect 26007 33408 26884 33436
rect 26007 33405 26019 33408
rect 25961 33399 26019 33405
rect 26878 33396 26884 33408
rect 26936 33436 26942 33448
rect 27246 33436 27252 33448
rect 26936 33408 27252 33436
rect 26936 33396 26942 33408
rect 27246 33396 27252 33408
rect 27304 33396 27310 33448
rect 21082 33368 21088 33380
rect 20456 33340 21088 33368
rect 21082 33328 21088 33340
rect 21140 33368 21146 33380
rect 24305 33371 24363 33377
rect 24305 33368 24317 33371
rect 21140 33340 24317 33368
rect 21140 33328 21146 33340
rect 24305 33337 24317 33340
rect 24351 33337 24363 33371
rect 24305 33331 24363 33337
rect 24394 33328 24400 33380
rect 24452 33368 24458 33380
rect 25225 33371 25283 33377
rect 25225 33368 25237 33371
rect 24452 33340 25237 33368
rect 24452 33328 24458 33340
rect 25225 33337 25237 33340
rect 25271 33368 25283 33371
rect 26970 33368 26976 33380
rect 25271 33340 26976 33368
rect 25271 33337 25283 33340
rect 25225 33331 25283 33337
rect 26970 33328 26976 33340
rect 27028 33368 27034 33380
rect 28920 33368 28948 33476
rect 29181 33473 29193 33476
rect 29227 33504 29239 33507
rect 30009 33507 30067 33513
rect 30009 33504 30021 33507
rect 29227 33476 30021 33504
rect 29227 33473 29239 33476
rect 29181 33467 29239 33473
rect 30009 33473 30021 33476
rect 30055 33473 30067 33507
rect 30009 33467 30067 33473
rect 30193 33507 30251 33513
rect 30193 33473 30205 33507
rect 30239 33504 30251 33507
rect 30282 33504 30288 33516
rect 30239 33476 30288 33504
rect 30239 33473 30251 33476
rect 30193 33467 30251 33473
rect 30282 33464 30288 33476
rect 30340 33464 30346 33516
rect 47854 33504 47860 33516
rect 47815 33476 47860 33504
rect 47854 33464 47860 33476
rect 47912 33464 47918 33516
rect 27028 33340 28948 33368
rect 27028 33328 27034 33340
rect 18785 33303 18843 33309
rect 18785 33269 18797 33303
rect 18831 33300 18843 33303
rect 21818 33300 21824 33312
rect 18831 33272 21824 33300
rect 18831 33269 18843 33272
rect 18785 33263 18843 33269
rect 21818 33260 21824 33272
rect 21876 33260 21882 33312
rect 22189 33303 22247 33309
rect 22189 33269 22201 33303
rect 22235 33300 22247 33303
rect 22554 33300 22560 33312
rect 22235 33272 22560 33300
rect 22235 33269 22247 33272
rect 22189 33263 22247 33269
rect 22554 33260 22560 33272
rect 22612 33260 22618 33312
rect 24121 33303 24179 33309
rect 24121 33269 24133 33303
rect 24167 33300 24179 33303
rect 24946 33300 24952 33312
rect 24167 33272 24952 33300
rect 24167 33269 24179 33272
rect 24121 33263 24179 33269
rect 24946 33260 24952 33272
rect 25004 33260 25010 33312
rect 28537 33303 28595 33309
rect 28537 33269 28549 33303
rect 28583 33300 28595 33303
rect 28994 33300 29000 33312
rect 28583 33272 29000 33300
rect 28583 33269 28595 33272
rect 28537 33263 28595 33269
rect 28994 33260 29000 33272
rect 29052 33260 29058 33312
rect 29638 33260 29644 33312
rect 29696 33300 29702 33312
rect 30101 33303 30159 33309
rect 30101 33300 30113 33303
rect 29696 33272 30113 33300
rect 29696 33260 29702 33272
rect 30101 33269 30113 33272
rect 30147 33269 30159 33303
rect 30101 33263 30159 33269
rect 41414 33260 41420 33312
rect 41472 33300 41478 33312
rect 48041 33303 48099 33309
rect 48041 33300 48053 33303
rect 41472 33272 48053 33300
rect 41472 33260 41478 33272
rect 48041 33269 48053 33272
rect 48087 33269 48099 33303
rect 48041 33263 48099 33269
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 16942 33096 16948 33108
rect 16903 33068 16948 33096
rect 16942 33056 16948 33068
rect 17000 33056 17006 33108
rect 17957 33099 18015 33105
rect 17957 33065 17969 33099
rect 18003 33096 18015 33099
rect 18690 33096 18696 33108
rect 18003 33068 18696 33096
rect 18003 33065 18015 33068
rect 17957 33059 18015 33065
rect 18690 33056 18696 33068
rect 18748 33056 18754 33108
rect 19242 33056 19248 33108
rect 19300 33096 19306 33108
rect 19300 33068 22416 33096
rect 19300 33056 19306 33068
rect 1486 33028 1492 33040
rect 1412 33000 1492 33028
rect 1412 32969 1440 33000
rect 1486 32988 1492 33000
rect 1544 32988 1550 33040
rect 22278 33028 22284 33040
rect 16684 33000 22284 33028
rect 1397 32963 1455 32969
rect 1397 32929 1409 32963
rect 1443 32929 1455 32963
rect 1578 32960 1584 32972
rect 1539 32932 1584 32960
rect 1397 32923 1455 32929
rect 1578 32920 1584 32932
rect 1636 32920 1642 32972
rect 16684 32904 16712 33000
rect 22278 32988 22284 33000
rect 22336 32988 22342 33040
rect 22388 33028 22416 33068
rect 22462 33056 22468 33108
rect 22520 33096 22526 33108
rect 23385 33099 23443 33105
rect 23385 33096 23397 33099
rect 22520 33068 23397 33096
rect 22520 33056 22526 33068
rect 23385 33065 23397 33068
rect 23431 33065 23443 33099
rect 23385 33059 23443 33065
rect 26142 33056 26148 33108
rect 26200 33096 26206 33108
rect 26697 33099 26755 33105
rect 26697 33096 26709 33099
rect 26200 33068 26709 33096
rect 26200 33056 26206 33068
rect 26697 33065 26709 33068
rect 26743 33065 26755 33099
rect 27890 33096 27896 33108
rect 27851 33068 27896 33096
rect 26697 33059 26755 33065
rect 27890 33056 27896 33068
rect 27948 33056 27954 33108
rect 23842 33028 23848 33040
rect 22388 33000 23848 33028
rect 23842 32988 23848 33000
rect 23900 33028 23906 33040
rect 24762 33028 24768 33040
rect 23900 33000 24768 33028
rect 23900 32988 23906 33000
rect 24762 32988 24768 33000
rect 24820 32988 24826 33040
rect 20364 32932 21496 32960
rect 16390 32892 16396 32904
rect 16351 32864 16396 32892
rect 16390 32852 16396 32864
rect 16448 32852 16454 32904
rect 16666 32892 16672 32904
rect 16579 32864 16672 32892
rect 16666 32852 16672 32864
rect 16724 32852 16730 32904
rect 16761 32895 16819 32901
rect 16761 32861 16773 32895
rect 16807 32892 16819 32895
rect 17678 32892 17684 32904
rect 16807 32864 17684 32892
rect 16807 32861 16819 32864
rect 16761 32855 16819 32861
rect 17678 32852 17684 32864
rect 17736 32852 17742 32904
rect 17770 32852 17776 32904
rect 17828 32892 17834 32904
rect 17957 32895 18015 32901
rect 17957 32892 17969 32895
rect 17828 32864 17969 32892
rect 17828 32852 17834 32864
rect 17957 32861 17969 32864
rect 18003 32861 18015 32895
rect 18138 32892 18144 32904
rect 18099 32864 18144 32892
rect 17957 32855 18015 32861
rect 18138 32852 18144 32864
rect 18196 32852 18202 32904
rect 3237 32827 3295 32833
rect 3237 32793 3249 32827
rect 3283 32824 3295 32827
rect 3970 32824 3976 32836
rect 3283 32796 3976 32824
rect 3283 32793 3295 32796
rect 3237 32787 3295 32793
rect 3970 32784 3976 32796
rect 4028 32784 4034 32836
rect 16577 32827 16635 32833
rect 16577 32793 16589 32827
rect 16623 32824 16635 32827
rect 16942 32824 16948 32836
rect 16623 32796 16948 32824
rect 16623 32793 16635 32796
rect 16577 32787 16635 32793
rect 16942 32784 16948 32796
rect 17000 32824 17006 32836
rect 18046 32824 18052 32836
rect 17000 32796 18052 32824
rect 17000 32784 17006 32796
rect 18046 32784 18052 32796
rect 18104 32784 18110 32836
rect 19702 32824 19708 32836
rect 19615 32796 19708 32824
rect 19702 32784 19708 32796
rect 19760 32824 19766 32836
rect 20162 32824 20168 32836
rect 19760 32796 20168 32824
rect 19760 32784 19766 32796
rect 20162 32784 20168 32796
rect 20220 32784 20226 32836
rect 19334 32716 19340 32768
rect 19392 32756 19398 32768
rect 19797 32759 19855 32765
rect 19797 32756 19809 32759
rect 19392 32728 19809 32756
rect 19392 32716 19398 32728
rect 19797 32725 19809 32728
rect 19843 32756 19855 32759
rect 20364 32756 20392 32932
rect 20717 32895 20775 32901
rect 20717 32861 20729 32895
rect 20763 32861 20775 32895
rect 20717 32855 20775 32861
rect 20732 32824 20760 32855
rect 21358 32824 21364 32836
rect 20732 32796 21364 32824
rect 21358 32784 21364 32796
rect 21416 32784 21422 32836
rect 21468 32824 21496 32932
rect 21726 32920 21732 32972
rect 21784 32960 21790 32972
rect 24302 32960 24308 32972
rect 21784 32932 24308 32960
rect 21784 32920 21790 32932
rect 24302 32920 24308 32932
rect 24360 32920 24366 32972
rect 26786 32920 26792 32972
rect 26844 32960 26850 32972
rect 27157 32963 27215 32969
rect 27157 32960 27169 32963
rect 26844 32932 27169 32960
rect 26844 32920 26850 32932
rect 27157 32929 27169 32932
rect 27203 32929 27215 32963
rect 27157 32923 27215 32929
rect 27890 32920 27896 32972
rect 27948 32960 27954 32972
rect 30561 32963 30619 32969
rect 30561 32960 30573 32963
rect 27948 32932 30573 32960
rect 27948 32920 27954 32932
rect 30561 32929 30573 32932
rect 30607 32929 30619 32963
rect 30561 32923 30619 32929
rect 21818 32852 21824 32904
rect 21876 32892 21882 32904
rect 22554 32892 22560 32904
rect 21876 32864 22560 32892
rect 21876 32852 21882 32864
rect 22554 32852 22560 32864
rect 22612 32852 22618 32904
rect 22649 32895 22707 32901
rect 22649 32861 22661 32895
rect 22695 32892 22707 32895
rect 23569 32895 23627 32901
rect 23569 32892 23581 32895
rect 22695 32864 23581 32892
rect 22695 32861 22707 32864
rect 22649 32855 22707 32861
rect 23569 32861 23581 32864
rect 23615 32861 23627 32895
rect 23569 32855 23627 32861
rect 23845 32895 23903 32901
rect 23845 32861 23857 32895
rect 23891 32892 23903 32895
rect 23934 32892 23940 32904
rect 23891 32864 23940 32892
rect 23891 32861 23903 32864
rect 23845 32855 23903 32861
rect 23584 32824 23612 32855
rect 23934 32852 23940 32864
rect 23992 32852 23998 32904
rect 26602 32852 26608 32904
rect 26660 32892 26666 32904
rect 26878 32892 26884 32904
rect 26660 32864 26884 32892
rect 26660 32852 26666 32864
rect 26878 32852 26884 32864
rect 26936 32852 26942 32904
rect 26973 32895 27031 32901
rect 26973 32861 26985 32895
rect 27019 32892 27031 32895
rect 27062 32892 27068 32904
rect 27019 32864 27068 32892
rect 27019 32861 27031 32864
rect 26973 32855 27031 32861
rect 27062 32852 27068 32864
rect 27120 32852 27126 32904
rect 27246 32892 27252 32904
rect 27207 32864 27252 32892
rect 27246 32852 27252 32864
rect 27304 32852 27310 32904
rect 29549 32895 29607 32901
rect 29549 32861 29561 32895
rect 29595 32892 29607 32895
rect 29638 32892 29644 32904
rect 29595 32864 29644 32892
rect 29595 32861 29607 32864
rect 29549 32855 29607 32861
rect 29638 32852 29644 32864
rect 29696 32852 29702 32904
rect 29733 32895 29791 32901
rect 29733 32861 29745 32895
rect 29779 32892 29791 32895
rect 30006 32892 30012 32904
rect 29779 32864 30012 32892
rect 29779 32861 29791 32864
rect 29733 32855 29791 32861
rect 30006 32852 30012 32864
rect 30064 32852 30070 32904
rect 46290 32892 46296 32904
rect 46251 32864 46296 32892
rect 46290 32852 46296 32864
rect 46348 32852 46354 32904
rect 25130 32824 25136 32836
rect 21468 32796 23520 32824
rect 23584 32796 25136 32824
rect 19843 32728 20392 32756
rect 19843 32725 19855 32728
rect 19797 32719 19855 32725
rect 20438 32716 20444 32768
rect 20496 32756 20502 32768
rect 20809 32759 20867 32765
rect 20809 32756 20821 32759
rect 20496 32728 20821 32756
rect 20496 32716 20502 32728
rect 20809 32725 20821 32728
rect 20855 32756 20867 32759
rect 22186 32756 22192 32768
rect 20855 32728 22192 32756
rect 20855 32725 20867 32728
rect 20809 32719 20867 32725
rect 22186 32716 22192 32728
rect 22244 32716 22250 32768
rect 22738 32756 22744 32768
rect 22699 32728 22744 32756
rect 22738 32716 22744 32728
rect 22796 32716 22802 32768
rect 23492 32756 23520 32796
rect 25130 32784 25136 32796
rect 25188 32784 25194 32836
rect 27338 32784 27344 32836
rect 27396 32824 27402 32836
rect 27801 32827 27859 32833
rect 27801 32824 27813 32827
rect 27396 32796 27813 32824
rect 27396 32784 27402 32796
rect 27801 32793 27813 32796
rect 27847 32793 27859 32827
rect 27801 32787 27859 32793
rect 30558 32784 30564 32836
rect 30616 32824 30622 32836
rect 30837 32827 30895 32833
rect 30837 32824 30849 32827
rect 30616 32796 30849 32824
rect 30616 32784 30622 32796
rect 30837 32793 30849 32796
rect 30883 32793 30895 32827
rect 30837 32787 30895 32793
rect 31386 32784 31392 32836
rect 31444 32784 31450 32836
rect 46477 32827 46535 32833
rect 46477 32793 46489 32827
rect 46523 32824 46535 32827
rect 47670 32824 47676 32836
rect 46523 32796 47676 32824
rect 46523 32793 46535 32796
rect 46477 32787 46535 32793
rect 47670 32784 47676 32796
rect 47728 32784 47734 32836
rect 48130 32824 48136 32836
rect 48091 32796 48136 32824
rect 48130 32784 48136 32796
rect 48188 32784 48194 32836
rect 23750 32756 23756 32768
rect 23492 32728 23756 32756
rect 23750 32716 23756 32728
rect 23808 32756 23814 32768
rect 24578 32756 24584 32768
rect 23808 32728 24584 32756
rect 23808 32716 23814 32728
rect 24578 32716 24584 32728
rect 24636 32716 24642 32768
rect 24762 32716 24768 32768
rect 24820 32756 24826 32768
rect 28166 32756 28172 32768
rect 24820 32728 28172 32756
rect 24820 32716 24826 32728
rect 28166 32716 28172 32728
rect 28224 32716 28230 32768
rect 29733 32759 29791 32765
rect 29733 32725 29745 32759
rect 29779 32756 29791 32759
rect 30006 32756 30012 32768
rect 29779 32728 30012 32756
rect 29779 32725 29791 32728
rect 29733 32719 29791 32725
rect 30006 32716 30012 32728
rect 30064 32716 30070 32768
rect 30282 32716 30288 32768
rect 30340 32756 30346 32768
rect 32309 32759 32367 32765
rect 32309 32756 32321 32759
rect 30340 32728 32321 32756
rect 30340 32716 30346 32728
rect 32309 32725 32321 32728
rect 32355 32725 32367 32759
rect 32309 32719 32367 32725
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 20162 32512 20168 32564
rect 20220 32552 20226 32564
rect 20220 32524 22508 32552
rect 20220 32512 20226 32524
rect 2498 32484 2504 32496
rect 2459 32456 2504 32484
rect 2498 32444 2504 32456
rect 2556 32444 2562 32496
rect 17034 32444 17040 32496
rect 17092 32484 17098 32496
rect 17092 32456 17816 32484
rect 17092 32444 17098 32456
rect 15286 32376 15292 32428
rect 15344 32416 15350 32428
rect 15381 32419 15439 32425
rect 15381 32416 15393 32419
rect 15344 32388 15393 32416
rect 15344 32376 15350 32388
rect 15381 32385 15393 32388
rect 15427 32385 15439 32419
rect 17126 32416 17132 32428
rect 17087 32388 17132 32416
rect 15381 32379 15439 32385
rect 17126 32376 17132 32388
rect 17184 32376 17190 32428
rect 17788 32425 17816 32456
rect 19978 32444 19984 32496
rect 20036 32484 20042 32496
rect 22097 32487 22155 32493
rect 22097 32484 22109 32487
rect 20036 32456 22109 32484
rect 20036 32444 20042 32456
rect 22097 32453 22109 32456
rect 22143 32453 22155 32487
rect 22480 32484 22508 32524
rect 22554 32512 22560 32564
rect 22612 32552 22618 32564
rect 23401 32555 23459 32561
rect 23401 32552 23413 32555
rect 22612 32524 23413 32552
rect 22612 32512 22618 32524
rect 23401 32521 23413 32524
rect 23447 32521 23459 32555
rect 24302 32552 24308 32564
rect 24263 32524 24308 32552
rect 23401 32515 23459 32521
rect 24302 32512 24308 32524
rect 24360 32552 24366 32564
rect 28350 32552 28356 32564
rect 24360 32524 28356 32552
rect 24360 32512 24366 32524
rect 28350 32512 28356 32524
rect 28408 32512 28414 32564
rect 30558 32552 30564 32564
rect 30519 32524 30564 32552
rect 30558 32512 30564 32524
rect 30616 32512 30622 32564
rect 31386 32552 31392 32564
rect 31347 32524 31392 32552
rect 31386 32512 31392 32524
rect 31444 32512 31450 32564
rect 47670 32552 47676 32564
rect 47631 32524 47676 32552
rect 47670 32512 47676 32524
rect 47728 32512 47734 32564
rect 23198 32484 23204 32496
rect 22480 32456 23204 32484
rect 22097 32447 22155 32453
rect 23198 32444 23204 32456
rect 23256 32444 23262 32496
rect 26053 32487 26111 32493
rect 26053 32484 26065 32487
rect 23400 32456 26065 32484
rect 23400 32428 23428 32456
rect 26053 32453 26065 32456
rect 26099 32453 26111 32487
rect 26418 32484 26424 32496
rect 26379 32456 26424 32484
rect 26053 32447 26111 32453
rect 26418 32444 26424 32456
rect 26476 32444 26482 32496
rect 30282 32484 30288 32496
rect 30243 32456 30288 32484
rect 30282 32444 30288 32456
rect 30340 32444 30346 32496
rect 31726 32456 35894 32484
rect 17773 32419 17831 32425
rect 17773 32385 17785 32419
rect 17819 32416 17831 32419
rect 17862 32416 17868 32428
rect 17819 32388 17868 32416
rect 17819 32385 17831 32388
rect 17773 32379 17831 32385
rect 17862 32376 17868 32388
rect 17920 32376 17926 32428
rect 17957 32419 18015 32425
rect 17957 32385 17969 32419
rect 18003 32416 18015 32419
rect 18230 32416 18236 32428
rect 18003 32388 18236 32416
rect 18003 32385 18015 32388
rect 17957 32379 18015 32385
rect 18230 32376 18236 32388
rect 18288 32376 18294 32428
rect 20438 32416 20444 32428
rect 20399 32388 20444 32416
rect 20438 32376 20444 32388
rect 20496 32376 20502 32428
rect 20530 32376 20536 32428
rect 20588 32416 20594 32428
rect 20901 32419 20959 32425
rect 20588 32388 20633 32416
rect 20588 32376 20594 32388
rect 20901 32385 20913 32419
rect 20947 32416 20959 32419
rect 21174 32416 21180 32428
rect 20947 32388 21180 32416
rect 20947 32385 20959 32388
rect 20901 32379 20959 32385
rect 21174 32376 21180 32388
rect 21232 32376 21238 32428
rect 21915 32419 21973 32425
rect 21915 32385 21927 32419
rect 21961 32385 21973 32419
rect 21915 32379 21973 32385
rect 2314 32348 2320 32360
rect 2275 32320 2320 32348
rect 2314 32308 2320 32320
rect 2372 32308 2378 32360
rect 3970 32348 3976 32360
rect 3931 32320 3976 32348
rect 3970 32308 3976 32320
rect 4028 32308 4034 32360
rect 20622 32348 20628 32360
rect 17972 32320 20628 32348
rect 17972 32292 18000 32320
rect 20622 32308 20628 32320
rect 20680 32308 20686 32360
rect 20714 32308 20720 32360
rect 20772 32348 20778 32360
rect 21726 32348 21732 32360
rect 20772 32320 20817 32348
rect 20916 32320 21732 32348
rect 20772 32308 20778 32320
rect 17954 32240 17960 32292
rect 18012 32240 18018 32292
rect 18046 32240 18052 32292
rect 18104 32280 18110 32292
rect 20916 32280 20944 32320
rect 21726 32308 21732 32320
rect 21784 32308 21790 32360
rect 21928 32348 21956 32379
rect 22370 32376 22376 32428
rect 22428 32416 22434 32428
rect 22557 32419 22615 32425
rect 22557 32416 22569 32419
rect 22428 32388 22569 32416
rect 22428 32376 22434 32388
rect 22557 32385 22569 32388
rect 22603 32385 22615 32419
rect 22557 32379 22615 32385
rect 23382 32376 23388 32428
rect 23440 32376 23446 32428
rect 24210 32416 24216 32428
rect 24171 32388 24216 32416
rect 24210 32376 24216 32388
rect 24268 32376 24274 32428
rect 24946 32416 24952 32428
rect 24907 32388 24952 32416
rect 24946 32376 24952 32388
rect 25004 32376 25010 32428
rect 27982 32376 27988 32428
rect 28040 32416 28046 32428
rect 28077 32419 28135 32425
rect 28077 32416 28089 32419
rect 28040 32388 28089 32416
rect 28040 32376 28046 32388
rect 28077 32385 28089 32388
rect 28123 32385 28135 32419
rect 29914 32416 29920 32428
rect 29875 32388 29920 32416
rect 28077 32379 28135 32385
rect 29914 32376 29920 32388
rect 29972 32376 29978 32428
rect 30006 32376 30012 32428
rect 30064 32416 30070 32428
rect 30190 32416 30196 32428
rect 30064 32388 30109 32416
rect 30151 32388 30196 32416
rect 30064 32376 30070 32388
rect 30190 32376 30196 32388
rect 30248 32376 30254 32428
rect 30382 32419 30440 32425
rect 30382 32416 30394 32419
rect 30300 32388 30394 32416
rect 25314 32348 25320 32360
rect 21928 32320 25320 32348
rect 25314 32308 25320 32320
rect 25372 32308 25378 32360
rect 26418 32308 26424 32360
rect 26476 32348 26482 32360
rect 28258 32348 28264 32360
rect 26476 32320 28264 32348
rect 26476 32308 26482 32320
rect 28258 32308 28264 32320
rect 28316 32308 28322 32360
rect 29730 32308 29736 32360
rect 29788 32348 29794 32360
rect 30300 32348 30328 32388
rect 30382 32385 30394 32388
rect 30428 32385 30440 32419
rect 31294 32416 31300 32428
rect 31255 32388 31300 32416
rect 30382 32379 30440 32385
rect 31294 32376 31300 32388
rect 31352 32376 31358 32428
rect 29788 32320 30328 32348
rect 29788 32308 29794 32320
rect 18104 32252 20944 32280
rect 18104 32240 18110 32252
rect 21450 32240 21456 32292
rect 21508 32280 21514 32292
rect 21508 32252 21956 32280
rect 21508 32240 21514 32252
rect 1394 32172 1400 32224
rect 1452 32212 1458 32224
rect 1857 32215 1915 32221
rect 1857 32212 1869 32215
rect 1452 32184 1869 32212
rect 1452 32172 1458 32184
rect 1857 32181 1869 32184
rect 1903 32181 1915 32215
rect 1857 32175 1915 32181
rect 15473 32215 15531 32221
rect 15473 32181 15485 32215
rect 15519 32212 15531 32215
rect 15654 32212 15660 32224
rect 15519 32184 15660 32212
rect 15519 32181 15531 32184
rect 15473 32175 15531 32181
rect 15654 32172 15660 32184
rect 15712 32172 15718 32224
rect 17218 32212 17224 32224
rect 17179 32184 17224 32212
rect 17218 32172 17224 32184
rect 17276 32172 17282 32224
rect 17773 32215 17831 32221
rect 17773 32181 17785 32215
rect 17819 32212 17831 32215
rect 18506 32212 18512 32224
rect 17819 32184 18512 32212
rect 17819 32181 17831 32184
rect 17773 32175 17831 32181
rect 18506 32172 18512 32184
rect 18564 32172 18570 32224
rect 20257 32215 20315 32221
rect 20257 32181 20269 32215
rect 20303 32212 20315 32215
rect 21818 32212 21824 32224
rect 20303 32184 21824 32212
rect 20303 32181 20315 32184
rect 20257 32175 20315 32181
rect 21818 32172 21824 32184
rect 21876 32172 21882 32224
rect 21928 32212 21956 32252
rect 23198 32240 23204 32292
rect 23256 32280 23262 32292
rect 31726 32280 31754 32456
rect 23256 32252 31754 32280
rect 35866 32280 35894 32456
rect 46290 32376 46296 32428
rect 46348 32416 46354 32428
rect 47029 32419 47087 32425
rect 47029 32416 47041 32419
rect 46348 32388 47041 32416
rect 46348 32376 46354 32388
rect 47029 32385 47041 32388
rect 47075 32385 47087 32419
rect 47029 32379 47087 32385
rect 47486 32376 47492 32428
rect 47544 32416 47550 32428
rect 47581 32419 47639 32425
rect 47581 32416 47593 32419
rect 47544 32388 47593 32416
rect 47544 32376 47550 32388
rect 47581 32385 47593 32388
rect 47627 32416 47639 32419
rect 47670 32416 47676 32428
rect 47627 32388 47676 32416
rect 47627 32385 47639 32388
rect 47581 32379 47639 32385
rect 47670 32376 47676 32388
rect 47728 32376 47734 32428
rect 41414 32280 41420 32292
rect 35866 32252 41420 32280
rect 23256 32240 23262 32252
rect 41414 32240 41420 32252
rect 41472 32240 41478 32292
rect 22649 32215 22707 32221
rect 22649 32212 22661 32215
rect 21928 32184 22661 32212
rect 22649 32181 22661 32184
rect 22695 32181 22707 32215
rect 22649 32175 22707 32181
rect 22738 32172 22744 32224
rect 22796 32212 22802 32224
rect 23385 32215 23443 32221
rect 23385 32212 23397 32215
rect 22796 32184 23397 32212
rect 22796 32172 22802 32184
rect 23385 32181 23397 32184
rect 23431 32181 23443 32215
rect 23566 32212 23572 32224
rect 23527 32184 23572 32212
rect 23385 32175 23443 32181
rect 23566 32172 23572 32184
rect 23624 32172 23630 32224
rect 25133 32215 25191 32221
rect 25133 32181 25145 32215
rect 25179 32212 25191 32215
rect 25222 32212 25228 32224
rect 25179 32184 25228 32212
rect 25179 32181 25191 32184
rect 25133 32175 25191 32181
rect 25222 32172 25228 32184
rect 25280 32212 25286 32224
rect 25682 32212 25688 32224
rect 25280 32184 25688 32212
rect 25280 32172 25286 32184
rect 25682 32172 25688 32184
rect 25740 32172 25746 32224
rect 28166 32212 28172 32224
rect 28079 32184 28172 32212
rect 28166 32172 28172 32184
rect 28224 32212 28230 32224
rect 29638 32212 29644 32224
rect 28224 32184 29644 32212
rect 28224 32172 28230 32184
rect 29638 32172 29644 32184
rect 29696 32172 29702 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 16025 32011 16083 32017
rect 16025 31977 16037 32011
rect 16071 32008 16083 32011
rect 17126 32008 17132 32020
rect 16071 31980 17132 32008
rect 16071 31977 16083 31980
rect 16025 31971 16083 31977
rect 17126 31968 17132 31980
rect 17184 31968 17190 32020
rect 17957 32011 18015 32017
rect 17957 31977 17969 32011
rect 18003 32008 18015 32011
rect 18322 32008 18328 32020
rect 18003 31980 18328 32008
rect 18003 31977 18015 31980
rect 17957 31971 18015 31977
rect 18322 31968 18328 31980
rect 18380 32008 18386 32020
rect 18601 32011 18659 32017
rect 18601 32008 18613 32011
rect 18380 31980 18613 32008
rect 18380 31968 18386 31980
rect 18601 31977 18613 31980
rect 18647 31977 18659 32011
rect 21358 32008 21364 32020
rect 21319 31980 21364 32008
rect 18601 31971 18659 31977
rect 21358 31968 21364 31980
rect 21416 31968 21422 32020
rect 21726 31968 21732 32020
rect 21784 32008 21790 32020
rect 23382 32008 23388 32020
rect 21784 31980 23388 32008
rect 21784 31968 21790 31980
rect 23382 31968 23388 31980
rect 23440 31968 23446 32020
rect 27341 32011 27399 32017
rect 27341 31977 27353 32011
rect 27387 32008 27399 32011
rect 27522 32008 27528 32020
rect 27387 31980 27528 32008
rect 27387 31977 27399 31980
rect 27341 31971 27399 31977
rect 27522 31968 27528 31980
rect 27580 31968 27586 32020
rect 29270 32008 29276 32020
rect 28184 31980 29276 32008
rect 28184 31952 28212 31980
rect 29270 31968 29276 31980
rect 29328 31968 29334 32020
rect 29914 31968 29920 32020
rect 29972 32008 29978 32020
rect 30009 32011 30067 32017
rect 30009 32008 30021 32011
rect 29972 31980 30021 32008
rect 29972 31968 29978 31980
rect 30009 31977 30021 31980
rect 30055 31977 30067 32011
rect 30009 31971 30067 31977
rect 16853 31943 16911 31949
rect 16853 31940 16865 31943
rect 15764 31912 16865 31940
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 1854 31872 1860 31884
rect 1815 31844 1860 31872
rect 1854 31832 1860 31844
rect 1912 31832 1918 31884
rect 14182 31832 14188 31884
rect 14240 31872 14246 31884
rect 14277 31875 14335 31881
rect 14277 31872 14289 31875
rect 14240 31844 14289 31872
rect 14240 31832 14246 31844
rect 14277 31841 14289 31844
rect 14323 31841 14335 31875
rect 14277 31835 14335 31841
rect 14553 31875 14611 31881
rect 14553 31841 14565 31875
rect 14599 31872 14611 31875
rect 15764 31872 15792 31912
rect 16853 31909 16865 31912
rect 16899 31909 16911 31943
rect 17405 31943 17463 31949
rect 17405 31940 17417 31943
rect 16853 31903 16911 31909
rect 16960 31912 17417 31940
rect 16758 31872 16764 31884
rect 14599 31844 15792 31872
rect 16719 31844 16764 31872
rect 14599 31841 14611 31844
rect 14553 31835 14611 31841
rect 16758 31832 16764 31844
rect 16816 31832 16822 31884
rect 16960 31881 16988 31912
rect 17405 31909 17417 31912
rect 17451 31909 17463 31943
rect 17405 31903 17463 31909
rect 17512 31912 18736 31940
rect 16945 31875 17003 31881
rect 16945 31841 16957 31875
rect 16991 31841 17003 31875
rect 17218 31872 17224 31884
rect 16945 31835 17003 31841
rect 17052 31844 17224 31872
rect 15654 31764 15660 31816
rect 15712 31764 15718 31816
rect 16669 31807 16727 31813
rect 16669 31773 16681 31807
rect 16715 31804 16727 31807
rect 17052 31804 17080 31844
rect 17218 31832 17224 31844
rect 17276 31872 17282 31884
rect 17512 31872 17540 31912
rect 17276 31844 17540 31872
rect 17276 31832 17282 31844
rect 17954 31832 17960 31884
rect 18012 31872 18018 31884
rect 18049 31875 18107 31881
rect 18049 31872 18061 31875
rect 18012 31844 18061 31872
rect 18012 31832 18018 31844
rect 18049 31841 18061 31844
rect 18095 31841 18107 31875
rect 18049 31835 18107 31841
rect 16715 31776 16749 31804
rect 16960 31776 17080 31804
rect 17586 31807 17644 31813
rect 16715 31773 16727 31776
rect 16669 31767 16727 31773
rect 1578 31736 1584 31748
rect 1539 31708 1584 31736
rect 1578 31696 1584 31708
rect 1636 31696 1642 31748
rect 16684 31736 16712 31767
rect 16960 31736 16988 31776
rect 17586 31773 17598 31807
rect 17632 31804 17644 31807
rect 18506 31804 18512 31816
rect 17632 31776 17908 31804
rect 18467 31776 18512 31804
rect 17632 31773 17644 31776
rect 17586 31767 17644 31773
rect 17880 31770 17908 31776
rect 17880 31742 18000 31770
rect 18506 31764 18512 31776
rect 18564 31764 18570 31816
rect 18708 31813 18736 31912
rect 25590 31900 25596 31952
rect 25648 31940 25654 31952
rect 25685 31943 25743 31949
rect 25685 31940 25697 31943
rect 25648 31912 25697 31940
rect 25648 31900 25654 31912
rect 25685 31909 25697 31912
rect 25731 31940 25743 31943
rect 28166 31940 28172 31952
rect 25731 31912 28172 31940
rect 25731 31909 25743 31912
rect 25685 31903 25743 31909
rect 28166 31900 28172 31912
rect 28224 31900 28230 31952
rect 28350 31900 28356 31952
rect 28408 31940 28414 31952
rect 29730 31940 29736 31952
rect 28408 31912 29736 31940
rect 28408 31900 28414 31912
rect 29730 31900 29736 31912
rect 29788 31940 29794 31952
rect 30190 31940 30196 31952
rect 29788 31912 30196 31940
rect 29788 31900 29794 31912
rect 30190 31900 30196 31912
rect 30248 31900 30254 31952
rect 19889 31875 19947 31881
rect 19889 31841 19901 31875
rect 19935 31872 19947 31875
rect 21818 31872 21824 31884
rect 19935 31844 21128 31872
rect 21779 31844 21824 31872
rect 19935 31841 19947 31844
rect 19889 31835 19947 31841
rect 18693 31807 18751 31813
rect 18693 31773 18705 31807
rect 18739 31773 18751 31807
rect 18693 31767 18751 31773
rect 19426 31764 19432 31816
rect 19484 31804 19490 31816
rect 19613 31807 19671 31813
rect 19613 31804 19625 31807
rect 19484 31776 19625 31804
rect 19484 31764 19490 31776
rect 19613 31773 19625 31776
rect 19659 31773 19671 31807
rect 21100 31804 21128 31844
rect 21818 31832 21824 31844
rect 21876 31832 21882 31884
rect 23569 31875 23627 31881
rect 23569 31841 23581 31875
rect 23615 31872 23627 31875
rect 24762 31872 24768 31884
rect 23615 31844 24768 31872
rect 23615 31841 23627 31844
rect 23569 31835 23627 31841
rect 24762 31832 24768 31844
rect 24820 31832 24826 31884
rect 46014 31872 46020 31884
rect 28092 31844 46020 31872
rect 22005 31807 22063 31813
rect 22005 31804 22017 31807
rect 21100 31776 22017 31804
rect 19613 31767 19671 31773
rect 22005 31773 22017 31776
rect 22051 31773 22063 31807
rect 22186 31804 22192 31816
rect 22147 31776 22192 31804
rect 22005 31767 22063 31773
rect 22186 31764 22192 31776
rect 22244 31764 22250 31816
rect 22281 31807 22339 31813
rect 22281 31773 22293 31807
rect 22327 31804 22339 31807
rect 22327 31776 22361 31804
rect 22327 31773 22339 31776
rect 22281 31767 22339 31773
rect 16684 31708 16988 31736
rect 17972 31736 18000 31742
rect 18322 31736 18328 31748
rect 17972 31708 18328 31736
rect 18322 31696 18328 31708
rect 18380 31736 18386 31748
rect 19242 31736 19248 31748
rect 18380 31708 19248 31736
rect 18380 31696 18386 31708
rect 19242 31696 19248 31708
rect 19300 31696 19306 31748
rect 21450 31736 21456 31748
rect 21114 31708 21456 31736
rect 21450 31696 21456 31708
rect 21508 31696 21514 31748
rect 22094 31696 22100 31748
rect 22152 31736 22158 31748
rect 22296 31736 22324 31767
rect 23198 31764 23204 31816
rect 23256 31804 23262 31816
rect 23477 31807 23535 31813
rect 23477 31804 23489 31807
rect 23256 31776 23489 31804
rect 23256 31764 23262 31776
rect 23477 31773 23489 31776
rect 23523 31773 23535 31807
rect 23477 31767 23535 31773
rect 24026 31764 24032 31816
rect 24084 31804 24090 31816
rect 24397 31807 24455 31813
rect 24397 31804 24409 31807
rect 24084 31776 24409 31804
rect 24084 31764 24090 31776
rect 24397 31773 24409 31776
rect 24443 31773 24455 31807
rect 24578 31804 24584 31816
rect 24539 31776 24584 31804
rect 24397 31767 24455 31773
rect 24578 31764 24584 31776
rect 24636 31764 24642 31816
rect 24854 31764 24860 31816
rect 24912 31804 24918 31816
rect 24949 31807 25007 31813
rect 24949 31804 24961 31807
rect 24912 31776 24961 31804
rect 24912 31764 24918 31776
rect 24949 31773 24961 31776
rect 24995 31804 25007 31807
rect 25501 31807 25559 31813
rect 25501 31804 25513 31807
rect 24995 31776 25513 31804
rect 24995 31773 25007 31776
rect 24949 31767 25007 31773
rect 25501 31773 25513 31776
rect 25547 31804 25559 31807
rect 25547 31776 25581 31804
rect 25547 31773 25559 31776
rect 25501 31767 25559 31773
rect 22152 31708 22324 31736
rect 25516 31736 25544 31767
rect 26142 31764 26148 31816
rect 26200 31804 26206 31816
rect 28092 31813 28120 31844
rect 46014 31832 46020 31844
rect 46072 31832 46078 31884
rect 47581 31875 47639 31881
rect 47581 31872 47593 31875
rect 46584 31844 47593 31872
rect 26237 31807 26295 31813
rect 26237 31804 26249 31807
rect 26200 31776 26249 31804
rect 26200 31764 26206 31776
rect 26237 31773 26249 31776
rect 26283 31804 26295 31807
rect 27249 31807 27307 31813
rect 27249 31804 27261 31807
rect 26283 31776 27261 31804
rect 26283 31773 26295 31776
rect 26237 31767 26295 31773
rect 27249 31773 27261 31776
rect 27295 31773 27307 31807
rect 27249 31767 27307 31773
rect 28077 31807 28135 31813
rect 28077 31773 28089 31807
rect 28123 31773 28135 31807
rect 28077 31767 28135 31773
rect 28166 31764 28172 31816
rect 28224 31804 28230 31816
rect 28350 31804 28356 31816
rect 28224 31776 28269 31804
rect 28311 31776 28356 31804
rect 28224 31764 28230 31776
rect 28350 31764 28356 31776
rect 28408 31764 28414 31816
rect 28445 31807 28503 31813
rect 28445 31773 28457 31807
rect 28491 31804 28503 31807
rect 28810 31804 28816 31816
rect 28491 31776 28816 31804
rect 28491 31773 28503 31776
rect 28445 31767 28503 31773
rect 28810 31764 28816 31776
rect 28868 31764 28874 31816
rect 29638 31804 29644 31816
rect 29599 31776 29644 31804
rect 29638 31764 29644 31776
rect 29696 31764 29702 31816
rect 29822 31804 29828 31816
rect 29783 31776 29828 31804
rect 29822 31764 29828 31776
rect 29880 31764 29886 31816
rect 44174 31764 44180 31816
rect 44232 31804 44238 31816
rect 46584 31804 46612 31844
rect 47581 31841 47593 31844
rect 47627 31841 47639 31875
rect 47581 31835 47639 31841
rect 47302 31804 47308 31816
rect 44232 31776 46612 31804
rect 47263 31776 47308 31804
rect 44232 31764 44238 31776
rect 47302 31764 47308 31776
rect 47360 31764 47366 31816
rect 27982 31736 27988 31748
rect 25516 31708 27988 31736
rect 22152 31696 22158 31708
rect 27982 31696 27988 31708
rect 28040 31696 28046 31748
rect 17402 31628 17408 31680
rect 17460 31668 17466 31680
rect 17589 31671 17647 31677
rect 17589 31668 17601 31671
rect 17460 31640 17601 31668
rect 17460 31628 17466 31640
rect 17589 31637 17601 31640
rect 17635 31637 17647 31671
rect 17589 31631 17647 31637
rect 17862 31628 17868 31680
rect 17920 31668 17926 31680
rect 18230 31668 18236 31680
rect 17920 31640 18236 31668
rect 17920 31628 17926 31640
rect 18230 31628 18236 31640
rect 18288 31628 18294 31680
rect 21174 31628 21180 31680
rect 21232 31668 21238 31680
rect 23474 31668 23480 31680
rect 21232 31640 23480 31668
rect 21232 31628 21238 31640
rect 23474 31628 23480 31640
rect 23532 31668 23538 31680
rect 24210 31668 24216 31680
rect 23532 31640 24216 31668
rect 23532 31628 23538 31640
rect 24210 31628 24216 31640
rect 24268 31668 24274 31680
rect 24581 31671 24639 31677
rect 24581 31668 24593 31671
rect 24268 31640 24593 31668
rect 24268 31628 24274 31640
rect 24581 31637 24593 31640
rect 24627 31637 24639 31671
rect 26418 31668 26424 31680
rect 26379 31640 26424 31668
rect 24581 31631 24639 31637
rect 26418 31628 26424 31640
rect 26476 31628 26482 31680
rect 27706 31628 27712 31680
rect 27764 31668 27770 31680
rect 27893 31671 27951 31677
rect 27893 31668 27905 31671
rect 27764 31640 27905 31668
rect 27764 31628 27770 31640
rect 27893 31637 27905 31640
rect 27939 31637 27951 31671
rect 27893 31631 27951 31637
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1578 31424 1584 31476
rect 1636 31464 1642 31476
rect 2225 31467 2283 31473
rect 2225 31464 2237 31467
rect 1636 31436 2237 31464
rect 1636 31424 1642 31436
rect 2225 31433 2237 31436
rect 2271 31433 2283 31467
rect 2225 31427 2283 31433
rect 15470 31424 15476 31476
rect 15528 31464 15534 31476
rect 19337 31467 19395 31473
rect 19337 31464 19349 31467
rect 15528 31436 19349 31464
rect 15528 31424 15534 31436
rect 19337 31433 19349 31436
rect 19383 31433 19395 31467
rect 19337 31427 19395 31433
rect 21269 31467 21327 31473
rect 21269 31433 21281 31467
rect 21315 31464 21327 31467
rect 21315 31436 22140 31464
rect 21315 31433 21327 31436
rect 21269 31427 21327 31433
rect 15654 31356 15660 31408
rect 15712 31356 15718 31408
rect 18874 31396 18880 31408
rect 17236 31368 18880 31396
rect 2130 31328 2136 31340
rect 2091 31300 2136 31328
rect 2130 31288 2136 31300
rect 2188 31328 2194 31340
rect 2406 31328 2412 31340
rect 2188 31300 2412 31328
rect 2188 31288 2194 31300
rect 2406 31288 2412 31300
rect 2464 31288 2470 31340
rect 16758 31288 16764 31340
rect 16816 31328 16822 31340
rect 16853 31331 16911 31337
rect 16853 31328 16865 31331
rect 16816 31300 16865 31328
rect 16816 31288 16822 31300
rect 16853 31297 16865 31300
rect 16899 31297 16911 31331
rect 16853 31291 16911 31297
rect 16945 31331 17003 31337
rect 16945 31297 16957 31331
rect 16991 31328 17003 31331
rect 17126 31328 17132 31340
rect 16991 31300 17132 31328
rect 16991 31297 17003 31300
rect 16945 31291 17003 31297
rect 14369 31263 14427 31269
rect 14369 31229 14381 31263
rect 14415 31229 14427 31263
rect 14369 31223 14427 31229
rect 14645 31263 14703 31269
rect 14645 31229 14657 31263
rect 14691 31260 14703 31263
rect 16669 31263 16727 31269
rect 16669 31260 16681 31263
rect 14691 31232 16681 31260
rect 14691 31229 14703 31232
rect 14645 31223 14703 31229
rect 16669 31229 16681 31232
rect 16715 31229 16727 31263
rect 16868 31260 16896 31291
rect 17126 31288 17132 31300
rect 17184 31288 17190 31340
rect 17236 31337 17264 31368
rect 18874 31356 18880 31368
rect 18932 31356 18938 31408
rect 20901 31399 20959 31405
rect 20901 31365 20913 31399
rect 20947 31396 20959 31399
rect 22002 31396 22008 31408
rect 20947 31368 22008 31396
rect 20947 31365 20959 31368
rect 20901 31359 20959 31365
rect 22002 31356 22008 31368
rect 22060 31356 22066 31408
rect 22112 31405 22140 31436
rect 24578 31424 24584 31476
rect 24636 31464 24642 31476
rect 24762 31464 24768 31476
rect 24636 31436 24768 31464
rect 24636 31424 24642 31436
rect 24762 31424 24768 31436
rect 24820 31424 24826 31476
rect 30190 31424 30196 31476
rect 30248 31424 30254 31476
rect 22097 31399 22155 31405
rect 22097 31365 22109 31399
rect 22143 31365 22155 31399
rect 22097 31359 22155 31365
rect 22738 31356 22744 31408
rect 22796 31356 22802 31408
rect 27982 31356 27988 31408
rect 28040 31396 28046 31408
rect 28353 31399 28411 31405
rect 28040 31368 28212 31396
rect 28040 31356 28046 31368
rect 17221 31331 17279 31337
rect 17221 31297 17233 31331
rect 17267 31297 17279 31331
rect 17221 31291 17279 31297
rect 17957 31331 18015 31337
rect 17957 31297 17969 31331
rect 18003 31328 18015 31331
rect 18506 31328 18512 31340
rect 18003 31300 18512 31328
rect 18003 31297 18015 31300
rect 17957 31291 18015 31297
rect 18506 31288 18512 31300
rect 18564 31288 18570 31340
rect 19153 31331 19211 31337
rect 19153 31297 19165 31331
rect 19199 31328 19211 31331
rect 20622 31328 20628 31340
rect 19199 31300 20300 31328
rect 20583 31300 20628 31328
rect 19199 31297 19211 31300
rect 19153 31291 19211 31297
rect 17773 31263 17831 31269
rect 17773 31260 17785 31263
rect 16868 31232 17785 31260
rect 16669 31223 16727 31229
rect 17773 31229 17785 31232
rect 17819 31229 17831 31263
rect 18046 31260 18052 31272
rect 18007 31232 18052 31260
rect 17773 31223 17831 31229
rect 14384 31124 14412 31223
rect 18046 31220 18052 31232
rect 18104 31220 18110 31272
rect 18141 31263 18199 31269
rect 18141 31229 18153 31263
rect 18187 31229 18199 31263
rect 18141 31223 18199 31229
rect 18233 31263 18291 31269
rect 18233 31229 18245 31263
rect 18279 31260 18291 31263
rect 18322 31260 18328 31272
rect 18279 31232 18328 31260
rect 18279 31229 18291 31232
rect 18233 31223 18291 31229
rect 16117 31195 16175 31201
rect 16117 31161 16129 31195
rect 16163 31192 16175 31195
rect 17954 31192 17960 31204
rect 16163 31164 17960 31192
rect 16163 31161 16175 31164
rect 16117 31155 16175 31161
rect 17954 31152 17960 31164
rect 18012 31152 18018 31204
rect 18156 31192 18184 31223
rect 18322 31220 18328 31232
rect 18380 31220 18386 31272
rect 19334 31220 19340 31272
rect 19392 31220 19398 31272
rect 19352 31192 19380 31220
rect 18156 31164 19380 31192
rect 20272 31192 20300 31300
rect 20622 31288 20628 31300
rect 20680 31288 20686 31340
rect 20714 31288 20720 31340
rect 20772 31328 20778 31340
rect 20990 31328 20996 31340
rect 20772 31300 20817 31328
rect 20951 31300 20996 31328
rect 20772 31288 20778 31300
rect 20990 31288 20996 31300
rect 21048 31288 21054 31340
rect 21090 31331 21148 31337
rect 21090 31297 21102 31331
rect 21136 31297 21148 31331
rect 21090 31291 21148 31297
rect 24029 31331 24087 31337
rect 24029 31297 24041 31331
rect 24075 31328 24087 31331
rect 24762 31328 24768 31340
rect 24075 31300 24768 31328
rect 24075 31297 24087 31300
rect 24029 31291 24087 31297
rect 20346 31220 20352 31272
rect 20404 31260 20410 31272
rect 21100 31260 21128 31291
rect 24762 31288 24768 31300
rect 24820 31288 24826 31340
rect 27341 31331 27399 31337
rect 27341 31297 27353 31331
rect 27387 31328 27399 31331
rect 27706 31328 27712 31340
rect 27387 31300 27712 31328
rect 27387 31297 27399 31300
rect 27341 31291 27399 31297
rect 27706 31288 27712 31300
rect 27764 31288 27770 31340
rect 28074 31328 28080 31340
rect 28035 31300 28080 31328
rect 28074 31288 28080 31300
rect 28132 31288 28138 31340
rect 28184 31328 28212 31368
rect 28353 31365 28365 31399
rect 28399 31396 28411 31399
rect 28399 31368 29132 31396
rect 28399 31365 28411 31368
rect 28353 31359 28411 31365
rect 28813 31331 28871 31337
rect 28813 31328 28825 31331
rect 28184 31300 28825 31328
rect 28813 31297 28825 31300
rect 28859 31297 28871 31331
rect 28813 31291 28871 31297
rect 28902 31288 28908 31340
rect 28960 31328 28966 31340
rect 29104 31337 29132 31368
rect 29270 31356 29276 31408
rect 29328 31396 29334 31408
rect 30101 31399 30159 31405
rect 29328 31368 30052 31396
rect 29328 31356 29334 31368
rect 28997 31331 29055 31337
rect 28997 31328 29009 31331
rect 28960 31300 29009 31328
rect 28960 31288 28966 31300
rect 28997 31297 29009 31300
rect 29043 31297 29055 31331
rect 28997 31291 29055 31297
rect 29089 31331 29147 31337
rect 29089 31297 29101 31331
rect 29135 31297 29147 31331
rect 29089 31291 29147 31297
rect 29917 31331 29975 31337
rect 29917 31297 29929 31331
rect 29963 31297 29975 31331
rect 30024 31328 30052 31368
rect 30101 31365 30113 31399
rect 30147 31396 30159 31399
rect 30208 31396 30236 31424
rect 30147 31368 30236 31396
rect 30147 31365 30159 31368
rect 30101 31359 30159 31365
rect 30193 31331 30251 31337
rect 30193 31328 30205 31331
rect 30024 31300 30205 31328
rect 29917 31291 29975 31297
rect 30193 31297 30205 31300
rect 30239 31297 30251 31331
rect 30193 31291 30251 31297
rect 30285 31331 30343 31337
rect 30285 31297 30297 31331
rect 30331 31297 30343 31331
rect 30285 31291 30343 31297
rect 20404 31232 21128 31260
rect 21821 31263 21879 31269
rect 20404 31220 20410 31232
rect 21821 31229 21833 31263
rect 21867 31229 21879 31263
rect 21821 31223 21879 31229
rect 21726 31192 21732 31204
rect 20272 31164 21732 31192
rect 21726 31152 21732 31164
rect 21784 31152 21790 31204
rect 16022 31124 16028 31136
rect 14384 31096 16028 31124
rect 16022 31084 16028 31096
rect 16080 31084 16086 31136
rect 16758 31084 16764 31136
rect 16816 31124 16822 31136
rect 17129 31127 17187 31133
rect 17129 31124 17141 31127
rect 16816 31096 17141 31124
rect 16816 31084 16822 31096
rect 17129 31093 17141 31096
rect 17175 31093 17187 31127
rect 17129 31087 17187 31093
rect 18046 31084 18052 31136
rect 18104 31124 18110 31136
rect 20898 31124 20904 31136
rect 18104 31096 20904 31124
rect 18104 31084 18110 31096
rect 20898 31084 20904 31096
rect 20956 31084 20962 31136
rect 21836 31124 21864 31223
rect 25314 31220 25320 31272
rect 25372 31260 25378 31272
rect 25774 31260 25780 31272
rect 25372 31232 25780 31260
rect 25372 31220 25378 31232
rect 25774 31220 25780 31232
rect 25832 31220 25838 31272
rect 27617 31263 27675 31269
rect 27617 31229 27629 31263
rect 27663 31260 27675 31263
rect 28166 31260 28172 31272
rect 27663 31232 28172 31260
rect 27663 31229 27675 31232
rect 27617 31223 27675 31229
rect 28166 31220 28172 31232
rect 28224 31260 28230 31272
rect 28353 31263 28411 31269
rect 28353 31260 28365 31263
rect 28224 31232 28365 31260
rect 28224 31220 28230 31232
rect 28353 31229 28365 31232
rect 28399 31229 28411 31263
rect 28353 31223 28411 31229
rect 27062 31192 27068 31204
rect 23492 31164 27068 31192
rect 23492 31124 23520 31164
rect 27062 31152 27068 31164
rect 27120 31152 27126 31204
rect 28810 31192 28816 31204
rect 28771 31164 28816 31192
rect 28810 31152 28816 31164
rect 28868 31152 28874 31204
rect 29932 31192 29960 31291
rect 30098 31220 30104 31272
rect 30156 31260 30162 31272
rect 30300 31260 30328 31291
rect 30156 31232 30328 31260
rect 30156 31220 30162 31232
rect 29932 31164 30144 31192
rect 30116 31136 30144 31164
rect 21836 31096 23520 31124
rect 23566 31084 23572 31136
rect 23624 31124 23630 31136
rect 23624 31096 23669 31124
rect 23624 31084 23630 31096
rect 26694 31084 26700 31136
rect 26752 31124 26758 31136
rect 27157 31127 27215 31133
rect 27157 31124 27169 31127
rect 26752 31096 27169 31124
rect 26752 31084 26758 31096
rect 27157 31093 27169 31096
rect 27203 31093 27215 31127
rect 27157 31087 27215 31093
rect 27525 31127 27583 31133
rect 27525 31093 27537 31127
rect 27571 31124 27583 31127
rect 27614 31124 27620 31136
rect 27571 31096 27620 31124
rect 27571 31093 27583 31096
rect 27525 31087 27583 31093
rect 27614 31084 27620 31096
rect 27672 31084 27678 31136
rect 28169 31127 28227 31133
rect 28169 31093 28181 31127
rect 28215 31124 28227 31127
rect 28626 31124 28632 31136
rect 28215 31096 28632 31124
rect 28215 31093 28227 31096
rect 28169 31087 28227 31093
rect 28626 31084 28632 31096
rect 28684 31084 28690 31136
rect 30098 31084 30104 31136
rect 30156 31084 30162 31136
rect 30469 31127 30527 31133
rect 30469 31093 30481 31127
rect 30515 31124 30527 31127
rect 31018 31124 31024 31136
rect 30515 31096 31024 31124
rect 30515 31093 30527 31096
rect 30469 31087 30527 31093
rect 31018 31084 31024 31096
rect 31076 31084 31082 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 15565 30923 15623 30929
rect 15565 30889 15577 30923
rect 15611 30920 15623 30923
rect 15654 30920 15660 30932
rect 15611 30892 15660 30920
rect 15611 30889 15623 30892
rect 15565 30883 15623 30889
rect 15654 30880 15660 30892
rect 15712 30880 15718 30932
rect 17126 30880 17132 30932
rect 17184 30920 17190 30932
rect 17865 30923 17923 30929
rect 17865 30920 17877 30923
rect 17184 30892 17877 30920
rect 17184 30880 17190 30892
rect 17865 30889 17877 30892
rect 17911 30889 17923 30923
rect 17865 30883 17923 30889
rect 20990 30880 20996 30932
rect 21048 30920 21054 30932
rect 22738 30920 22744 30932
rect 21048 30892 22094 30920
rect 22699 30892 22744 30920
rect 21048 30880 21054 30892
rect 20622 30812 20628 30864
rect 20680 30852 20686 30864
rect 21729 30855 21787 30861
rect 21729 30852 21741 30855
rect 20680 30824 21741 30852
rect 20680 30812 20686 30824
rect 21729 30821 21741 30824
rect 21775 30821 21787 30855
rect 21729 30815 21787 30821
rect 21821 30855 21879 30861
rect 21821 30821 21833 30855
rect 21867 30852 21879 30855
rect 21910 30852 21916 30864
rect 21867 30824 21916 30852
rect 21867 30821 21879 30824
rect 21821 30815 21879 30821
rect 21910 30812 21916 30824
rect 21968 30812 21974 30864
rect 22066 30852 22094 30892
rect 22738 30880 22744 30892
rect 22796 30880 22802 30932
rect 27062 30880 27068 30932
rect 27120 30920 27126 30932
rect 28166 30920 28172 30932
rect 27120 30892 28028 30920
rect 28127 30892 28172 30920
rect 27120 30880 27126 30892
rect 23106 30852 23112 30864
rect 22066 30824 23112 30852
rect 23106 30812 23112 30824
rect 23164 30852 23170 30864
rect 23845 30855 23903 30861
rect 23845 30852 23857 30855
rect 23164 30824 23857 30852
rect 23164 30812 23170 30824
rect 23845 30821 23857 30824
rect 23891 30821 23903 30855
rect 23845 30815 23903 30821
rect 14550 30744 14556 30796
rect 14608 30784 14614 30796
rect 20809 30787 20867 30793
rect 14608 30756 17264 30784
rect 14608 30744 14614 30756
rect 15470 30716 15476 30728
rect 15431 30688 15476 30716
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 16850 30716 16856 30728
rect 16811 30688 16856 30716
rect 16850 30676 16856 30688
rect 16908 30676 16914 30728
rect 16942 30676 16948 30728
rect 17000 30716 17006 30728
rect 17236 30725 17264 30756
rect 20809 30753 20821 30787
rect 20855 30784 20867 30787
rect 22094 30784 22100 30796
rect 20855 30756 22100 30784
rect 20855 30753 20867 30756
rect 20809 30747 20867 30753
rect 22094 30744 22100 30756
rect 22152 30744 22158 30796
rect 24854 30784 24860 30796
rect 23676 30756 24860 30784
rect 17037 30719 17095 30725
rect 17037 30716 17049 30719
rect 17000 30688 17049 30716
rect 17000 30676 17006 30688
rect 17037 30685 17049 30688
rect 17083 30685 17095 30719
rect 17037 30679 17095 30685
rect 17221 30719 17279 30725
rect 17221 30685 17233 30719
rect 17267 30685 17279 30719
rect 17221 30679 17279 30685
rect 17954 30676 17960 30728
rect 18012 30716 18018 30728
rect 18049 30719 18107 30725
rect 18049 30716 18061 30719
rect 18012 30688 18061 30716
rect 18012 30676 18018 30688
rect 18049 30685 18061 30688
rect 18095 30685 18107 30719
rect 18230 30716 18236 30728
rect 18191 30688 18236 30716
rect 18049 30679 18107 30685
rect 18230 30676 18236 30688
rect 18288 30676 18294 30728
rect 18325 30719 18383 30725
rect 18325 30685 18337 30719
rect 18371 30716 18383 30719
rect 20993 30719 21051 30725
rect 20993 30716 21005 30719
rect 18371 30688 21005 30716
rect 18371 30685 18383 30688
rect 18325 30679 18383 30685
rect 20993 30685 21005 30688
rect 21039 30716 21051 30719
rect 21174 30716 21180 30728
rect 21039 30688 21180 30716
rect 21039 30685 21051 30688
rect 20993 30679 21051 30685
rect 21174 30676 21180 30688
rect 21232 30676 21238 30728
rect 21269 30719 21327 30725
rect 21269 30685 21281 30719
rect 21315 30716 21327 30719
rect 21729 30719 21787 30725
rect 21729 30716 21741 30719
rect 21315 30688 21741 30716
rect 21315 30685 21327 30688
rect 21269 30679 21327 30685
rect 21729 30685 21741 30688
rect 21775 30716 21787 30719
rect 21910 30716 21916 30728
rect 21775 30688 21916 30716
rect 21775 30685 21787 30688
rect 21729 30679 21787 30685
rect 21910 30676 21916 30688
rect 21968 30676 21974 30728
rect 22370 30676 22376 30728
rect 22428 30716 22434 30728
rect 23676 30725 23704 30756
rect 24854 30744 24860 30756
rect 24912 30784 24918 30796
rect 25225 30787 25283 30793
rect 25225 30784 25237 30787
rect 24912 30756 25237 30784
rect 24912 30744 24918 30756
rect 25225 30753 25237 30756
rect 25271 30753 25283 30787
rect 25225 30747 25283 30753
rect 26421 30787 26479 30793
rect 26421 30753 26433 30787
rect 26467 30784 26479 30787
rect 27890 30784 27896 30796
rect 26467 30756 27896 30784
rect 26467 30753 26479 30756
rect 26421 30747 26479 30753
rect 27890 30744 27896 30756
rect 27948 30744 27954 30796
rect 28000 30784 28028 30892
rect 28166 30880 28172 30892
rect 28224 30880 28230 30932
rect 28810 30920 28816 30932
rect 28771 30892 28816 30920
rect 28810 30880 28816 30892
rect 28868 30880 28874 30932
rect 28074 30812 28080 30864
rect 28132 30852 28138 30864
rect 28828 30852 28856 30880
rect 28132 30824 28856 30852
rect 28132 30812 28138 30824
rect 30193 30787 30251 30793
rect 30193 30784 30205 30787
rect 28000 30756 30205 30784
rect 30193 30753 30205 30756
rect 30239 30753 30251 30787
rect 30193 30747 30251 30753
rect 22649 30719 22707 30725
rect 22649 30716 22661 30719
rect 22428 30688 22661 30716
rect 22428 30676 22434 30688
rect 22649 30685 22661 30688
rect 22695 30685 22707 30719
rect 22649 30679 22707 30685
rect 23661 30719 23719 30725
rect 23661 30685 23673 30719
rect 23707 30685 23719 30719
rect 23661 30679 23719 30685
rect 24949 30719 25007 30725
rect 24949 30685 24961 30719
rect 24995 30716 25007 30719
rect 25130 30716 25136 30728
rect 24995 30688 25136 30716
rect 24995 30685 25007 30688
rect 24949 30679 25007 30685
rect 25130 30676 25136 30688
rect 25188 30676 25194 30728
rect 28626 30716 28632 30728
rect 28587 30688 28632 30716
rect 28626 30676 28632 30688
rect 28684 30676 28690 30728
rect 28721 30719 28779 30725
rect 28721 30685 28733 30719
rect 28767 30685 28779 30719
rect 28721 30679 28779 30685
rect 16666 30608 16672 30660
rect 16724 30648 16730 30660
rect 17129 30651 17187 30657
rect 17129 30648 17141 30651
rect 16724 30620 17141 30648
rect 16724 30608 16730 30620
rect 17129 30617 17141 30620
rect 17175 30617 17187 30651
rect 17129 30611 17187 30617
rect 20714 30608 20720 30660
rect 20772 30648 20778 30660
rect 22002 30648 22008 30660
rect 20772 30620 22008 30648
rect 20772 30608 20778 30620
rect 22002 30608 22008 30620
rect 22060 30648 22066 30660
rect 23566 30648 23572 30660
rect 22060 30620 23572 30648
rect 22060 30608 22066 30620
rect 23566 30608 23572 30620
rect 23624 30608 23630 30660
rect 26694 30648 26700 30660
rect 26655 30620 26700 30648
rect 26694 30608 26700 30620
rect 26752 30608 26758 30660
rect 27706 30608 27712 30660
rect 27764 30608 27770 30660
rect 28166 30608 28172 30660
rect 28224 30648 28230 30660
rect 28736 30648 28764 30679
rect 30466 30648 30472 30660
rect 28224 30620 28764 30648
rect 30427 30620 30472 30648
rect 28224 30608 28230 30620
rect 30466 30608 30472 30620
rect 30524 30608 30530 30660
rect 31110 30608 31116 30660
rect 31168 30608 31174 30660
rect 17310 30540 17316 30592
rect 17368 30580 17374 30592
rect 17405 30583 17463 30589
rect 17405 30580 17417 30583
rect 17368 30552 17417 30580
rect 17368 30540 17374 30552
rect 17405 30549 17417 30552
rect 17451 30549 17463 30583
rect 17405 30543 17463 30549
rect 21177 30583 21235 30589
rect 21177 30549 21189 30583
rect 21223 30580 21235 30583
rect 21266 30580 21272 30592
rect 21223 30552 21272 30580
rect 21223 30549 21235 30552
rect 21177 30543 21235 30549
rect 21266 30540 21272 30552
rect 21324 30540 21330 30592
rect 28350 30540 28356 30592
rect 28408 30580 28414 30592
rect 28902 30580 28908 30592
rect 28408 30552 28908 30580
rect 28408 30540 28414 30552
rect 28902 30540 28908 30552
rect 28960 30580 28966 30592
rect 28997 30583 29055 30589
rect 28997 30580 29009 30583
rect 28960 30552 29009 30580
rect 28960 30540 28966 30552
rect 28997 30549 29009 30552
rect 29043 30549 29055 30583
rect 28997 30543 29055 30549
rect 30098 30540 30104 30592
rect 30156 30580 30162 30592
rect 31941 30583 31999 30589
rect 31941 30580 31953 30583
rect 30156 30552 31953 30580
rect 30156 30540 30162 30552
rect 31941 30549 31953 30552
rect 31987 30549 31999 30583
rect 31941 30543 31999 30549
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 24581 30379 24639 30385
rect 21836 30348 22324 30376
rect 19705 30311 19763 30317
rect 19705 30277 19717 30311
rect 19751 30308 19763 30311
rect 19978 30308 19984 30320
rect 19751 30280 19984 30308
rect 19751 30277 19763 30280
rect 19705 30271 19763 30277
rect 19978 30268 19984 30280
rect 20036 30268 20042 30320
rect 20530 30308 20536 30320
rect 20491 30280 20536 30308
rect 20530 30268 20536 30280
rect 20588 30268 20594 30320
rect 20714 30268 20720 30320
rect 20772 30308 20778 30320
rect 21836 30308 21864 30348
rect 20772 30280 21864 30308
rect 20772 30268 20778 30280
rect 21910 30268 21916 30320
rect 21968 30308 21974 30320
rect 22189 30311 22247 30317
rect 22189 30308 22201 30311
rect 21968 30280 22201 30308
rect 21968 30268 21974 30280
rect 22189 30277 22201 30280
rect 22235 30277 22247 30311
rect 22296 30308 22324 30348
rect 24581 30345 24593 30379
rect 24627 30345 24639 30379
rect 26142 30376 26148 30388
rect 24581 30339 24639 30345
rect 25700 30348 26148 30376
rect 23842 30308 23848 30320
rect 22296 30280 23848 30308
rect 22189 30271 22247 30277
rect 23842 30268 23848 30280
rect 23900 30268 23906 30320
rect 24596 30308 24624 30339
rect 25590 30308 25596 30320
rect 24504 30280 25596 30308
rect 20346 30240 20352 30252
rect 20307 30212 20352 30240
rect 20346 30200 20352 30212
rect 20404 30200 20410 30252
rect 20548 30240 20576 30268
rect 21821 30243 21879 30249
rect 21821 30240 21833 30243
rect 20548 30212 21833 30240
rect 21821 30209 21833 30212
rect 21867 30209 21879 30243
rect 21821 30203 21879 30209
rect 22005 30243 22063 30249
rect 22005 30209 22017 30243
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 23753 30243 23811 30249
rect 23753 30209 23765 30243
rect 23799 30240 23811 30243
rect 24504 30240 24532 30280
rect 25590 30268 25596 30280
rect 25648 30308 25654 30320
rect 25700 30308 25728 30348
rect 26142 30336 26148 30348
rect 26200 30336 26206 30388
rect 28626 30376 28632 30388
rect 27632 30348 28632 30376
rect 25648 30280 25728 30308
rect 25648 30268 25654 30280
rect 25774 30268 25780 30320
rect 25832 30308 25838 30320
rect 27065 30311 27123 30317
rect 27065 30308 27077 30311
rect 25832 30280 27077 30308
rect 25832 30268 25838 30280
rect 27065 30277 27077 30280
rect 27111 30277 27123 30311
rect 27065 30271 27123 30277
rect 27249 30311 27307 30317
rect 27249 30277 27261 30311
rect 27295 30308 27307 30311
rect 27338 30308 27344 30320
rect 27295 30280 27344 30308
rect 27295 30277 27307 30280
rect 27249 30271 27307 30277
rect 27338 30268 27344 30280
rect 27396 30268 27402 30320
rect 23799 30212 24532 30240
rect 23799 30209 23811 30212
rect 23753 30203 23811 30209
rect 12986 30172 12992 30184
rect 12947 30144 12992 30172
rect 12986 30132 12992 30144
rect 13044 30132 13050 30184
rect 13173 30175 13231 30181
rect 13173 30141 13185 30175
rect 13219 30172 13231 30175
rect 13446 30172 13452 30184
rect 13219 30144 13452 30172
rect 13219 30141 13231 30144
rect 13173 30135 13231 30141
rect 13446 30132 13452 30144
rect 13504 30132 13510 30184
rect 13541 30175 13599 30181
rect 13541 30141 13553 30175
rect 13587 30141 13599 30175
rect 13541 30135 13599 30141
rect 8294 30064 8300 30116
rect 8352 30104 8358 30116
rect 13556 30104 13584 30135
rect 18230 30132 18236 30184
rect 18288 30172 18294 30184
rect 21266 30172 21272 30184
rect 18288 30144 21272 30172
rect 18288 30132 18294 30144
rect 21266 30132 21272 30144
rect 21324 30132 21330 30184
rect 21358 30132 21364 30184
rect 21416 30172 21422 30184
rect 22020 30172 22048 30203
rect 24578 30200 24584 30252
rect 24636 30240 24642 30252
rect 24765 30243 24823 30249
rect 24765 30240 24777 30243
rect 24636 30212 24777 30240
rect 24636 30200 24642 30212
rect 24765 30209 24777 30212
rect 24811 30209 24823 30243
rect 24765 30203 24823 30209
rect 25409 30243 25467 30249
rect 25409 30209 25421 30243
rect 25455 30209 25467 30243
rect 25409 30203 25467 30209
rect 24397 30175 24455 30181
rect 24397 30172 24409 30175
rect 21416 30144 22048 30172
rect 23032 30144 24409 30172
rect 21416 30132 21422 30144
rect 8352 30076 13584 30104
rect 8352 30064 8358 30076
rect 18966 30064 18972 30116
rect 19024 30104 19030 30116
rect 19024 30076 20852 30104
rect 19024 30064 19030 30076
rect 19426 29996 19432 30048
rect 19484 30036 19490 30048
rect 19797 30039 19855 30045
rect 19797 30036 19809 30039
rect 19484 30008 19809 30036
rect 19484 29996 19490 30008
rect 19797 30005 19809 30008
rect 19843 30005 19855 30039
rect 19797 29999 19855 30005
rect 20438 29996 20444 30048
rect 20496 30036 20502 30048
rect 20717 30039 20775 30045
rect 20717 30036 20729 30039
rect 20496 30008 20729 30036
rect 20496 29996 20502 30008
rect 20717 30005 20729 30008
rect 20763 30005 20775 30039
rect 20824 30036 20852 30076
rect 21542 30064 21548 30116
rect 21600 30104 21606 30116
rect 22554 30104 22560 30116
rect 21600 30076 22560 30104
rect 21600 30064 21606 30076
rect 22554 30064 22560 30076
rect 22612 30104 22618 30116
rect 23032 30104 23060 30144
rect 24397 30141 24409 30144
rect 24443 30141 24455 30175
rect 24397 30135 24455 30141
rect 25424 30104 25452 30203
rect 25498 30200 25504 30252
rect 25556 30240 25562 30252
rect 25685 30243 25743 30249
rect 25685 30240 25697 30243
rect 25556 30212 25697 30240
rect 25556 30200 25562 30212
rect 25685 30209 25697 30212
rect 25731 30240 25743 30243
rect 27632 30240 27660 30348
rect 28626 30336 28632 30348
rect 28684 30336 28690 30388
rect 30466 30336 30472 30388
rect 30524 30376 30530 30388
rect 30837 30379 30895 30385
rect 30837 30376 30849 30379
rect 30524 30348 30849 30376
rect 30524 30336 30530 30348
rect 30837 30345 30849 30348
rect 30883 30345 30895 30379
rect 30837 30339 30895 30345
rect 27709 30311 27767 30317
rect 27709 30277 27721 30311
rect 27755 30308 27767 30311
rect 28166 30308 28172 30320
rect 27755 30280 28172 30308
rect 27755 30277 27767 30280
rect 27709 30271 27767 30277
rect 28166 30268 28172 30280
rect 28224 30268 28230 30320
rect 29089 30311 29147 30317
rect 29089 30277 29101 30311
rect 29135 30308 29147 30311
rect 30374 30308 30380 30320
rect 29135 30280 30380 30308
rect 29135 30277 29147 30280
rect 29089 30271 29147 30277
rect 30374 30268 30380 30280
rect 30432 30268 30438 30320
rect 31205 30311 31263 30317
rect 31205 30308 31217 30311
rect 30484 30280 31217 30308
rect 25731 30212 27660 30240
rect 27893 30243 27951 30249
rect 25731 30209 25743 30212
rect 25685 30203 25743 30209
rect 27893 30209 27905 30243
rect 27939 30240 27951 30243
rect 28534 30240 28540 30252
rect 27939 30212 28540 30240
rect 27939 30209 27951 30212
rect 27893 30203 27951 30209
rect 28534 30200 28540 30212
rect 28592 30200 28598 30252
rect 28810 30200 28816 30252
rect 28868 30240 28874 30252
rect 28905 30243 28963 30249
rect 28905 30240 28917 30243
rect 28868 30212 28917 30240
rect 28868 30200 28874 30212
rect 28905 30209 28917 30212
rect 28951 30240 28963 30243
rect 30009 30243 30067 30249
rect 30009 30240 30021 30243
rect 28951 30212 30021 30240
rect 28951 30209 28963 30212
rect 28905 30203 28963 30209
rect 30009 30209 30021 30212
rect 30055 30240 30067 30243
rect 30098 30240 30104 30252
rect 30055 30212 30104 30240
rect 30055 30209 30067 30212
rect 30009 30203 30067 30209
rect 30098 30200 30104 30212
rect 30156 30200 30162 30252
rect 30282 30200 30288 30252
rect 30340 30240 30346 30252
rect 30484 30240 30512 30280
rect 31205 30277 31217 30280
rect 31251 30277 31263 30311
rect 31205 30271 31263 30277
rect 31018 30240 31024 30252
rect 30340 30212 30512 30240
rect 30979 30212 31024 30240
rect 30340 30200 30346 30212
rect 31018 30200 31024 30212
rect 31076 30200 31082 30252
rect 31297 30243 31355 30249
rect 31297 30209 31309 30243
rect 31343 30209 31355 30243
rect 31297 30203 31355 30209
rect 25593 30175 25651 30181
rect 25593 30141 25605 30175
rect 25639 30172 25651 30175
rect 26050 30172 26056 30184
rect 25639 30144 26056 30172
rect 25639 30141 25651 30144
rect 25593 30135 25651 30141
rect 26050 30132 26056 30144
rect 26108 30172 26114 30184
rect 29273 30175 29331 30181
rect 29273 30172 29285 30175
rect 26108 30144 29285 30172
rect 26108 30132 26114 30144
rect 29273 30141 29285 30144
rect 29319 30141 29331 30175
rect 29273 30135 29331 30141
rect 29917 30175 29975 30181
rect 29917 30141 29929 30175
rect 29963 30141 29975 30175
rect 31312 30172 31340 30203
rect 29917 30135 29975 30141
rect 30392 30144 31340 30172
rect 26142 30104 26148 30116
rect 22612 30076 23060 30104
rect 23768 30076 25452 30104
rect 25700 30076 26148 30104
rect 22612 30064 22618 30076
rect 23768 30036 23796 30076
rect 20824 30008 23796 30036
rect 20717 29999 20775 30005
rect 23842 29996 23848 30048
rect 23900 30036 23906 30048
rect 24949 30039 25007 30045
rect 23900 30008 23945 30036
rect 23900 29996 23906 30008
rect 24949 30005 24961 30039
rect 24995 30036 25007 30039
rect 25130 30036 25136 30048
rect 24995 30008 25136 30036
rect 24995 30005 25007 30008
rect 24949 29999 25007 30005
rect 25130 29996 25136 30008
rect 25188 29996 25194 30048
rect 25700 30045 25728 30076
rect 26142 30064 26148 30076
rect 26200 30104 26206 30116
rect 28077 30107 28135 30113
rect 28077 30104 28089 30107
rect 26200 30076 28089 30104
rect 26200 30064 26206 30076
rect 28077 30073 28089 30076
rect 28123 30073 28135 30107
rect 28077 30067 28135 30073
rect 28626 30064 28632 30116
rect 28684 30104 28690 30116
rect 29932 30104 29960 30135
rect 30392 30113 30420 30144
rect 28684 30076 29960 30104
rect 30377 30107 30435 30113
rect 28684 30064 28690 30076
rect 30377 30073 30389 30107
rect 30423 30073 30435 30107
rect 30377 30067 30435 30073
rect 25685 30039 25743 30045
rect 25685 30005 25697 30039
rect 25731 30005 25743 30039
rect 25866 30036 25872 30048
rect 25827 30008 25872 30036
rect 25685 29999 25743 30005
rect 25866 29996 25872 30008
rect 25924 29996 25930 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 20901 29835 20959 29841
rect 20901 29801 20913 29835
rect 20947 29832 20959 29835
rect 21545 29835 21603 29841
rect 21545 29832 21557 29835
rect 20947 29804 21557 29832
rect 20947 29801 20959 29804
rect 20901 29795 20959 29801
rect 21545 29801 21557 29804
rect 21591 29801 21603 29835
rect 21910 29832 21916 29844
rect 21871 29804 21916 29832
rect 21545 29795 21603 29801
rect 21910 29792 21916 29804
rect 21968 29792 21974 29844
rect 25498 29832 25504 29844
rect 25459 29804 25504 29832
rect 25498 29792 25504 29804
rect 25556 29792 25562 29844
rect 26142 29832 26148 29844
rect 26103 29804 26148 29832
rect 26142 29792 26148 29804
rect 26200 29792 26206 29844
rect 27062 29832 27068 29844
rect 27023 29804 27068 29832
rect 27062 29792 27068 29804
rect 27120 29792 27126 29844
rect 27706 29832 27712 29844
rect 27667 29804 27712 29832
rect 27706 29792 27712 29804
rect 27764 29792 27770 29844
rect 31110 29832 31116 29844
rect 31071 29804 31116 29832
rect 31110 29792 31116 29804
rect 31168 29792 31174 29844
rect 24210 29764 24216 29776
rect 21008 29736 24216 29764
rect 21008 29696 21036 29736
rect 24210 29724 24216 29736
rect 24268 29724 24274 29776
rect 24946 29724 24952 29776
rect 25004 29764 25010 29776
rect 26421 29767 26479 29773
rect 26421 29764 26433 29767
rect 25004 29736 26433 29764
rect 25004 29724 25010 29736
rect 26421 29733 26433 29736
rect 26467 29733 26479 29767
rect 26421 29727 26479 29733
rect 18156 29668 21036 29696
rect 27632 29668 30880 29696
rect 13814 29588 13820 29640
rect 13872 29628 13878 29640
rect 14185 29631 14243 29637
rect 14185 29628 14197 29631
rect 13872 29600 14197 29628
rect 13872 29588 13878 29600
rect 14185 29597 14197 29600
rect 14231 29628 14243 29631
rect 14829 29631 14887 29637
rect 14829 29628 14841 29631
rect 14231 29600 14841 29628
rect 14231 29597 14243 29600
rect 14185 29591 14243 29597
rect 14829 29597 14841 29600
rect 14875 29597 14887 29631
rect 17310 29628 17316 29640
rect 17271 29600 17316 29628
rect 14829 29591 14887 29597
rect 17310 29588 17316 29600
rect 17368 29588 17374 29640
rect 17586 29628 17592 29640
rect 17547 29600 17592 29628
rect 17586 29588 17592 29600
rect 17644 29588 17650 29640
rect 17497 29563 17555 29569
rect 17497 29529 17509 29563
rect 17543 29560 17555 29563
rect 18156 29560 18184 29668
rect 18230 29588 18236 29640
rect 18288 29628 18294 29640
rect 20254 29628 20260 29640
rect 18288 29600 20260 29628
rect 18288 29588 18294 29600
rect 20254 29588 20260 29600
rect 20312 29588 20318 29640
rect 20438 29588 20444 29640
rect 20496 29628 20502 29640
rect 20533 29631 20591 29637
rect 20533 29628 20545 29631
rect 20496 29600 20545 29628
rect 20496 29588 20502 29600
rect 20533 29597 20545 29600
rect 20579 29597 20591 29631
rect 20533 29591 20591 29597
rect 20714 29588 20720 29640
rect 20772 29628 20778 29640
rect 20809 29631 20867 29637
rect 20809 29628 20821 29631
rect 20772 29600 20821 29628
rect 20772 29588 20778 29600
rect 20809 29597 20821 29600
rect 20855 29597 20867 29631
rect 20809 29591 20867 29597
rect 21729 29631 21787 29637
rect 21729 29597 21741 29631
rect 21775 29597 21787 29631
rect 22002 29628 22008 29640
rect 21963 29600 22008 29628
rect 21729 29591 21787 29597
rect 21174 29560 21180 29572
rect 17543 29532 18184 29560
rect 19904 29532 21180 29560
rect 17543 29529 17555 29532
rect 17497 29523 17555 29529
rect 14274 29492 14280 29504
rect 14235 29464 14280 29492
rect 14274 29452 14280 29464
rect 14332 29452 14338 29504
rect 14918 29492 14924 29504
rect 14879 29464 14924 29492
rect 14918 29452 14924 29464
rect 14976 29452 14982 29504
rect 16666 29452 16672 29504
rect 16724 29492 16730 29504
rect 17129 29495 17187 29501
rect 17129 29492 17141 29495
rect 16724 29464 17141 29492
rect 16724 29452 16730 29464
rect 17129 29461 17141 29464
rect 17175 29461 17187 29495
rect 17129 29455 17187 29461
rect 18598 29452 18604 29504
rect 18656 29492 18662 29504
rect 18874 29492 18880 29504
rect 18656 29464 18880 29492
rect 18656 29452 18662 29464
rect 18874 29452 18880 29464
rect 18932 29492 18938 29504
rect 19904 29492 19932 29532
rect 21174 29520 21180 29532
rect 21232 29520 21238 29572
rect 21744 29560 21772 29591
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 22370 29588 22376 29640
rect 22428 29628 22434 29640
rect 22465 29631 22523 29637
rect 22465 29628 22477 29631
rect 22428 29600 22477 29628
rect 22428 29588 22434 29600
rect 22465 29597 22477 29600
rect 22511 29597 22523 29631
rect 22465 29591 22523 29597
rect 23658 29588 23664 29640
rect 23716 29628 23722 29640
rect 24397 29631 24455 29637
rect 24397 29628 24409 29631
rect 23716 29600 24409 29628
rect 23716 29588 23722 29600
rect 24397 29597 24409 29600
rect 24443 29597 24455 29631
rect 25866 29628 25872 29640
rect 24397 29591 24455 29597
rect 24504 29600 25872 29628
rect 22094 29560 22100 29572
rect 21744 29532 22100 29560
rect 22094 29520 22100 29532
rect 22152 29520 22158 29572
rect 24504 29560 24532 29600
rect 25866 29588 25872 29600
rect 25924 29588 25930 29640
rect 26050 29628 26056 29640
rect 26011 29600 26056 29628
rect 26050 29588 26056 29600
rect 26108 29588 26114 29640
rect 26142 29588 26148 29640
rect 26200 29628 26206 29640
rect 26973 29631 27031 29637
rect 26200 29600 26245 29628
rect 26200 29588 26206 29600
rect 26973 29597 26985 29631
rect 27019 29628 27031 29631
rect 27338 29628 27344 29640
rect 27019 29600 27344 29628
rect 27019 29597 27031 29600
rect 26973 29591 27031 29597
rect 27338 29588 27344 29600
rect 27396 29588 27402 29640
rect 27632 29637 27660 29668
rect 30852 29640 30880 29668
rect 27617 29631 27675 29637
rect 27617 29597 27629 29631
rect 27663 29597 27675 29631
rect 27617 29591 27675 29597
rect 28350 29588 28356 29640
rect 28408 29628 28414 29640
rect 28445 29631 28503 29637
rect 28445 29628 28457 29631
rect 28408 29600 28457 29628
rect 28408 29588 28414 29600
rect 28445 29597 28457 29600
rect 28491 29597 28503 29631
rect 28626 29628 28632 29640
rect 28587 29600 28632 29628
rect 28445 29591 28503 29597
rect 28626 29588 28632 29600
rect 28684 29588 28690 29640
rect 28994 29588 29000 29640
rect 29052 29628 29058 29640
rect 30282 29628 30288 29640
rect 29052 29600 30288 29628
rect 29052 29588 29058 29600
rect 30282 29588 30288 29600
rect 30340 29588 30346 29640
rect 30834 29588 30840 29640
rect 30892 29628 30898 29640
rect 31021 29631 31079 29637
rect 31021 29628 31033 29631
rect 30892 29600 31033 29628
rect 30892 29588 30898 29600
rect 31021 29597 31033 29600
rect 31067 29597 31079 29631
rect 47302 29628 47308 29640
rect 47263 29600 47308 29628
rect 31021 29591 31079 29597
rect 47302 29588 47308 29600
rect 47360 29588 47366 29640
rect 47394 29588 47400 29640
rect 47452 29628 47458 29640
rect 47581 29631 47639 29637
rect 47581 29628 47593 29631
rect 47452 29600 47593 29628
rect 47452 29588 47458 29600
rect 47581 29597 47593 29600
rect 47627 29597 47639 29631
rect 47581 29591 47639 29597
rect 22388 29532 24532 29560
rect 25409 29563 25467 29569
rect 18932 29464 19932 29492
rect 18932 29452 18938 29464
rect 20530 29452 20536 29504
rect 20588 29492 20594 29504
rect 21085 29495 21143 29501
rect 21085 29492 21097 29495
rect 20588 29464 21097 29492
rect 20588 29452 20594 29464
rect 21085 29461 21097 29464
rect 21131 29461 21143 29495
rect 21085 29455 21143 29461
rect 21266 29452 21272 29504
rect 21324 29492 21330 29504
rect 22388 29492 22416 29532
rect 25409 29529 25421 29563
rect 25455 29560 25467 29563
rect 26160 29560 26188 29588
rect 29012 29560 29040 29588
rect 25455 29532 26188 29560
rect 26896 29532 29040 29560
rect 25455 29529 25467 29532
rect 25409 29523 25467 29529
rect 22554 29492 22560 29504
rect 21324 29464 22416 29492
rect 22515 29464 22560 29492
rect 21324 29452 21330 29464
rect 22554 29452 22560 29464
rect 22612 29452 22618 29504
rect 24210 29452 24216 29504
rect 24268 29492 24274 29504
rect 24581 29495 24639 29501
rect 24581 29492 24593 29495
rect 24268 29464 24593 29492
rect 24268 29452 24274 29464
rect 24581 29461 24593 29464
rect 24627 29492 24639 29495
rect 26896 29492 26924 29532
rect 24627 29464 26924 29492
rect 28537 29495 28595 29501
rect 24627 29461 24639 29464
rect 24581 29455 24639 29461
rect 28537 29461 28549 29495
rect 28583 29492 28595 29495
rect 28994 29492 29000 29504
rect 28583 29464 29000 29492
rect 28583 29461 28595 29464
rect 28537 29455 28595 29461
rect 28994 29452 29000 29464
rect 29052 29452 29058 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 13446 29288 13452 29300
rect 13407 29260 13452 29288
rect 13446 29248 13452 29260
rect 13504 29248 13510 29300
rect 17586 29288 17592 29300
rect 17547 29260 17592 29288
rect 17586 29248 17592 29260
rect 17644 29248 17650 29300
rect 20438 29288 20444 29300
rect 17972 29260 20444 29288
rect 14274 29220 14280 29232
rect 14235 29192 14280 29220
rect 14274 29180 14280 29192
rect 14332 29180 14338 29232
rect 15930 29220 15936 29232
rect 15891 29192 15936 29220
rect 15930 29180 15936 29192
rect 15988 29180 15994 29232
rect 17972 29220 18000 29260
rect 19794 29220 19800 29232
rect 16776 29192 18000 29220
rect 18064 29192 19800 29220
rect 13357 29155 13415 29161
rect 13357 29121 13369 29155
rect 13403 29152 13415 29155
rect 13814 29152 13820 29164
rect 13403 29124 13820 29152
rect 13403 29121 13415 29124
rect 13357 29115 13415 29121
rect 13814 29112 13820 29124
rect 13872 29112 13878 29164
rect 11698 29044 11704 29096
rect 11756 29084 11762 29096
rect 14093 29087 14151 29093
rect 14093 29084 14105 29087
rect 11756 29056 14105 29084
rect 11756 29044 11762 29056
rect 14093 29053 14105 29056
rect 14139 29053 14151 29087
rect 16776 29084 16804 29192
rect 16850 29112 16856 29164
rect 16908 29152 16914 29164
rect 17221 29155 17279 29161
rect 17221 29152 17233 29155
rect 16908 29124 17233 29152
rect 16908 29112 16914 29124
rect 17221 29121 17233 29124
rect 17267 29152 17279 29155
rect 17954 29152 17960 29164
rect 17267 29124 17960 29152
rect 17267 29121 17279 29124
rect 17221 29115 17279 29121
rect 17954 29112 17960 29124
rect 18012 29112 18018 29164
rect 18064 29161 18092 29192
rect 19794 29180 19800 29192
rect 19852 29180 19858 29232
rect 18049 29155 18107 29161
rect 18049 29121 18061 29155
rect 18095 29121 18107 29155
rect 18230 29152 18236 29164
rect 18191 29124 18236 29152
rect 18049 29115 18107 29121
rect 18230 29112 18236 29124
rect 18288 29112 18294 29164
rect 18325 29155 18383 29161
rect 18325 29121 18337 29155
rect 18371 29152 18383 29155
rect 18371 29124 18552 29152
rect 18371 29121 18383 29124
rect 18325 29115 18383 29121
rect 17129 29087 17187 29093
rect 17129 29084 17141 29087
rect 16776 29056 17141 29084
rect 14093 29047 14151 29053
rect 17129 29053 17141 29056
rect 17175 29053 17187 29087
rect 17129 29047 17187 29053
rect 18417 29087 18475 29093
rect 18417 29053 18429 29087
rect 18463 29053 18475 29087
rect 18524 29084 18552 29124
rect 18598 29112 18604 29164
rect 18656 29152 18662 29164
rect 19429 29155 19487 29161
rect 18656 29124 18701 29152
rect 18656 29112 18662 29124
rect 19429 29121 19441 29155
rect 19475 29121 19487 29155
rect 19429 29115 19487 29121
rect 19613 29155 19671 29161
rect 19613 29121 19625 29155
rect 19659 29152 19671 29155
rect 19904 29152 19932 29260
rect 20438 29248 20444 29260
rect 20496 29248 20502 29300
rect 30377 29291 30435 29297
rect 30377 29288 30389 29291
rect 28092 29260 30389 29288
rect 20254 29180 20260 29232
rect 20312 29220 20318 29232
rect 20312 29192 20760 29220
rect 20312 29180 20318 29192
rect 20530 29152 20536 29164
rect 19659 29124 19932 29152
rect 20491 29124 20536 29152
rect 19659 29121 19671 29124
rect 19613 29115 19671 29121
rect 19150 29084 19156 29096
rect 18524 29056 19156 29084
rect 18417 29047 18475 29053
rect 7834 28976 7840 29028
rect 7892 29016 7898 29028
rect 18432 29016 18460 29047
rect 19150 29044 19156 29056
rect 19208 29084 19214 29096
rect 19444 29084 19472 29115
rect 20530 29112 20536 29124
rect 20588 29112 20594 29164
rect 20732 29161 20760 29192
rect 20824 29192 22048 29220
rect 20824 29161 20852 29192
rect 20717 29155 20775 29161
rect 20717 29121 20729 29155
rect 20763 29121 20775 29155
rect 20717 29115 20775 29121
rect 20809 29155 20867 29161
rect 20809 29121 20821 29155
rect 20855 29121 20867 29155
rect 20809 29115 20867 29121
rect 21085 29155 21143 29161
rect 21085 29121 21097 29155
rect 21131 29152 21143 29155
rect 21174 29152 21180 29164
rect 21131 29124 21180 29152
rect 21131 29121 21143 29124
rect 21085 29115 21143 29121
rect 21174 29112 21180 29124
rect 21232 29112 21238 29164
rect 21358 29112 21364 29164
rect 21416 29152 21422 29164
rect 22020 29161 22048 29192
rect 21821 29155 21879 29161
rect 21821 29152 21833 29155
rect 21416 29124 21833 29152
rect 21416 29112 21422 29124
rect 21821 29121 21833 29124
rect 21867 29121 21879 29155
rect 21821 29115 21879 29121
rect 22005 29155 22063 29161
rect 22005 29121 22017 29155
rect 22051 29152 22063 29155
rect 22094 29152 22100 29164
rect 22051 29124 22100 29152
rect 22051 29121 22063 29124
rect 22005 29115 22063 29121
rect 22094 29112 22100 29124
rect 22152 29152 22158 29164
rect 22646 29152 22652 29164
rect 22152 29124 22652 29152
rect 22152 29112 22158 29124
rect 22646 29112 22652 29124
rect 22704 29112 22710 29164
rect 25317 29155 25375 29161
rect 25317 29121 25329 29155
rect 25363 29152 25375 29155
rect 25498 29152 25504 29164
rect 25363 29124 25504 29152
rect 25363 29121 25375 29124
rect 25317 29115 25375 29121
rect 25498 29112 25504 29124
rect 25556 29112 25562 29164
rect 28092 29152 28120 29260
rect 30377 29257 30389 29260
rect 30423 29257 30435 29291
rect 30377 29251 30435 29257
rect 28629 29223 28687 29229
rect 28629 29189 28641 29223
rect 28675 29189 28687 29223
rect 28629 29183 28687 29189
rect 29380 29192 30328 29220
rect 28169 29155 28227 29161
rect 28169 29152 28181 29155
rect 28092 29124 28181 29152
rect 28169 29121 28181 29124
rect 28215 29121 28227 29155
rect 28537 29155 28595 29161
rect 28537 29152 28549 29155
rect 28169 29115 28227 29121
rect 28276 29124 28549 29152
rect 19208 29056 19472 29084
rect 19705 29087 19763 29093
rect 19208 29044 19214 29056
rect 19705 29053 19717 29087
rect 19751 29053 19763 29087
rect 19705 29047 19763 29053
rect 20901 29087 20959 29093
rect 20901 29053 20913 29087
rect 20947 29053 20959 29087
rect 20901 29047 20959 29053
rect 7892 28988 18460 29016
rect 19245 29019 19303 29025
rect 7892 28976 7898 28988
rect 19245 28985 19257 29019
rect 19291 29016 19303 29019
rect 19334 29016 19340 29028
rect 19291 28988 19340 29016
rect 19291 28985 19303 28988
rect 19245 28979 19303 28985
rect 19334 28976 19340 28988
rect 19392 28976 19398 29028
rect 18046 28908 18052 28960
rect 18104 28948 18110 28960
rect 18785 28951 18843 28957
rect 18785 28948 18797 28951
rect 18104 28920 18797 28948
rect 18104 28908 18110 28920
rect 18785 28917 18797 28920
rect 18831 28917 18843 28951
rect 18785 28911 18843 28917
rect 19058 28908 19064 28960
rect 19116 28948 19122 28960
rect 19720 28948 19748 29047
rect 20916 29016 20944 29047
rect 23842 29044 23848 29096
rect 23900 29084 23906 29096
rect 25593 29087 25651 29093
rect 25593 29084 25605 29087
rect 23900 29056 25605 29084
rect 23900 29044 23906 29056
rect 25593 29053 25605 29056
rect 25639 29053 25651 29087
rect 25593 29047 25651 29053
rect 25682 29044 25688 29096
rect 25740 29084 25746 29096
rect 28276 29084 28304 29124
rect 28537 29121 28549 29124
rect 28583 29121 28595 29155
rect 28644 29152 28672 29183
rect 29089 29155 29147 29161
rect 29089 29152 29101 29155
rect 28644 29124 29101 29152
rect 28537 29115 28595 29121
rect 29089 29121 29101 29124
rect 29135 29121 29147 29155
rect 29089 29115 29147 29121
rect 29178 29112 29184 29164
rect 29236 29152 29242 29164
rect 29380 29161 29408 29192
rect 30300 29161 30328 29192
rect 29273 29155 29331 29161
rect 29273 29152 29285 29155
rect 29236 29124 29285 29152
rect 29236 29112 29242 29124
rect 29273 29121 29285 29124
rect 29319 29121 29331 29155
rect 29273 29115 29331 29121
rect 29365 29155 29423 29161
rect 29365 29121 29377 29155
rect 29411 29121 29423 29155
rect 29365 29115 29423 29121
rect 29641 29155 29699 29161
rect 29641 29121 29653 29155
rect 29687 29121 29699 29155
rect 29641 29115 29699 29121
rect 30285 29155 30343 29161
rect 30285 29121 30297 29155
rect 30331 29152 30343 29155
rect 30374 29152 30380 29164
rect 30331 29124 30380 29152
rect 30331 29121 30343 29124
rect 30285 29115 30343 29121
rect 25740 29056 28304 29084
rect 28445 29087 28503 29093
rect 25740 29044 25746 29056
rect 28445 29053 28457 29087
rect 28491 29084 28503 29087
rect 28902 29084 28908 29096
rect 28491 29056 28908 29084
rect 28491 29053 28503 29056
rect 28445 29047 28503 29053
rect 28902 29044 28908 29056
rect 28960 29044 28966 29096
rect 29454 29044 29460 29096
rect 29512 29084 29518 29096
rect 29512 29056 29557 29084
rect 29512 29044 29518 29056
rect 21726 29016 21732 29028
rect 20916 28988 21732 29016
rect 21726 28976 21732 28988
rect 21784 28976 21790 29028
rect 21818 28976 21824 29028
rect 21876 29016 21882 29028
rect 22189 29019 22247 29025
rect 22189 29016 22201 29019
rect 21876 28988 22201 29016
rect 21876 28976 21882 28988
rect 22189 28985 22201 28988
rect 22235 28985 22247 29019
rect 22189 28979 22247 28985
rect 25869 29019 25927 29025
rect 25869 28985 25881 29019
rect 25915 29016 25927 29019
rect 26418 29016 26424 29028
rect 25915 28988 26424 29016
rect 25915 28985 25927 28988
rect 25869 28979 25927 28985
rect 26418 28976 26424 28988
rect 26476 28976 26482 29028
rect 27246 28976 27252 29028
rect 27304 29016 27310 29028
rect 28261 29019 28319 29025
rect 27304 28988 28212 29016
rect 27304 28976 27310 28988
rect 19116 28920 19748 28948
rect 19116 28908 19122 28920
rect 21174 28908 21180 28960
rect 21232 28948 21238 28960
rect 21269 28951 21327 28957
rect 21269 28948 21281 28951
rect 21232 28920 21281 28948
rect 21232 28908 21238 28920
rect 21269 28917 21281 28920
rect 21315 28917 21327 28951
rect 22002 28948 22008 28960
rect 21963 28920 22008 28948
rect 21269 28911 21327 28917
rect 22002 28908 22008 28920
rect 22060 28908 22066 28960
rect 25406 28948 25412 28960
rect 25367 28920 25412 28948
rect 25406 28908 25412 28920
rect 25464 28908 25470 28960
rect 28184 28948 28212 28988
rect 28261 28985 28273 29019
rect 28307 29016 28319 29019
rect 28994 29016 29000 29028
rect 28307 28988 29000 29016
rect 28307 28985 28319 28988
rect 28261 28979 28319 28985
rect 28994 28976 29000 28988
rect 29052 28976 29058 29028
rect 29656 29016 29684 29115
rect 30374 29112 30380 29124
rect 30432 29152 30438 29164
rect 31662 29152 31668 29164
rect 30432 29124 31668 29152
rect 30432 29112 30438 29124
rect 31662 29112 31668 29124
rect 31720 29112 31726 29164
rect 29104 28988 29684 29016
rect 29104 28948 29132 28988
rect 28184 28920 29132 28948
rect 29825 28951 29883 28957
rect 29825 28917 29837 28951
rect 29871 28948 29883 28951
rect 30190 28948 30196 28960
rect 29871 28920 30196 28948
rect 29871 28917 29883 28920
rect 29825 28911 29883 28917
rect 30190 28908 30196 28920
rect 30248 28908 30254 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 11974 28744 11980 28756
rect 10428 28716 11980 28744
rect 10428 28549 10456 28716
rect 11974 28704 11980 28716
rect 12032 28744 12038 28756
rect 12989 28747 13047 28753
rect 12989 28744 13001 28747
rect 12032 28716 13001 28744
rect 12032 28704 12038 28716
rect 12989 28713 13001 28716
rect 13035 28713 13047 28747
rect 12989 28707 13047 28713
rect 10505 28611 10563 28617
rect 10505 28577 10517 28611
rect 10551 28608 10563 28611
rect 11606 28608 11612 28620
rect 10551 28580 11612 28608
rect 10551 28577 10563 28580
rect 10505 28571 10563 28577
rect 11606 28568 11612 28580
rect 11664 28568 11670 28620
rect 13004 28608 13032 28707
rect 17954 28704 17960 28756
rect 18012 28744 18018 28756
rect 18141 28747 18199 28753
rect 18141 28744 18153 28747
rect 18012 28716 18153 28744
rect 18012 28704 18018 28716
rect 18141 28713 18153 28716
rect 18187 28744 18199 28747
rect 19058 28744 19064 28756
rect 18187 28716 19064 28744
rect 18187 28713 18199 28716
rect 18141 28707 18199 28713
rect 19058 28704 19064 28716
rect 19116 28704 19122 28756
rect 19334 28744 19340 28756
rect 19295 28716 19340 28744
rect 19334 28704 19340 28716
rect 19392 28704 19398 28756
rect 19794 28744 19800 28756
rect 19755 28716 19800 28744
rect 19794 28704 19800 28716
rect 19852 28704 19858 28756
rect 20346 28704 20352 28756
rect 20404 28744 20410 28756
rect 21818 28744 21824 28756
rect 20404 28716 21824 28744
rect 20404 28704 20410 28716
rect 21818 28704 21824 28716
rect 21876 28704 21882 28756
rect 22646 28744 22652 28756
rect 22607 28716 22652 28744
rect 22646 28704 22652 28716
rect 22704 28704 22710 28756
rect 25406 28744 25412 28756
rect 25367 28716 25412 28744
rect 25406 28704 25412 28716
rect 25464 28704 25470 28756
rect 29288 28716 35894 28744
rect 23584 28648 24532 28676
rect 13262 28608 13268 28620
rect 13004 28580 13268 28608
rect 13262 28568 13268 28580
rect 13320 28608 13326 28620
rect 14093 28611 14151 28617
rect 14093 28608 14105 28611
rect 13320 28580 14105 28608
rect 13320 28568 13326 28580
rect 14093 28577 14105 28580
rect 14139 28577 14151 28611
rect 14093 28571 14151 28577
rect 14277 28611 14335 28617
rect 14277 28577 14289 28611
rect 14323 28608 14335 28611
rect 14918 28608 14924 28620
rect 14323 28580 14924 28608
rect 14323 28577 14335 28580
rect 14277 28571 14335 28577
rect 14918 28568 14924 28580
rect 14976 28568 14982 28620
rect 16022 28568 16028 28620
rect 16080 28608 16086 28620
rect 16393 28611 16451 28617
rect 16393 28608 16405 28611
rect 16080 28580 16405 28608
rect 16080 28568 16086 28580
rect 16393 28577 16405 28580
rect 16439 28577 16451 28611
rect 16666 28608 16672 28620
rect 16627 28580 16672 28608
rect 16393 28571 16451 28577
rect 16666 28568 16672 28580
rect 16724 28568 16730 28620
rect 19426 28568 19432 28620
rect 19484 28608 19490 28620
rect 20898 28608 20904 28620
rect 19484 28580 20904 28608
rect 19484 28568 19490 28580
rect 20898 28568 20904 28580
rect 20956 28568 20962 28620
rect 21174 28608 21180 28620
rect 21135 28580 21180 28608
rect 21174 28568 21180 28580
rect 21232 28568 21238 28620
rect 23474 28568 23480 28620
rect 23532 28608 23538 28620
rect 23584 28617 23612 28648
rect 23569 28611 23627 28617
rect 23569 28608 23581 28611
rect 23532 28580 23581 28608
rect 23532 28568 23538 28580
rect 23569 28577 23581 28580
rect 23615 28577 23627 28611
rect 23750 28608 23756 28620
rect 23711 28580 23756 28608
rect 23569 28571 23627 28577
rect 23750 28568 23756 28580
rect 23808 28568 23814 28620
rect 10413 28543 10471 28549
rect 10413 28509 10425 28543
rect 10459 28509 10471 28543
rect 10413 28503 10471 28509
rect 10870 28500 10876 28552
rect 10928 28540 10934 28552
rect 11241 28543 11299 28549
rect 11241 28540 11253 28543
rect 10928 28512 11253 28540
rect 10928 28500 10934 28512
rect 11241 28509 11253 28512
rect 11287 28509 11299 28543
rect 11241 28503 11299 28509
rect 19245 28543 19303 28549
rect 19245 28509 19257 28543
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 19613 28543 19671 28549
rect 19613 28509 19625 28543
rect 19659 28540 19671 28543
rect 20714 28540 20720 28552
rect 19659 28512 20720 28540
rect 19659 28509 19671 28512
rect 19613 28503 19671 28509
rect 11517 28475 11575 28481
rect 11517 28441 11529 28475
rect 11563 28441 11575 28475
rect 11517 28435 11575 28441
rect 10781 28407 10839 28413
rect 10781 28373 10793 28407
rect 10827 28404 10839 28407
rect 11532 28404 11560 28435
rect 12526 28432 12532 28484
rect 12584 28432 12590 28484
rect 15933 28475 15991 28481
rect 15933 28441 15945 28475
rect 15979 28472 15991 28475
rect 16574 28472 16580 28484
rect 15979 28444 16580 28472
rect 15979 28441 15991 28444
rect 15933 28435 15991 28441
rect 16574 28432 16580 28444
rect 16632 28432 16638 28484
rect 17402 28432 17408 28484
rect 17460 28432 17466 28484
rect 10827 28376 11560 28404
rect 19260 28404 19288 28503
rect 20714 28500 20720 28512
rect 20772 28500 20778 28552
rect 24394 28540 24400 28552
rect 24355 28512 24400 28540
rect 24394 28500 24400 28512
rect 24452 28500 24458 28552
rect 24504 28540 24532 28648
rect 25869 28611 25927 28617
rect 25869 28608 25881 28611
rect 25240 28580 25881 28608
rect 24765 28543 24823 28549
rect 24765 28540 24777 28543
rect 24504 28512 24777 28540
rect 24765 28509 24777 28512
rect 24811 28509 24823 28543
rect 24765 28503 24823 28509
rect 25240 28484 25268 28580
rect 25869 28577 25881 28580
rect 25915 28577 25927 28611
rect 25869 28571 25927 28577
rect 26789 28611 26847 28617
rect 26789 28577 26801 28611
rect 26835 28608 26847 28611
rect 29288 28608 29316 28716
rect 31662 28676 31668 28688
rect 31623 28648 31668 28676
rect 31662 28636 31668 28648
rect 31720 28636 31726 28688
rect 30190 28608 30196 28620
rect 26835 28580 29316 28608
rect 30151 28580 30196 28608
rect 26835 28577 26847 28580
rect 26789 28571 26847 28577
rect 30190 28568 30196 28580
rect 30248 28568 30254 28620
rect 35866 28608 35894 28716
rect 40402 28608 40408 28620
rect 35866 28580 40408 28608
rect 40402 28568 40408 28580
rect 40460 28568 40466 28620
rect 46477 28611 46535 28617
rect 46477 28577 46489 28611
rect 46523 28608 46535 28611
rect 47394 28608 47400 28620
rect 46523 28580 47400 28608
rect 46523 28577 46535 28580
rect 46477 28571 46535 28577
rect 47394 28568 47400 28580
rect 47452 28568 47458 28620
rect 47854 28608 47860 28620
rect 47815 28580 47860 28608
rect 47854 28568 47860 28580
rect 47912 28568 47918 28620
rect 25593 28543 25651 28549
rect 25593 28509 25605 28543
rect 25639 28509 25651 28543
rect 25774 28540 25780 28552
rect 25735 28512 25780 28540
rect 25593 28503 25651 28509
rect 22554 28472 22560 28484
rect 22402 28444 22560 28472
rect 22554 28432 22560 28444
rect 22612 28432 22618 28484
rect 23477 28475 23535 28481
rect 23477 28441 23489 28475
rect 23523 28472 23535 28475
rect 23658 28472 23664 28484
rect 23523 28444 23664 28472
rect 23523 28441 23535 28444
rect 23477 28435 23535 28441
rect 23658 28432 23664 28444
rect 23716 28432 23722 28484
rect 24210 28432 24216 28484
rect 24268 28472 24274 28484
rect 24581 28475 24639 28481
rect 24581 28472 24593 28475
rect 24268 28444 24593 28472
rect 24268 28432 24274 28444
rect 24581 28441 24593 28444
rect 24627 28441 24639 28475
rect 24581 28435 24639 28441
rect 24673 28475 24731 28481
rect 24673 28441 24685 28475
rect 24719 28472 24731 28475
rect 25222 28472 25228 28484
rect 24719 28444 25228 28472
rect 24719 28441 24731 28444
rect 24673 28435 24731 28441
rect 25222 28432 25228 28444
rect 25280 28432 25286 28484
rect 25608 28472 25636 28503
rect 25774 28500 25780 28512
rect 25832 28500 25838 28552
rect 26418 28540 26424 28552
rect 26379 28512 26424 28540
rect 26418 28500 26424 28512
rect 26476 28500 26482 28552
rect 26602 28540 26608 28552
rect 26563 28512 26608 28540
rect 26602 28500 26608 28512
rect 26660 28500 26666 28552
rect 26694 28500 26700 28552
rect 26752 28540 26758 28552
rect 26973 28543 27031 28549
rect 26973 28540 26985 28543
rect 26752 28512 26797 28540
rect 26896 28512 26985 28540
rect 26752 28500 26758 28512
rect 26712 28472 26740 28500
rect 25608 28444 26740 28472
rect 20714 28404 20720 28416
rect 19260 28376 20720 28404
rect 10827 28373 10839 28376
rect 10781 28367 10839 28373
rect 20714 28364 20720 28376
rect 20772 28364 20778 28416
rect 22922 28364 22928 28416
rect 22980 28404 22986 28416
rect 23109 28407 23167 28413
rect 23109 28404 23121 28407
rect 22980 28376 23121 28404
rect 22980 28364 22986 28376
rect 23109 28373 23121 28376
rect 23155 28373 23167 28407
rect 23109 28367 23167 28373
rect 24486 28364 24492 28416
rect 24544 28404 24550 28416
rect 24949 28407 25007 28413
rect 24949 28404 24961 28407
rect 24544 28376 24961 28404
rect 24544 28364 24550 28376
rect 24949 28373 24961 28376
rect 24995 28373 25007 28407
rect 24949 28367 25007 28373
rect 26234 28364 26240 28416
rect 26292 28404 26298 28416
rect 26896 28404 26924 28512
rect 26973 28509 26985 28512
rect 27019 28540 27031 28543
rect 27246 28540 27252 28552
rect 27019 28512 27252 28540
rect 27019 28509 27031 28512
rect 26973 28503 27031 28509
rect 27246 28500 27252 28512
rect 27304 28500 27310 28552
rect 28169 28543 28227 28549
rect 28169 28509 28181 28543
rect 28215 28509 28227 28543
rect 28350 28540 28356 28552
rect 28311 28512 28356 28540
rect 28169 28503 28227 28509
rect 28184 28472 28212 28503
rect 28350 28500 28356 28512
rect 28408 28500 28414 28552
rect 29086 28500 29092 28552
rect 29144 28540 29150 28552
rect 29917 28543 29975 28549
rect 29917 28540 29929 28543
rect 29144 28512 29929 28540
rect 29144 28500 29150 28512
rect 29917 28509 29929 28512
rect 29963 28509 29975 28543
rect 46290 28540 46296 28552
rect 46251 28512 46296 28540
rect 29917 28503 29975 28509
rect 46290 28500 46296 28512
rect 46348 28500 46354 28552
rect 28626 28472 28632 28484
rect 28184 28444 28632 28472
rect 28626 28432 28632 28444
rect 28684 28432 28690 28484
rect 30926 28432 30932 28484
rect 30984 28432 30990 28484
rect 26292 28376 26924 28404
rect 27157 28407 27215 28413
rect 26292 28364 26298 28376
rect 27157 28373 27169 28407
rect 27203 28404 27215 28407
rect 27246 28404 27252 28416
rect 27203 28376 27252 28404
rect 27203 28373 27215 28376
rect 27157 28367 27215 28373
rect 27246 28364 27252 28376
rect 27304 28364 27310 28416
rect 28537 28407 28595 28413
rect 28537 28373 28549 28407
rect 28583 28404 28595 28407
rect 29178 28404 29184 28416
rect 28583 28376 29184 28404
rect 28583 28373 28595 28376
rect 28537 28367 28595 28373
rect 29178 28364 29184 28376
rect 29236 28364 29242 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 1670 28160 1676 28212
rect 1728 28200 1734 28212
rect 10870 28200 10876 28212
rect 1728 28172 6914 28200
rect 10831 28172 10876 28200
rect 1728 28160 1734 28172
rect 6886 28132 6914 28172
rect 10870 28160 10876 28172
rect 10928 28160 10934 28212
rect 11606 28200 11612 28212
rect 11567 28172 11612 28200
rect 11606 28160 11612 28172
rect 11664 28160 11670 28212
rect 12526 28200 12532 28212
rect 12487 28172 12532 28200
rect 12526 28160 12532 28172
rect 12584 28160 12590 28212
rect 19242 28200 19248 28212
rect 17512 28172 19248 28200
rect 6886 28104 15976 28132
rect 10502 28024 10508 28076
rect 10560 28064 10566 28076
rect 10781 28067 10839 28073
rect 10781 28064 10793 28067
rect 10560 28036 10793 28064
rect 10560 28024 10566 28036
rect 10781 28033 10793 28036
rect 10827 28033 10839 28067
rect 11514 28064 11520 28076
rect 11475 28036 11520 28064
rect 10781 28027 10839 28033
rect 11514 28024 11520 28036
rect 11572 28024 11578 28076
rect 11698 28064 11704 28076
rect 11659 28036 11704 28064
rect 11698 28024 11704 28036
rect 11756 28024 11762 28076
rect 12342 28024 12348 28076
rect 12400 28064 12406 28076
rect 12437 28067 12495 28073
rect 12437 28064 12449 28067
rect 12400 28036 12449 28064
rect 12400 28024 12406 28036
rect 12437 28033 12449 28036
rect 12483 28033 12495 28067
rect 12437 28027 12495 28033
rect 14090 27956 14096 28008
rect 14148 27996 14154 28008
rect 14277 27999 14335 28005
rect 14277 27996 14289 27999
rect 14148 27968 14289 27996
rect 14148 27956 14154 27968
rect 14277 27965 14289 27968
rect 14323 27965 14335 27999
rect 14458 27996 14464 28008
rect 14419 27968 14464 27996
rect 14277 27959 14335 27965
rect 14458 27956 14464 27968
rect 14516 27956 14522 28008
rect 14737 27999 14795 28005
rect 14737 27965 14749 27999
rect 14783 27965 14795 27999
rect 15948 27996 15976 28104
rect 16022 28024 16028 28076
rect 16080 28064 16086 28076
rect 17512 28073 17540 28172
rect 19242 28160 19248 28172
rect 19300 28200 19306 28212
rect 19426 28200 19432 28212
rect 19300 28172 19432 28200
rect 19300 28160 19306 28172
rect 19426 28160 19432 28172
rect 19484 28160 19490 28212
rect 20714 28160 20720 28212
rect 20772 28200 20778 28212
rect 20901 28203 20959 28209
rect 20901 28200 20913 28203
rect 20772 28172 20913 28200
rect 20772 28160 20778 28172
rect 20901 28169 20913 28172
rect 20947 28200 20959 28203
rect 21910 28200 21916 28212
rect 20947 28172 21916 28200
rect 20947 28169 20959 28172
rect 20901 28163 20959 28169
rect 21910 28160 21916 28172
rect 21968 28160 21974 28212
rect 22646 28160 22652 28212
rect 22704 28200 22710 28212
rect 23106 28200 23112 28212
rect 22704 28172 23112 28200
rect 22704 28160 22710 28172
rect 23106 28160 23112 28172
rect 23164 28160 23170 28212
rect 24394 28160 24400 28212
rect 24452 28200 24458 28212
rect 24857 28203 24915 28209
rect 24857 28200 24869 28203
rect 24452 28172 24869 28200
rect 24452 28160 24458 28172
rect 24857 28169 24869 28172
rect 24903 28169 24915 28203
rect 24857 28163 24915 28169
rect 25869 28203 25927 28209
rect 25869 28169 25881 28203
rect 25915 28200 25927 28203
rect 26142 28200 26148 28212
rect 25915 28172 26148 28200
rect 25915 28169 25927 28172
rect 25869 28163 25927 28169
rect 26142 28160 26148 28172
rect 26200 28160 26206 28212
rect 26694 28160 26700 28212
rect 26752 28200 26758 28212
rect 28721 28203 28779 28209
rect 28721 28200 28733 28203
rect 26752 28172 28733 28200
rect 26752 28160 26758 28172
rect 28721 28169 28733 28172
rect 28767 28169 28779 28203
rect 30926 28200 30932 28212
rect 30887 28172 30932 28200
rect 28721 28163 28779 28169
rect 30926 28160 30932 28172
rect 30984 28160 30990 28212
rect 47854 28200 47860 28212
rect 35866 28172 47860 28200
rect 17773 28135 17831 28141
rect 17773 28101 17785 28135
rect 17819 28132 17831 28135
rect 18046 28132 18052 28144
rect 17819 28104 18052 28132
rect 17819 28101 17831 28104
rect 17773 28095 17831 28101
rect 18046 28092 18052 28104
rect 18104 28092 18110 28144
rect 18506 28092 18512 28144
rect 18564 28092 18570 28144
rect 19058 28092 19064 28144
rect 19116 28132 19122 28144
rect 19705 28135 19763 28141
rect 19705 28132 19717 28135
rect 19116 28104 19717 28132
rect 19116 28092 19122 28104
rect 19705 28101 19717 28104
rect 19751 28101 19763 28135
rect 19705 28095 19763 28101
rect 17497 28067 17555 28073
rect 17497 28064 17509 28067
rect 16080 28036 17509 28064
rect 16080 28024 16086 28036
rect 17497 28033 17509 28036
rect 17543 28033 17555 28067
rect 17497 28027 17555 28033
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28033 19947 28067
rect 19889 28027 19947 28033
rect 20073 28067 20131 28073
rect 20073 28033 20085 28067
rect 20119 28064 20131 28067
rect 20530 28064 20536 28076
rect 20119 28036 20536 28064
rect 20119 28033 20131 28036
rect 20073 28027 20131 28033
rect 15948 27968 18828 27996
rect 14737 27959 14795 27965
rect 3326 27888 3332 27940
rect 3384 27928 3390 27940
rect 14182 27928 14188 27940
rect 3384 27900 14188 27928
rect 3384 27888 3390 27900
rect 14182 27888 14188 27900
rect 14240 27888 14246 27940
rect 14366 27888 14372 27940
rect 14424 27928 14430 27940
rect 14752 27928 14780 27959
rect 14424 27900 14780 27928
rect 18800 27928 18828 27968
rect 19150 27956 19156 28008
rect 19208 27996 19214 28008
rect 19245 27999 19303 28005
rect 19245 27996 19257 27999
rect 19208 27968 19257 27996
rect 19208 27956 19214 27968
rect 19245 27965 19257 27968
rect 19291 27996 19303 27999
rect 19904 27996 19932 28027
rect 20530 28024 20536 28036
rect 20588 28024 20594 28076
rect 20622 28024 20628 28076
rect 20680 28064 20686 28076
rect 21818 28064 21824 28076
rect 20680 28036 20725 28064
rect 21779 28036 21824 28064
rect 20680 28024 20686 28036
rect 21818 28024 21824 28036
rect 21876 28024 21882 28076
rect 22922 28064 22928 28076
rect 22883 28036 22928 28064
rect 22922 28024 22928 28036
rect 22980 28024 22986 28076
rect 23201 28067 23259 28073
rect 23201 28033 23213 28067
rect 23247 28033 23259 28067
rect 23201 28027 23259 28033
rect 24489 28067 24547 28073
rect 24489 28033 24501 28067
rect 24535 28064 24547 28067
rect 25222 28064 25228 28076
rect 24535 28036 25228 28064
rect 24535 28033 24547 28036
rect 24489 28027 24547 28033
rect 19291 27968 19932 27996
rect 19291 27965 19303 27968
rect 19245 27959 19303 27965
rect 23216 27928 23244 28027
rect 25222 28024 25228 28036
rect 25280 28024 25286 28076
rect 25406 28064 25412 28076
rect 25367 28036 25412 28064
rect 25406 28024 25412 28036
rect 25464 28024 25470 28076
rect 25685 28067 25743 28073
rect 25685 28033 25697 28067
rect 25731 28064 25743 28067
rect 26712 28064 26740 28160
rect 27246 28132 27252 28144
rect 27207 28104 27252 28132
rect 27246 28092 27252 28104
rect 27304 28092 27310 28144
rect 27982 28092 27988 28144
rect 28040 28092 28046 28144
rect 26970 28064 26976 28076
rect 25731 28036 26740 28064
rect 26931 28036 26976 28064
rect 25731 28033 25743 28036
rect 25685 28027 25743 28033
rect 26970 28024 26976 28036
rect 27028 28024 27034 28076
rect 29178 28064 29184 28076
rect 29139 28036 29184 28064
rect 29178 28024 29184 28036
rect 29236 28024 29242 28076
rect 30834 28064 30840 28076
rect 30795 28036 30840 28064
rect 30834 28024 30840 28036
rect 30892 28024 30898 28076
rect 24581 27999 24639 28005
rect 24581 27965 24593 27999
rect 24627 27965 24639 27999
rect 25590 27996 25596 28008
rect 25551 27968 25596 27996
rect 24581 27959 24639 27965
rect 18800 27900 23244 27928
rect 24596 27928 24624 27959
rect 25590 27956 25596 27968
rect 25648 27956 25654 28008
rect 25866 27956 25872 28008
rect 25924 27996 25930 28008
rect 29273 27999 29331 28005
rect 29273 27996 29285 27999
rect 25924 27968 29285 27996
rect 25924 27956 25930 27968
rect 29273 27965 29285 27968
rect 29319 27965 29331 27999
rect 35866 27996 35894 28172
rect 47854 28160 47860 28172
rect 47912 28160 47918 28212
rect 47210 28024 47216 28076
rect 47268 28064 47274 28076
rect 47581 28067 47639 28073
rect 47581 28064 47593 28067
rect 47268 28036 47593 28064
rect 47268 28024 47274 28036
rect 47581 28033 47593 28036
rect 47627 28033 47639 28067
rect 47581 28027 47639 28033
rect 29273 27959 29331 27965
rect 31726 27968 35894 27996
rect 25774 27928 25780 27940
rect 24596 27900 25780 27928
rect 14424 27888 14430 27900
rect 25774 27888 25780 27900
rect 25832 27888 25838 27940
rect 28902 27888 28908 27940
rect 28960 27928 28966 27940
rect 31726 27928 31754 27968
rect 28960 27900 31754 27928
rect 28960 27888 28966 27900
rect 20346 27820 20352 27872
rect 20404 27860 20410 27872
rect 20533 27863 20591 27869
rect 20533 27860 20545 27863
rect 20404 27832 20545 27860
rect 20404 27820 20410 27832
rect 20533 27829 20545 27832
rect 20579 27829 20591 27863
rect 20533 27823 20591 27829
rect 21174 27820 21180 27872
rect 21232 27860 21238 27872
rect 21542 27860 21548 27872
rect 21232 27832 21548 27860
rect 21232 27820 21238 27832
rect 21542 27820 21548 27832
rect 21600 27860 21606 27872
rect 22005 27863 22063 27869
rect 22005 27860 22017 27863
rect 21600 27832 22017 27860
rect 21600 27820 21606 27832
rect 22005 27829 22017 27832
rect 22051 27829 22063 27863
rect 22738 27860 22744 27872
rect 22699 27832 22744 27860
rect 22005 27823 22063 27829
rect 22738 27820 22744 27832
rect 22796 27820 22802 27872
rect 25222 27820 25228 27872
rect 25280 27860 25286 27872
rect 25409 27863 25467 27869
rect 25409 27860 25421 27863
rect 25280 27832 25421 27860
rect 25280 27820 25286 27832
rect 25409 27829 25421 27832
rect 25455 27829 25467 27863
rect 25409 27823 25467 27829
rect 28994 27820 29000 27872
rect 29052 27860 29058 27872
rect 29181 27863 29239 27869
rect 29181 27860 29193 27863
rect 29052 27832 29193 27860
rect 29052 27820 29058 27832
rect 29181 27829 29193 27832
rect 29227 27829 29239 27863
rect 29546 27860 29552 27872
rect 29507 27832 29552 27860
rect 29181 27823 29239 27829
rect 29546 27820 29552 27832
rect 29604 27820 29610 27872
rect 47026 27860 47032 27872
rect 46987 27832 47032 27860
rect 47026 27820 47032 27832
rect 47084 27820 47090 27872
rect 47670 27860 47676 27872
rect 47631 27832 47676 27860
rect 47670 27820 47676 27832
rect 47728 27820 47734 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 14458 27616 14464 27668
rect 14516 27656 14522 27668
rect 14829 27659 14887 27665
rect 14829 27656 14841 27659
rect 14516 27628 14841 27656
rect 14516 27616 14522 27628
rect 14829 27625 14841 27628
rect 14875 27625 14887 27659
rect 14829 27619 14887 27625
rect 20346 27616 20352 27668
rect 20404 27656 20410 27668
rect 20533 27659 20591 27665
rect 20533 27656 20545 27659
rect 20404 27628 20545 27656
rect 20404 27616 20410 27628
rect 20533 27625 20545 27628
rect 20579 27625 20591 27659
rect 20533 27619 20591 27625
rect 22360 27659 22418 27665
rect 22360 27625 22372 27659
rect 22406 27656 22418 27659
rect 22738 27656 22744 27668
rect 22406 27628 22744 27656
rect 22406 27625 22418 27628
rect 22360 27619 22418 27625
rect 22738 27616 22744 27628
rect 22796 27616 22802 27668
rect 25961 27659 26019 27665
rect 25961 27625 25973 27659
rect 26007 27656 26019 27659
rect 26510 27656 26516 27668
rect 26007 27628 26516 27656
rect 26007 27625 26019 27628
rect 25961 27619 26019 27625
rect 26510 27616 26516 27628
rect 26568 27616 26574 27668
rect 26970 27616 26976 27668
rect 27028 27656 27034 27668
rect 29086 27656 29092 27668
rect 27028 27628 29092 27656
rect 27028 27616 27034 27628
rect 29086 27616 29092 27628
rect 29144 27616 29150 27668
rect 32214 27616 32220 27668
rect 32272 27656 32278 27668
rect 45554 27656 45560 27668
rect 32272 27628 45560 27656
rect 32272 27616 32278 27628
rect 45554 27616 45560 27628
rect 45612 27616 45618 27668
rect 17402 27548 17408 27600
rect 17460 27588 17466 27600
rect 17497 27591 17555 27597
rect 17497 27588 17509 27591
rect 17460 27560 17509 27588
rect 17460 27548 17466 27560
rect 17497 27557 17509 27560
rect 17543 27557 17555 27591
rect 18506 27588 18512 27600
rect 18467 27560 18512 27588
rect 17497 27551 17555 27557
rect 18506 27548 18512 27560
rect 18564 27548 18570 27600
rect 20993 27591 21051 27597
rect 20993 27557 21005 27591
rect 21039 27588 21051 27591
rect 21818 27588 21824 27600
rect 21039 27560 21824 27588
rect 21039 27557 21051 27560
rect 20993 27551 21051 27557
rect 21818 27548 21824 27560
rect 21876 27548 21882 27600
rect 23382 27548 23388 27600
rect 23440 27588 23446 27600
rect 23440 27560 27476 27588
rect 23440 27548 23446 27560
rect 13814 27480 13820 27532
rect 13872 27520 13878 27532
rect 13872 27492 14780 27520
rect 13872 27480 13878 27492
rect 14752 27464 14780 27492
rect 20530 27480 20536 27532
rect 20588 27520 20594 27532
rect 20625 27523 20683 27529
rect 20625 27520 20637 27523
rect 20588 27492 20637 27520
rect 20588 27480 20594 27492
rect 20625 27489 20637 27492
rect 20671 27489 20683 27523
rect 20625 27483 20683 27489
rect 20898 27480 20904 27532
rect 20956 27520 20962 27532
rect 22097 27523 22155 27529
rect 22097 27520 22109 27523
rect 20956 27492 22109 27520
rect 20956 27480 20962 27492
rect 22097 27489 22109 27492
rect 22143 27489 22155 27523
rect 22097 27483 22155 27489
rect 23750 27480 23756 27532
rect 23808 27520 23814 27532
rect 23845 27523 23903 27529
rect 23845 27520 23857 27523
rect 23808 27492 23857 27520
rect 23808 27480 23814 27492
rect 23845 27489 23857 27492
rect 23891 27520 23903 27523
rect 25406 27520 25412 27532
rect 23891 27492 25412 27520
rect 23891 27489 23903 27492
rect 23845 27483 23903 27489
rect 11146 27452 11152 27464
rect 11107 27424 11152 27452
rect 11146 27412 11152 27424
rect 11204 27412 11210 27464
rect 11333 27455 11391 27461
rect 11333 27421 11345 27455
rect 11379 27421 11391 27455
rect 11333 27415 11391 27421
rect 11977 27455 12035 27461
rect 11977 27421 11989 27455
rect 12023 27452 12035 27455
rect 12342 27452 12348 27464
rect 12023 27424 12348 27452
rect 12023 27421 12035 27424
rect 11977 27415 12035 27421
rect 11348 27384 11376 27415
rect 12342 27412 12348 27424
rect 12400 27452 12406 27464
rect 13906 27452 13912 27464
rect 12400 27424 13912 27452
rect 12400 27412 12406 27424
rect 13906 27412 13912 27424
rect 13964 27452 13970 27464
rect 14093 27455 14151 27461
rect 14093 27452 14105 27455
rect 13964 27424 14105 27452
rect 13964 27412 13970 27424
rect 14093 27421 14105 27424
rect 14139 27421 14151 27455
rect 14734 27452 14740 27464
rect 14695 27424 14740 27452
rect 14093 27415 14151 27421
rect 14734 27412 14740 27424
rect 14792 27412 14798 27464
rect 17405 27455 17463 27461
rect 17405 27421 17417 27455
rect 17451 27452 17463 27455
rect 18417 27455 18475 27461
rect 18417 27452 18429 27455
rect 17451 27424 18429 27452
rect 17451 27421 17463 27424
rect 17405 27415 17463 27421
rect 18417 27421 18429 27424
rect 18463 27452 18475 27455
rect 19058 27452 19064 27464
rect 18463 27424 19064 27452
rect 18463 27421 18475 27424
rect 18417 27415 18475 27421
rect 19058 27412 19064 27424
rect 19116 27412 19122 27464
rect 20809 27455 20867 27461
rect 20809 27421 20821 27455
rect 20855 27452 20867 27455
rect 21082 27452 21088 27464
rect 20855 27424 21088 27452
rect 20855 27421 20867 27424
rect 20809 27415 20867 27421
rect 21082 27412 21088 27424
rect 21140 27412 21146 27464
rect 24780 27461 24808 27492
rect 25406 27480 25412 27492
rect 25464 27520 25470 27532
rect 25464 27492 26096 27520
rect 25464 27480 25470 27492
rect 24765 27455 24823 27461
rect 24765 27421 24777 27455
rect 24811 27421 24823 27455
rect 24765 27415 24823 27421
rect 25133 27455 25191 27461
rect 25133 27421 25145 27455
rect 25179 27452 25191 27455
rect 25593 27455 25651 27461
rect 25593 27452 25605 27455
rect 25179 27424 25605 27452
rect 25179 27421 25191 27424
rect 25133 27415 25191 27421
rect 25593 27421 25605 27424
rect 25639 27452 25651 27455
rect 25774 27452 25780 27464
rect 25639 27424 25780 27452
rect 25639 27421 25651 27424
rect 25593 27415 25651 27421
rect 25774 27412 25780 27424
rect 25832 27412 25838 27464
rect 25866 27412 25872 27464
rect 25924 27452 25930 27464
rect 25924 27424 25969 27452
rect 25924 27412 25930 27424
rect 12434 27384 12440 27396
rect 11348 27356 12440 27384
rect 12434 27344 12440 27356
rect 12492 27344 12498 27396
rect 20533 27387 20591 27393
rect 20533 27353 20545 27387
rect 20579 27384 20591 27387
rect 20714 27384 20720 27396
rect 20579 27356 20720 27384
rect 20579 27353 20591 27356
rect 20533 27347 20591 27353
rect 20714 27344 20720 27356
rect 20772 27344 20778 27396
rect 23658 27384 23664 27396
rect 23598 27356 23664 27384
rect 23658 27344 23664 27356
rect 23716 27344 23722 27396
rect 24949 27387 25007 27393
rect 24949 27353 24961 27387
rect 24995 27384 25007 27387
rect 26068 27384 26096 27492
rect 26510 27480 26516 27532
rect 26568 27520 26574 27532
rect 26973 27523 27031 27529
rect 26973 27520 26985 27523
rect 26568 27492 26985 27520
rect 26568 27480 26574 27492
rect 26973 27489 26985 27492
rect 27019 27489 27031 27523
rect 26973 27483 27031 27489
rect 26694 27452 26700 27464
rect 26655 27424 26700 27452
rect 26694 27412 26700 27424
rect 26752 27412 26758 27464
rect 27448 27461 27476 27560
rect 28442 27548 28448 27600
rect 28500 27548 28506 27600
rect 28534 27548 28540 27600
rect 28592 27548 28598 27600
rect 28810 27548 28816 27600
rect 28868 27588 28874 27600
rect 29270 27588 29276 27600
rect 28868 27560 29276 27588
rect 28868 27548 28874 27560
rect 29270 27548 29276 27560
rect 29328 27548 29334 27600
rect 26789 27455 26847 27461
rect 26789 27421 26801 27455
rect 26835 27421 26847 27455
rect 26789 27415 26847 27421
rect 27433 27455 27491 27461
rect 27433 27421 27445 27455
rect 27479 27421 27491 27455
rect 27433 27415 27491 27421
rect 26804 27384 26832 27415
rect 28166 27412 28172 27464
rect 28224 27430 28230 27464
rect 28460 27463 28488 27548
rect 28552 27520 28580 27548
rect 28629 27523 28687 27529
rect 28629 27520 28641 27523
rect 28552 27492 28641 27520
rect 28629 27489 28641 27492
rect 28675 27489 28687 27523
rect 28629 27483 28687 27489
rect 28948 27480 28954 27532
rect 29006 27520 29012 27532
rect 29546 27520 29552 27532
rect 29006 27492 29552 27520
rect 29006 27480 29012 27492
rect 29546 27480 29552 27492
rect 29604 27480 29610 27532
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27520 46351 27523
rect 47026 27520 47032 27532
rect 46339 27492 47032 27520
rect 46339 27489 46351 27492
rect 46293 27483 46351 27489
rect 47026 27480 47032 27492
rect 47084 27480 47090 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 28433 27457 28491 27463
rect 28261 27433 28319 27439
rect 28261 27430 28273 27433
rect 28224 27412 28273 27430
rect 28184 27402 28273 27412
rect 28261 27399 28273 27402
rect 28307 27399 28319 27433
rect 28433 27423 28445 27457
rect 28479 27423 28491 27457
rect 28433 27417 28491 27423
rect 28534 27412 28540 27464
rect 28592 27452 28598 27464
rect 28813 27455 28871 27461
rect 28592 27424 28637 27452
rect 28592 27412 28598 27424
rect 28813 27421 28825 27455
rect 28859 27421 28871 27455
rect 28813 27415 28871 27421
rect 30193 27455 30251 27461
rect 30193 27421 30205 27455
rect 30239 27452 30251 27455
rect 30834 27452 30840 27464
rect 30239 27424 30840 27452
rect 30239 27421 30251 27424
rect 30193 27415 30251 27421
rect 28261 27393 28319 27399
rect 28828 27384 28856 27415
rect 30208 27384 30236 27415
rect 30834 27412 30840 27424
rect 30892 27412 30898 27464
rect 24995 27356 25636 27384
rect 26068 27356 26832 27384
rect 28736 27356 28856 27384
rect 28920 27356 30236 27384
rect 46477 27387 46535 27393
rect 24995 27353 25007 27356
rect 24949 27347 25007 27353
rect 25608 27328 25636 27356
rect 10778 27276 10784 27328
rect 10836 27316 10842 27328
rect 11241 27319 11299 27325
rect 11241 27316 11253 27319
rect 10836 27288 11253 27316
rect 10836 27276 10842 27288
rect 11241 27285 11253 27288
rect 11287 27285 11299 27319
rect 12066 27316 12072 27328
rect 12027 27288 12072 27316
rect 11241 27279 11299 27285
rect 12066 27276 12072 27288
rect 12124 27276 12130 27328
rect 14182 27316 14188 27328
rect 14143 27288 14188 27316
rect 14182 27276 14188 27288
rect 14240 27276 14246 27328
rect 25590 27276 25596 27328
rect 25648 27276 25654 27328
rect 25682 27276 25688 27328
rect 25740 27316 25746 27328
rect 26145 27319 26203 27325
rect 26145 27316 26157 27319
rect 25740 27288 26157 27316
rect 25740 27276 25746 27288
rect 26145 27285 26157 27288
rect 26191 27285 26203 27319
rect 26145 27279 26203 27285
rect 27617 27319 27675 27325
rect 27617 27285 27629 27319
rect 27663 27316 27675 27319
rect 27890 27316 27896 27328
rect 27663 27288 27896 27316
rect 27663 27285 27675 27288
rect 27617 27279 27675 27285
rect 27890 27276 27896 27288
rect 27948 27276 27954 27328
rect 28442 27276 28448 27328
rect 28500 27316 28506 27328
rect 28736 27316 28764 27356
rect 28920 27328 28948 27356
rect 46477 27353 46489 27387
rect 46523 27384 46535 27387
rect 47670 27384 47676 27396
rect 46523 27356 47676 27384
rect 46523 27353 46535 27356
rect 46477 27347 46535 27353
rect 47670 27344 47676 27356
rect 47728 27344 47734 27396
rect 28500 27288 28764 27316
rect 28500 27276 28506 27288
rect 28902 27276 28908 27328
rect 28960 27276 28966 27328
rect 28997 27319 29055 27325
rect 28997 27285 29009 27319
rect 29043 27316 29055 27319
rect 29362 27316 29368 27328
rect 29043 27288 29368 27316
rect 29043 27285 29055 27288
rect 28997 27279 29055 27285
rect 29362 27276 29368 27288
rect 29420 27276 29426 27328
rect 30285 27319 30343 27325
rect 30285 27285 30297 27319
rect 30331 27316 30343 27319
rect 30374 27316 30380 27328
rect 30331 27288 30380 27316
rect 30331 27285 30343 27288
rect 30285 27279 30343 27285
rect 30374 27276 30380 27288
rect 30432 27276 30438 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 11514 27072 11520 27124
rect 11572 27112 11578 27124
rect 11977 27115 12035 27121
rect 11977 27112 11989 27115
rect 11572 27084 11989 27112
rect 11572 27072 11578 27084
rect 11977 27081 11989 27084
rect 12023 27081 12035 27115
rect 11977 27075 12035 27081
rect 12161 27115 12219 27121
rect 12161 27081 12173 27115
rect 12207 27112 12219 27115
rect 12434 27112 12440 27124
rect 12207 27084 12440 27112
rect 12207 27081 12219 27084
rect 12161 27075 12219 27081
rect 11422 27004 11428 27056
rect 11480 27044 11486 27056
rect 11698 27044 11704 27056
rect 11480 27016 11704 27044
rect 11480 27004 11486 27016
rect 11698 27004 11704 27016
rect 11756 27044 11762 27056
rect 11885 27047 11943 27053
rect 11885 27044 11897 27047
rect 11756 27016 11897 27044
rect 11756 27004 11762 27016
rect 11885 27013 11897 27016
rect 11931 27013 11943 27047
rect 11992 27044 12020 27075
rect 12434 27072 12440 27084
rect 12492 27112 12498 27124
rect 13078 27112 13084 27124
rect 12492 27084 13084 27112
rect 12492 27072 12498 27084
rect 13078 27072 13084 27084
rect 13136 27072 13142 27124
rect 13170 27072 13176 27124
rect 13228 27112 13234 27124
rect 14645 27115 14703 27121
rect 14645 27112 14657 27115
rect 13228 27084 14657 27112
rect 13228 27072 13234 27084
rect 14645 27081 14657 27084
rect 14691 27081 14703 27115
rect 27982 27112 27988 27124
rect 14645 27075 14703 27081
rect 18248 27084 22508 27112
rect 27943 27084 27988 27112
rect 13446 27044 13452 27056
rect 11992 27016 13452 27044
rect 11885 27007 11943 27013
rect 13446 27004 13452 27016
rect 13504 27004 13510 27056
rect 14182 27004 14188 27056
rect 14240 27004 14246 27056
rect 18248 27053 18276 27084
rect 18233 27047 18291 27053
rect 18233 27044 18245 27047
rect 15764 27016 18245 27044
rect 10502 26976 10508 26988
rect 10463 26948 10508 26976
rect 10502 26936 10508 26948
rect 10560 26936 10566 26988
rect 11793 26979 11851 26985
rect 11793 26945 11805 26979
rect 11839 26976 11851 26979
rect 11974 26976 11980 26988
rect 11839 26948 11980 26976
rect 11839 26945 11851 26948
rect 11793 26939 11851 26945
rect 11974 26936 11980 26948
rect 12032 26936 12038 26988
rect 15764 26985 15792 27016
rect 18233 27013 18245 27016
rect 18279 27013 18291 27047
rect 18233 27007 18291 27013
rect 21818 27004 21824 27056
rect 21876 27044 21882 27056
rect 22480 27053 22508 27084
rect 27982 27072 27988 27084
rect 28040 27072 28046 27124
rect 28534 27072 28540 27124
rect 28592 27112 28598 27124
rect 30837 27115 30895 27121
rect 30837 27112 30849 27115
rect 28592 27084 30849 27112
rect 28592 27072 28598 27084
rect 30837 27081 30849 27084
rect 30883 27081 30895 27115
rect 30837 27075 30895 27081
rect 45830 27072 45836 27124
rect 45888 27112 45894 27124
rect 46198 27112 46204 27124
rect 45888 27084 46204 27112
rect 45888 27072 45894 27084
rect 46198 27072 46204 27084
rect 46256 27072 46262 27124
rect 22281 27047 22339 27053
rect 22281 27044 22293 27047
rect 21876 27016 22293 27044
rect 21876 27004 21882 27016
rect 22281 27013 22293 27016
rect 22327 27013 22339 27047
rect 22281 27007 22339 27013
rect 22465 27047 22523 27053
rect 22465 27013 22477 27047
rect 22511 27044 22523 27047
rect 24026 27044 24032 27056
rect 22511 27016 24032 27044
rect 22511 27013 22523 27016
rect 22465 27007 22523 27013
rect 24026 27004 24032 27016
rect 24084 27004 24090 27056
rect 26602 27044 26608 27056
rect 25884 27016 26608 27044
rect 15749 26979 15807 26985
rect 15749 26945 15761 26979
rect 15795 26945 15807 26979
rect 15749 26939 15807 26945
rect 15838 26936 15844 26988
rect 15896 26976 15902 26988
rect 15933 26979 15991 26985
rect 15933 26976 15945 26979
rect 15896 26948 15945 26976
rect 15896 26936 15902 26948
rect 15933 26945 15945 26948
rect 15979 26945 15991 26979
rect 20254 26976 20260 26988
rect 20215 26948 20260 26976
rect 15933 26939 15991 26945
rect 20254 26936 20260 26948
rect 20312 26936 20318 26988
rect 20441 26979 20499 26985
rect 20441 26945 20453 26979
rect 20487 26976 20499 26979
rect 20530 26976 20536 26988
rect 20487 26948 20536 26976
rect 20487 26945 20499 26948
rect 20441 26939 20499 26945
rect 20530 26936 20536 26948
rect 20588 26936 20594 26988
rect 20717 26979 20775 26985
rect 20717 26945 20729 26979
rect 20763 26976 20775 26979
rect 21082 26976 21088 26988
rect 20763 26948 21088 26976
rect 20763 26945 20775 26948
rect 20717 26939 20775 26945
rect 21082 26936 21088 26948
rect 21140 26936 21146 26988
rect 25682 26976 25688 26988
rect 25643 26948 25688 26976
rect 25682 26936 25688 26948
rect 25740 26936 25746 26988
rect 25884 26985 25912 27016
rect 26602 27004 26608 27016
rect 26660 27004 26666 27056
rect 28442 27044 28448 27056
rect 27816 27016 28448 27044
rect 25869 26979 25927 26985
rect 25869 26945 25881 26979
rect 25915 26945 25927 26979
rect 26234 26976 26240 26988
rect 26195 26948 26240 26976
rect 25869 26939 25927 26945
rect 26234 26936 26240 26948
rect 26292 26976 26298 26988
rect 27816 26976 27844 27016
rect 28442 27004 28448 27016
rect 28500 27004 28506 27056
rect 29362 27044 29368 27056
rect 29323 27016 29368 27044
rect 29362 27004 29368 27016
rect 29420 27004 29426 27056
rect 30374 27004 30380 27056
rect 30432 27004 30438 27056
rect 26292 26948 27844 26976
rect 26292 26936 26298 26948
rect 27890 26936 27896 26988
rect 27948 26976 27954 26988
rect 28810 26976 28816 26988
rect 27948 26948 28816 26976
rect 27948 26936 27954 26948
rect 28810 26936 28816 26948
rect 28868 26936 28874 26988
rect 29086 26976 29092 26988
rect 29047 26948 29092 26976
rect 29086 26936 29092 26948
rect 29144 26936 29150 26988
rect 45830 26936 45836 26988
rect 45888 26976 45894 26988
rect 46109 26979 46167 26985
rect 46109 26976 46121 26979
rect 45888 26948 46121 26976
rect 45888 26936 45894 26948
rect 46109 26945 46121 26948
rect 46155 26945 46167 26979
rect 46109 26939 46167 26945
rect 12897 26911 12955 26917
rect 12897 26877 12909 26911
rect 12943 26877 12955 26911
rect 13170 26908 13176 26920
rect 13131 26880 13176 26908
rect 12897 26871 12955 26877
rect 11609 26843 11667 26849
rect 11609 26809 11621 26843
rect 11655 26840 11667 26843
rect 11882 26840 11888 26852
rect 11655 26812 11888 26840
rect 11655 26809 11667 26812
rect 11609 26803 11667 26809
rect 11882 26800 11888 26812
rect 11940 26840 11946 26852
rect 12250 26840 12256 26852
rect 11940 26812 12256 26840
rect 11940 26800 11946 26812
rect 12250 26800 12256 26812
rect 12308 26800 12314 26852
rect 10502 26772 10508 26784
rect 10463 26744 10508 26772
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 12912 26772 12940 26871
rect 13170 26868 13176 26880
rect 13228 26868 13234 26920
rect 19981 26911 20039 26917
rect 19981 26877 19993 26911
rect 20027 26908 20039 26911
rect 20806 26908 20812 26920
rect 20027 26880 20812 26908
rect 20027 26877 20039 26880
rect 19981 26871 20039 26877
rect 20806 26868 20812 26880
rect 20864 26868 20870 26920
rect 25590 26868 25596 26920
rect 25648 26908 25654 26920
rect 25961 26911 26019 26917
rect 25961 26908 25973 26911
rect 25648 26880 25973 26908
rect 25648 26868 25654 26880
rect 25961 26877 25973 26880
rect 26007 26877 26019 26911
rect 25961 26871 26019 26877
rect 20349 26843 20407 26849
rect 20349 26809 20361 26843
rect 20395 26840 20407 26843
rect 20714 26840 20720 26852
rect 20395 26812 20720 26840
rect 20395 26809 20407 26812
rect 20349 26803 20407 26809
rect 20714 26800 20720 26812
rect 20772 26840 20778 26852
rect 21266 26840 21272 26852
rect 20772 26812 21272 26840
rect 20772 26800 20778 26812
rect 21266 26800 21272 26812
rect 21324 26800 21330 26852
rect 25976 26840 26004 26871
rect 26050 26868 26056 26920
rect 26108 26908 26114 26920
rect 26108 26880 26153 26908
rect 26108 26868 26114 26880
rect 32122 26868 32128 26920
rect 32180 26908 32186 26920
rect 46385 26911 46443 26917
rect 46385 26908 46397 26911
rect 32180 26880 46397 26908
rect 32180 26868 32186 26880
rect 46385 26877 46397 26880
rect 46431 26908 46443 26911
rect 47486 26908 47492 26920
rect 46431 26880 47492 26908
rect 46431 26877 46443 26880
rect 46385 26871 46443 26877
rect 47486 26868 47492 26880
rect 47544 26868 47550 26920
rect 26694 26840 26700 26852
rect 25976 26812 26700 26840
rect 26694 26800 26700 26812
rect 26752 26800 26758 26852
rect 13814 26772 13820 26784
rect 12912 26744 13820 26772
rect 13814 26732 13820 26744
rect 13872 26732 13878 26784
rect 16114 26772 16120 26784
rect 16075 26744 16120 26772
rect 16114 26732 16120 26744
rect 16172 26732 16178 26784
rect 18230 26732 18236 26784
rect 18288 26772 18294 26784
rect 18325 26775 18383 26781
rect 18325 26772 18337 26775
rect 18288 26744 18337 26772
rect 18288 26732 18294 26744
rect 18325 26741 18337 26744
rect 18371 26741 18383 26775
rect 18325 26735 18383 26741
rect 20438 26732 20444 26784
rect 20496 26772 20502 26784
rect 20533 26775 20591 26781
rect 20533 26772 20545 26775
rect 20496 26744 20545 26772
rect 20496 26732 20502 26744
rect 20533 26741 20545 26744
rect 20579 26741 20591 26775
rect 26418 26772 26424 26784
rect 26379 26744 26424 26772
rect 20533 26735 20591 26741
rect 26418 26732 26424 26744
rect 26476 26732 26482 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 12250 26568 12256 26580
rect 12211 26540 12256 26568
rect 12250 26528 12256 26540
rect 12308 26528 12314 26580
rect 23658 26568 23664 26580
rect 21560 26540 22692 26568
rect 23619 26540 23664 26568
rect 16114 26500 16120 26512
rect 14108 26472 16120 26500
rect 10502 26432 10508 26444
rect 10463 26404 10508 26432
rect 10502 26392 10508 26404
rect 10560 26392 10566 26444
rect 10778 26432 10784 26444
rect 10739 26404 10784 26432
rect 10778 26392 10784 26404
rect 10836 26392 10842 26444
rect 13446 26392 13452 26444
rect 13504 26432 13510 26444
rect 14108 26432 14136 26472
rect 13504 26404 14136 26432
rect 13504 26392 13510 26404
rect 13173 26367 13231 26373
rect 13173 26364 13185 26367
rect 12406 26336 13185 26364
rect 12066 26296 12072 26308
rect 12006 26268 12072 26296
rect 12066 26256 12072 26268
rect 12124 26256 12130 26308
rect 12250 26256 12256 26308
rect 12308 26296 12314 26308
rect 12406 26296 12434 26336
rect 13173 26333 13185 26336
rect 13219 26333 13231 26367
rect 13173 26327 13231 26333
rect 13262 26324 13268 26376
rect 13320 26364 13326 26376
rect 14108 26373 14136 26404
rect 15580 26373 15608 26472
rect 16114 26460 16120 26472
rect 16172 26460 16178 26512
rect 16209 26503 16267 26509
rect 16209 26469 16221 26503
rect 16255 26469 16267 26503
rect 16209 26463 16267 26469
rect 16224 26432 16252 26463
rect 16224 26404 16988 26432
rect 14093 26367 14151 26373
rect 13320 26336 13365 26364
rect 13320 26324 13326 26336
rect 14093 26333 14105 26367
rect 14139 26333 14151 26367
rect 14093 26327 14151 26333
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26333 14335 26367
rect 14277 26327 14335 26333
rect 15565 26367 15623 26373
rect 15565 26333 15577 26367
rect 15611 26333 15623 26367
rect 15746 26364 15752 26376
rect 15707 26336 15752 26364
rect 15565 26327 15623 26333
rect 12986 26296 12992 26308
rect 12308 26268 12434 26296
rect 12947 26268 12992 26296
rect 12308 26256 12314 26268
rect 12986 26256 12992 26268
rect 13044 26256 13050 26308
rect 13446 26256 13452 26308
rect 13504 26296 13510 26308
rect 14185 26299 14243 26305
rect 14185 26296 14197 26299
rect 13504 26268 14197 26296
rect 13504 26256 13510 26268
rect 14185 26265 14197 26268
rect 14231 26265 14243 26299
rect 14185 26259 14243 26265
rect 11422 26188 11428 26240
rect 11480 26228 11486 26240
rect 13357 26231 13415 26237
rect 13357 26228 13369 26231
rect 11480 26200 13369 26228
rect 11480 26188 11486 26200
rect 13357 26197 13369 26200
rect 13403 26197 13415 26231
rect 13357 26191 13415 26197
rect 13541 26231 13599 26237
rect 13541 26197 13553 26231
rect 13587 26228 13599 26231
rect 14292 26228 14320 26327
rect 15746 26324 15752 26336
rect 15804 26364 15810 26376
rect 16960 26373 16988 26404
rect 16485 26367 16543 26373
rect 16485 26364 16497 26367
rect 15804 26336 16497 26364
rect 15804 26324 15810 26336
rect 16485 26333 16497 26336
rect 16531 26333 16543 26367
rect 16485 26327 16543 26333
rect 16945 26367 17003 26373
rect 16945 26333 16957 26367
rect 16991 26333 17003 26367
rect 16945 26327 17003 26333
rect 17129 26367 17187 26373
rect 17129 26333 17141 26367
rect 17175 26364 17187 26367
rect 20806 26364 20812 26376
rect 17175 26336 20812 26364
rect 17175 26333 17187 26336
rect 17129 26327 17187 26333
rect 20806 26324 20812 26336
rect 20864 26324 20870 26376
rect 21450 26324 21456 26376
rect 21508 26364 21514 26376
rect 21560 26373 21588 26540
rect 21729 26503 21787 26509
rect 21729 26469 21741 26503
rect 21775 26500 21787 26503
rect 21910 26500 21916 26512
rect 21775 26472 21916 26500
rect 21775 26469 21787 26472
rect 21729 26463 21787 26469
rect 21910 26460 21916 26472
rect 21968 26500 21974 26512
rect 22465 26503 22523 26509
rect 22465 26500 22477 26503
rect 21968 26472 22477 26500
rect 21968 26460 21974 26472
rect 22465 26469 22477 26472
rect 22511 26469 22523 26503
rect 22465 26463 22523 26469
rect 22664 26441 22692 26540
rect 23658 26528 23664 26540
rect 23716 26528 23722 26580
rect 26234 26500 26240 26512
rect 26195 26472 26240 26500
rect 26234 26460 26240 26472
rect 26292 26460 26298 26512
rect 22649 26435 22707 26441
rect 21652 26404 22094 26432
rect 21652 26376 21680 26404
rect 21545 26367 21603 26373
rect 21545 26364 21557 26367
rect 21508 26336 21557 26364
rect 21508 26324 21514 26336
rect 21545 26333 21557 26336
rect 21591 26333 21603 26367
rect 21545 26327 21603 26333
rect 21634 26324 21640 26376
rect 21692 26364 21698 26376
rect 21692 26336 21737 26364
rect 21692 26324 21698 26336
rect 21818 26324 21824 26376
rect 21876 26364 21882 26376
rect 22066 26364 22094 26404
rect 22649 26401 22661 26435
rect 22695 26401 22707 26435
rect 24578 26432 24584 26444
rect 22649 26395 22707 26401
rect 23124 26404 24584 26432
rect 22373 26367 22431 26373
rect 22373 26364 22385 26367
rect 21876 26336 21921 26364
rect 22066 26336 22385 26364
rect 21876 26324 21882 26336
rect 22373 26333 22385 26336
rect 22419 26364 22431 26367
rect 23124 26364 23152 26404
rect 24578 26392 24584 26404
rect 24636 26392 24642 26444
rect 45002 26392 45008 26444
rect 45060 26432 45066 26444
rect 45465 26435 45523 26441
rect 45465 26432 45477 26435
rect 45060 26404 45477 26432
rect 45060 26392 45066 26404
rect 45465 26401 45477 26404
rect 45511 26432 45523 26435
rect 46382 26432 46388 26444
rect 45511 26404 46388 26432
rect 45511 26401 45523 26404
rect 45465 26395 45523 26401
rect 46382 26392 46388 26404
rect 46440 26392 46446 26444
rect 48038 26432 48044 26444
rect 47999 26404 48044 26432
rect 48038 26392 48044 26404
rect 48096 26392 48102 26444
rect 22419 26336 23152 26364
rect 22419 26333 22431 26336
rect 22373 26327 22431 26333
rect 23198 26324 23204 26376
rect 23256 26364 23262 26376
rect 23569 26367 23627 26373
rect 23569 26364 23581 26367
rect 23256 26336 23581 26364
rect 23256 26324 23262 26336
rect 23569 26333 23581 26336
rect 23615 26333 23627 26367
rect 23569 26327 23627 26333
rect 45097 26367 45155 26373
rect 45097 26333 45109 26367
rect 45143 26364 45155 26367
rect 45830 26364 45836 26376
rect 45143 26336 45836 26364
rect 45143 26333 45155 26336
rect 45097 26327 45155 26333
rect 45830 26324 45836 26336
rect 45888 26324 45894 26376
rect 46014 26324 46020 26376
rect 46072 26364 46078 26376
rect 46201 26367 46259 26373
rect 46201 26364 46213 26367
rect 46072 26336 46213 26364
rect 46072 26324 46078 26336
rect 46201 26333 46213 26336
rect 46247 26333 46259 26367
rect 46201 26327 46259 26333
rect 16206 26296 16212 26308
rect 16167 26268 16212 26296
rect 16206 26256 16212 26268
rect 16264 26256 16270 26308
rect 21361 26299 21419 26305
rect 21361 26265 21373 26299
rect 21407 26296 21419 26299
rect 22278 26296 22284 26308
rect 21407 26268 22284 26296
rect 21407 26265 21419 26268
rect 21361 26259 21419 26265
rect 22278 26256 22284 26268
rect 22336 26256 22342 26308
rect 26053 26299 26111 26305
rect 26053 26296 26065 26299
rect 22572 26268 26065 26296
rect 15930 26228 15936 26240
rect 13587 26200 15936 26228
rect 13587 26197 13599 26200
rect 13541 26191 13599 26197
rect 15930 26188 15936 26200
rect 15988 26188 15994 26240
rect 16390 26228 16396 26240
rect 16351 26200 16396 26228
rect 16390 26188 16396 26200
rect 16448 26188 16454 26240
rect 17034 26228 17040 26240
rect 16995 26200 17040 26228
rect 17034 26188 17040 26200
rect 17092 26188 17098 26240
rect 18874 26188 18880 26240
rect 18932 26228 18938 26240
rect 20990 26228 20996 26240
rect 18932 26200 20996 26228
rect 18932 26188 18938 26200
rect 20990 26188 20996 26200
rect 21048 26188 21054 26240
rect 22186 26188 22192 26240
rect 22244 26228 22250 26240
rect 22572 26228 22600 26268
rect 26053 26265 26065 26268
rect 26099 26265 26111 26299
rect 46382 26296 46388 26308
rect 46343 26268 46388 26296
rect 26053 26259 26111 26265
rect 46382 26256 46388 26268
rect 46440 26256 46446 26308
rect 22244 26200 22600 26228
rect 22649 26231 22707 26237
rect 22244 26188 22250 26200
rect 22649 26197 22661 26231
rect 22695 26228 22707 26231
rect 22830 26228 22836 26240
rect 22695 26200 22836 26228
rect 22695 26197 22707 26200
rect 22649 26191 22707 26197
rect 22830 26188 22836 26200
rect 22888 26188 22894 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 11146 25984 11152 26036
rect 11204 26024 11210 26036
rect 11793 26027 11851 26033
rect 11793 26024 11805 26027
rect 11204 25996 11805 26024
rect 11204 25984 11210 25996
rect 11793 25993 11805 25996
rect 11839 25993 11851 26027
rect 11793 25987 11851 25993
rect 12805 26027 12863 26033
rect 12805 25993 12817 26027
rect 12851 26024 12863 26027
rect 13170 26024 13176 26036
rect 12851 25996 13176 26024
rect 12851 25993 12863 25996
rect 12805 25987 12863 25993
rect 13170 25984 13176 25996
rect 13228 25984 13234 26036
rect 13814 26024 13820 26036
rect 13775 25996 13820 26024
rect 13814 25984 13820 25996
rect 13872 25984 13878 26036
rect 15933 26027 15991 26033
rect 15933 25993 15945 26027
rect 15979 26024 15991 26027
rect 16390 26024 16396 26036
rect 15979 25996 16396 26024
rect 15979 25993 15991 25996
rect 15933 25987 15991 25993
rect 16390 25984 16396 25996
rect 16448 25984 16454 26036
rect 20254 26024 20260 26036
rect 16868 25996 20260 26024
rect 11422 25916 11428 25968
rect 11480 25956 11486 25968
rect 11609 25959 11667 25965
rect 11609 25956 11621 25959
rect 11480 25928 11621 25956
rect 11480 25916 11486 25928
rect 11609 25925 11621 25928
rect 11655 25925 11667 25959
rect 13446 25956 13452 25968
rect 11609 25919 11667 25925
rect 13004 25928 13452 25956
rect 9493 25891 9551 25897
rect 9493 25857 9505 25891
rect 9539 25888 9551 25891
rect 10410 25888 10416 25900
rect 9539 25860 10416 25888
rect 9539 25857 9551 25860
rect 9493 25851 9551 25857
rect 10410 25848 10416 25860
rect 10468 25848 10474 25900
rect 10962 25848 10968 25900
rect 11020 25888 11026 25900
rect 11517 25891 11575 25897
rect 11517 25888 11529 25891
rect 11020 25860 11529 25888
rect 11020 25848 11026 25860
rect 11517 25857 11529 25860
rect 11563 25857 11575 25891
rect 11882 25888 11888 25900
rect 11843 25860 11888 25888
rect 11517 25851 11575 25857
rect 11882 25848 11888 25860
rect 11940 25848 11946 25900
rect 12802 25848 12808 25900
rect 12860 25888 12866 25900
rect 13004 25897 13032 25928
rect 13446 25916 13452 25928
rect 13504 25916 13510 25968
rect 15654 25916 15660 25968
rect 15712 25956 15718 25968
rect 15841 25959 15899 25965
rect 15841 25956 15853 25959
rect 15712 25928 15853 25956
rect 15712 25916 15718 25928
rect 15841 25925 15853 25928
rect 15887 25925 15899 25959
rect 15841 25919 15899 25925
rect 16117 25959 16175 25965
rect 16117 25925 16129 25959
rect 16163 25956 16175 25959
rect 16868 25956 16896 25996
rect 20254 25984 20260 25996
rect 20312 25984 20318 26036
rect 21266 26024 21272 26036
rect 21227 25996 21272 26024
rect 21266 25984 21272 25996
rect 21324 25984 21330 26036
rect 22278 26024 22284 26036
rect 22239 25996 22284 26024
rect 22278 25984 22284 25996
rect 22336 25984 22342 26036
rect 22370 25984 22376 26036
rect 22428 26024 22434 26036
rect 27430 26024 27436 26036
rect 22428 25996 27436 26024
rect 22428 25984 22434 25996
rect 27430 25984 27436 25996
rect 27488 25984 27494 26036
rect 44729 26027 44787 26033
rect 44729 25993 44741 26027
rect 44775 26024 44787 26027
rect 46382 26024 46388 26036
rect 44775 25996 46388 26024
rect 44775 25993 44787 25996
rect 44729 25987 44787 25993
rect 46382 25984 46388 25996
rect 46440 25984 46446 26036
rect 46658 25984 46664 26036
rect 46716 26024 46722 26036
rect 46753 26027 46811 26033
rect 46753 26024 46765 26027
rect 46716 25996 46765 26024
rect 46716 25984 46722 25996
rect 46753 25993 46765 25996
rect 46799 26024 46811 26027
rect 47578 26024 47584 26036
rect 46799 25996 47584 26024
rect 46799 25993 46811 25996
rect 46753 25987 46811 25993
rect 47578 25984 47584 25996
rect 47636 25984 47642 26036
rect 16163 25928 16896 25956
rect 16945 25959 17003 25965
rect 16163 25925 16175 25928
rect 16117 25919 16175 25925
rect 16945 25925 16957 25959
rect 16991 25956 17003 25959
rect 17034 25956 17040 25968
rect 16991 25928 17040 25956
rect 16991 25925 17003 25928
rect 16945 25919 17003 25925
rect 17034 25916 17040 25928
rect 17092 25916 17098 25968
rect 17954 25916 17960 25968
rect 18012 25916 18018 25968
rect 20990 25916 20996 25968
rect 21048 25956 21054 25968
rect 21085 25959 21143 25965
rect 21085 25956 21097 25959
rect 21048 25928 21097 25956
rect 21048 25916 21054 25928
rect 21085 25925 21097 25928
rect 21131 25956 21143 25959
rect 21818 25956 21824 25968
rect 21131 25928 21824 25956
rect 21131 25925 21143 25928
rect 21085 25919 21143 25925
rect 21818 25916 21824 25928
rect 21876 25916 21882 25968
rect 12989 25891 13047 25897
rect 12989 25888 13001 25891
rect 12860 25860 13001 25888
rect 12860 25848 12866 25860
rect 12989 25857 13001 25860
rect 13035 25857 13047 25891
rect 12989 25851 13047 25857
rect 13078 25848 13084 25900
rect 13136 25888 13142 25900
rect 13173 25891 13231 25897
rect 13173 25888 13185 25891
rect 13136 25860 13185 25888
rect 13136 25848 13142 25860
rect 13173 25857 13185 25860
rect 13219 25857 13231 25891
rect 13173 25851 13231 25857
rect 13725 25891 13783 25897
rect 13725 25857 13737 25891
rect 13771 25888 13783 25891
rect 13998 25888 14004 25900
rect 13771 25860 14004 25888
rect 13771 25857 13783 25860
rect 13725 25851 13783 25857
rect 13998 25848 14004 25860
rect 14056 25848 14062 25900
rect 15562 25848 15568 25900
rect 15620 25888 15626 25900
rect 15749 25891 15807 25897
rect 15749 25888 15761 25891
rect 15620 25860 15761 25888
rect 15620 25848 15626 25860
rect 15749 25857 15761 25860
rect 15795 25857 15807 25891
rect 18874 25888 18880 25900
rect 18835 25860 18880 25888
rect 15749 25851 15807 25857
rect 18874 25848 18880 25860
rect 18932 25848 18938 25900
rect 19797 25891 19855 25897
rect 19797 25857 19809 25891
rect 19843 25857 19855 25891
rect 19797 25851 19855 25857
rect 11701 25823 11759 25829
rect 11701 25789 11713 25823
rect 11747 25820 11759 25823
rect 11974 25820 11980 25832
rect 11747 25792 11980 25820
rect 11747 25789 11759 25792
rect 11701 25783 11759 25789
rect 11974 25780 11980 25792
rect 12032 25780 12038 25832
rect 13265 25823 13323 25829
rect 13265 25789 13277 25823
rect 13311 25789 13323 25823
rect 13265 25783 13323 25789
rect 12986 25712 12992 25764
rect 13044 25752 13050 25764
rect 13280 25752 13308 25783
rect 16574 25780 16580 25832
rect 16632 25820 16638 25832
rect 16669 25823 16727 25829
rect 16669 25820 16681 25823
rect 16632 25792 16681 25820
rect 16632 25780 16638 25792
rect 16669 25789 16681 25792
rect 16715 25789 16727 25823
rect 19812 25820 19840 25851
rect 19978 25848 19984 25900
rect 20036 25888 20042 25900
rect 20257 25891 20315 25897
rect 20257 25888 20269 25891
rect 20036 25860 20269 25888
rect 20036 25848 20042 25860
rect 20257 25857 20269 25860
rect 20303 25857 20315 25891
rect 20257 25851 20315 25857
rect 20901 25891 20959 25897
rect 20901 25857 20913 25891
rect 20947 25888 20959 25891
rect 21450 25888 21456 25900
rect 20947 25860 21456 25888
rect 20947 25857 20959 25860
rect 20901 25851 20959 25857
rect 21450 25848 21456 25860
rect 21508 25888 21514 25900
rect 21910 25888 21916 25900
rect 21508 25860 21916 25888
rect 21508 25848 21514 25860
rect 21910 25848 21916 25860
rect 21968 25848 21974 25900
rect 22189 25891 22247 25897
rect 22189 25857 22201 25891
rect 22235 25888 22247 25891
rect 23106 25888 23112 25900
rect 22235 25860 23112 25888
rect 22235 25857 22247 25860
rect 22189 25851 22247 25857
rect 23106 25848 23112 25860
rect 23164 25848 23170 25900
rect 23198 25848 23204 25900
rect 23256 25888 23262 25900
rect 24489 25891 24547 25897
rect 24489 25888 24501 25891
rect 23256 25860 24501 25888
rect 23256 25848 23262 25860
rect 24489 25857 24501 25860
rect 24535 25888 24547 25891
rect 25501 25891 25559 25897
rect 25501 25888 25513 25891
rect 24535 25860 25513 25888
rect 24535 25857 24547 25860
rect 24489 25851 24547 25857
rect 25501 25857 25513 25860
rect 25547 25857 25559 25891
rect 25501 25851 25559 25857
rect 44637 25891 44695 25897
rect 44637 25857 44649 25891
rect 44683 25888 44695 25891
rect 45281 25891 45339 25897
rect 45281 25888 45293 25891
rect 44683 25860 45293 25888
rect 44683 25857 44695 25860
rect 44637 25851 44695 25857
rect 45281 25857 45293 25860
rect 45327 25888 45339 25891
rect 45830 25888 45836 25900
rect 45327 25860 45836 25888
rect 45327 25857 45339 25860
rect 45281 25851 45339 25857
rect 45830 25848 45836 25860
rect 45888 25888 45894 25900
rect 47581 25891 47639 25897
rect 47581 25888 47593 25891
rect 45888 25860 47593 25888
rect 45888 25848 45894 25860
rect 47581 25857 47593 25860
rect 47627 25857 47639 25891
rect 47581 25851 47639 25857
rect 19812 25792 21864 25820
rect 16669 25783 16727 25789
rect 13044 25724 13308 25752
rect 13044 25712 13050 25724
rect 14090 25712 14096 25764
rect 14148 25752 14154 25764
rect 15565 25755 15623 25761
rect 15565 25752 15577 25755
rect 14148 25724 15577 25752
rect 14148 25712 14154 25724
rect 15565 25721 15577 25724
rect 15611 25752 15623 25755
rect 16206 25752 16212 25764
rect 15611 25724 16212 25752
rect 15611 25721 15623 25724
rect 15565 25715 15623 25721
rect 16206 25712 16212 25724
rect 16264 25712 16270 25764
rect 19058 25752 19064 25764
rect 18971 25724 19064 25752
rect 19058 25712 19064 25724
rect 19116 25752 19122 25764
rect 19978 25752 19984 25764
rect 19116 25724 19984 25752
rect 19116 25712 19122 25724
rect 19978 25712 19984 25724
rect 20036 25712 20042 25764
rect 21836 25761 21864 25792
rect 22278 25780 22284 25832
rect 22336 25820 22342 25832
rect 22373 25823 22431 25829
rect 22373 25820 22385 25823
rect 22336 25792 22385 25820
rect 22336 25780 22342 25792
rect 22373 25789 22385 25792
rect 22419 25789 22431 25823
rect 22373 25783 22431 25789
rect 47210 25780 47216 25832
rect 47268 25820 47274 25832
rect 47765 25823 47823 25829
rect 47765 25820 47777 25823
rect 47268 25792 47777 25820
rect 47268 25780 47274 25792
rect 47765 25789 47777 25792
rect 47811 25789 47823 25823
rect 47765 25783 47823 25789
rect 21821 25755 21879 25761
rect 21821 25721 21833 25755
rect 21867 25721 21879 25755
rect 21821 25715 21879 25721
rect 9398 25644 9404 25696
rect 9456 25684 9462 25696
rect 9493 25687 9551 25693
rect 9493 25684 9505 25687
rect 9456 25656 9505 25684
rect 9456 25644 9462 25656
rect 9493 25653 9505 25656
rect 9539 25653 9551 25687
rect 16224 25684 16252 25712
rect 18417 25687 18475 25693
rect 18417 25684 18429 25687
rect 16224 25656 18429 25684
rect 9493 25647 9551 25653
rect 18417 25653 18429 25656
rect 18463 25653 18475 25687
rect 18417 25647 18475 25653
rect 19518 25644 19524 25696
rect 19576 25684 19582 25696
rect 19613 25687 19671 25693
rect 19613 25684 19625 25687
rect 19576 25656 19625 25684
rect 19576 25644 19582 25656
rect 19613 25653 19625 25656
rect 19659 25653 19671 25687
rect 19613 25647 19671 25653
rect 20254 25644 20260 25696
rect 20312 25684 20318 25696
rect 20349 25687 20407 25693
rect 20349 25684 20361 25687
rect 20312 25656 20361 25684
rect 20312 25644 20318 25656
rect 20349 25653 20361 25656
rect 20395 25653 20407 25687
rect 20349 25647 20407 25653
rect 24581 25687 24639 25693
rect 24581 25653 24593 25687
rect 24627 25684 24639 25687
rect 24854 25684 24860 25696
rect 24627 25656 24860 25684
rect 24627 25653 24639 25656
rect 24581 25647 24639 25653
rect 24854 25644 24860 25656
rect 24912 25644 24918 25696
rect 25593 25687 25651 25693
rect 25593 25653 25605 25687
rect 25639 25684 25651 25687
rect 26050 25684 26056 25696
rect 25639 25656 26056 25684
rect 25639 25653 25651 25656
rect 25593 25647 25651 25653
rect 26050 25644 26056 25656
rect 26108 25644 26114 25696
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 16574 25480 16580 25492
rect 16535 25452 16580 25480
rect 16574 25440 16580 25452
rect 16632 25440 16638 25492
rect 20990 25480 20996 25492
rect 20951 25452 20996 25480
rect 20990 25440 20996 25452
rect 21048 25440 21054 25492
rect 21634 25480 21640 25492
rect 21595 25452 21640 25480
rect 21634 25440 21640 25452
rect 21692 25440 21698 25492
rect 26694 25440 26700 25492
rect 26752 25480 26758 25492
rect 27065 25483 27123 25489
rect 27065 25480 27077 25483
rect 26752 25452 27077 25480
rect 26752 25440 26758 25452
rect 27065 25449 27077 25452
rect 27111 25449 27123 25483
rect 27065 25443 27123 25449
rect 18874 25412 18880 25424
rect 13556 25384 18880 25412
rect 9398 25344 9404 25356
rect 9359 25316 9404 25344
rect 9398 25304 9404 25316
rect 9456 25304 9462 25356
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 13357 25279 13415 25285
rect 13357 25245 13369 25279
rect 13403 25276 13415 25279
rect 13556 25276 13584 25384
rect 18874 25372 18880 25384
rect 18932 25372 18938 25424
rect 22002 25372 22008 25424
rect 22060 25372 22066 25424
rect 22186 25372 22192 25424
rect 22244 25412 22250 25424
rect 22649 25415 22707 25421
rect 22649 25412 22661 25415
rect 22244 25384 22661 25412
rect 22244 25372 22250 25384
rect 22649 25381 22661 25384
rect 22695 25381 22707 25415
rect 45830 25412 45836 25424
rect 45791 25384 45836 25412
rect 22649 25375 22707 25381
rect 45830 25372 45836 25384
rect 45888 25372 45894 25424
rect 13630 25304 13636 25356
rect 13688 25344 13694 25356
rect 15562 25344 15568 25356
rect 13688 25316 15568 25344
rect 13688 25304 13694 25316
rect 15562 25304 15568 25316
rect 15620 25304 15626 25356
rect 19242 25344 19248 25356
rect 19203 25316 19248 25344
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 19518 25344 19524 25356
rect 19479 25316 19524 25344
rect 19518 25304 19524 25316
rect 19576 25304 19582 25356
rect 21821 25347 21879 25353
rect 21821 25313 21833 25347
rect 21867 25344 21879 25347
rect 22020 25344 22048 25372
rect 21867 25316 22048 25344
rect 21867 25313 21879 25316
rect 21821 25307 21879 25313
rect 23474 25304 23480 25356
rect 23532 25344 23538 25356
rect 25317 25347 25375 25353
rect 25317 25344 25329 25347
rect 23532 25316 25329 25344
rect 23532 25304 23538 25316
rect 25317 25313 25329 25316
rect 25363 25344 25375 25347
rect 26970 25344 26976 25356
rect 25363 25316 26976 25344
rect 25363 25313 25375 25316
rect 25317 25307 25375 25313
rect 26970 25304 26976 25316
rect 27028 25304 27034 25356
rect 48130 25344 48136 25356
rect 48091 25316 48136 25344
rect 48130 25304 48136 25316
rect 48188 25304 48194 25356
rect 13403 25248 13584 25276
rect 13403 25245 13415 25248
rect 13357 25239 13415 25245
rect 13906 25236 13912 25288
rect 13964 25276 13970 25288
rect 14093 25279 14151 25285
rect 14093 25276 14105 25279
rect 13964 25248 14105 25276
rect 13964 25236 13970 25248
rect 14093 25245 14105 25248
rect 14139 25245 14151 25279
rect 14093 25239 14151 25245
rect 15654 25236 15660 25288
rect 15712 25276 15718 25288
rect 15749 25279 15807 25285
rect 15749 25276 15761 25279
rect 15712 25248 15761 25276
rect 15712 25236 15718 25248
rect 15749 25245 15761 25248
rect 15795 25245 15807 25279
rect 15749 25239 15807 25245
rect 16393 25279 16451 25285
rect 16393 25245 16405 25279
rect 16439 25245 16451 25279
rect 16393 25239 16451 25245
rect 1670 25208 1676 25220
rect 1631 25180 1676 25208
rect 1670 25168 1676 25180
rect 1728 25168 1734 25220
rect 9674 25208 9680 25220
rect 9635 25180 9680 25208
rect 9674 25168 9680 25180
rect 9732 25168 9738 25220
rect 10410 25168 10416 25220
rect 10468 25168 10474 25220
rect 11422 25208 11428 25220
rect 11383 25180 11428 25208
rect 11422 25168 11428 25180
rect 11480 25168 11486 25220
rect 13541 25211 13599 25217
rect 13541 25177 13553 25211
rect 13587 25208 13599 25211
rect 13722 25208 13728 25220
rect 13587 25180 13728 25208
rect 13587 25177 13599 25180
rect 13541 25171 13599 25177
rect 13722 25168 13728 25180
rect 13780 25168 13786 25220
rect 13998 25168 14004 25220
rect 14056 25208 14062 25220
rect 16408 25208 16436 25239
rect 20990 25236 20996 25288
rect 21048 25276 21054 25288
rect 21545 25279 21603 25285
rect 21545 25276 21557 25279
rect 21048 25248 21557 25276
rect 21048 25236 21054 25248
rect 21545 25245 21557 25248
rect 21591 25245 21603 25279
rect 21545 25239 21603 25245
rect 21910 25236 21916 25288
rect 21968 25276 21974 25288
rect 22005 25279 22063 25285
rect 22005 25276 22017 25279
rect 21968 25248 22017 25276
rect 21968 25236 21974 25248
rect 22005 25245 22017 25248
rect 22051 25245 22063 25279
rect 22925 25279 22983 25285
rect 22925 25276 22937 25279
rect 22005 25239 22063 25245
rect 22204 25248 22937 25276
rect 16574 25208 16580 25220
rect 14056 25180 16580 25208
rect 14056 25168 14062 25180
rect 16574 25168 16580 25180
rect 16632 25168 16638 25220
rect 20254 25168 20260 25220
rect 20312 25168 20318 25220
rect 14090 25100 14096 25152
rect 14148 25140 14154 25152
rect 14185 25143 14243 25149
rect 14185 25140 14197 25143
rect 14148 25112 14197 25140
rect 14148 25100 14154 25112
rect 14185 25109 14197 25112
rect 14231 25109 14243 25143
rect 14185 25103 14243 25109
rect 15838 25100 15844 25152
rect 15896 25140 15902 25152
rect 22204 25149 22232 25248
rect 22925 25245 22937 25248
rect 22971 25245 22983 25279
rect 22925 25239 22983 25245
rect 24486 25236 24492 25288
rect 24544 25276 24550 25288
rect 24581 25279 24639 25285
rect 24581 25276 24593 25279
rect 24544 25248 24593 25276
rect 24544 25236 24550 25248
rect 24581 25245 24593 25248
rect 24627 25245 24639 25279
rect 24581 25239 24639 25245
rect 24857 25279 24915 25285
rect 24857 25245 24869 25279
rect 24903 25276 24915 25279
rect 25038 25276 25044 25288
rect 24903 25248 25044 25276
rect 24903 25245 24915 25248
rect 24857 25239 24915 25245
rect 25038 25236 25044 25248
rect 25096 25236 25102 25288
rect 45649 25279 45707 25285
rect 45649 25245 45661 25279
rect 45695 25276 45707 25279
rect 45738 25276 45744 25288
rect 45695 25248 45744 25276
rect 45695 25245 45707 25248
rect 45649 25239 45707 25245
rect 45738 25236 45744 25248
rect 45796 25236 45802 25288
rect 46290 25276 46296 25288
rect 46251 25248 46296 25276
rect 46290 25236 46296 25248
rect 46348 25236 46354 25288
rect 22646 25208 22652 25220
rect 22607 25180 22652 25208
rect 22646 25168 22652 25180
rect 22704 25168 22710 25220
rect 22830 25208 22836 25220
rect 22791 25180 22836 25208
rect 22830 25168 22836 25180
rect 22888 25168 22894 25220
rect 24765 25211 24823 25217
rect 24765 25208 24777 25211
rect 23124 25180 24777 25208
rect 15933 25143 15991 25149
rect 15933 25140 15945 25143
rect 15896 25112 15945 25140
rect 15896 25100 15902 25112
rect 15933 25109 15945 25112
rect 15979 25109 15991 25143
rect 15933 25103 15991 25109
rect 22189 25143 22247 25149
rect 22189 25109 22201 25143
rect 22235 25109 22247 25143
rect 22664 25140 22692 25168
rect 23124 25140 23152 25180
rect 24765 25177 24777 25180
rect 24811 25177 24823 25211
rect 24765 25171 24823 25177
rect 25593 25211 25651 25217
rect 25593 25177 25605 25211
rect 25639 25177 25651 25211
rect 25593 25171 25651 25177
rect 22664 25112 23152 25140
rect 22189 25103 22247 25109
rect 23750 25100 23756 25152
rect 23808 25140 23814 25152
rect 24397 25143 24455 25149
rect 24397 25140 24409 25143
rect 23808 25112 24409 25140
rect 23808 25100 23814 25112
rect 24397 25109 24409 25112
rect 24443 25109 24455 25143
rect 25608 25140 25636 25171
rect 26050 25168 26056 25220
rect 26108 25168 26114 25220
rect 46477 25211 46535 25217
rect 46477 25177 46489 25211
rect 46523 25208 46535 25211
rect 47670 25208 47676 25220
rect 46523 25180 47676 25208
rect 46523 25177 46535 25180
rect 46477 25171 46535 25177
rect 47670 25168 47676 25180
rect 47728 25168 47734 25220
rect 26418 25140 26424 25152
rect 25608 25112 26424 25140
rect 24397 25103 24455 25109
rect 26418 25100 26424 25112
rect 26476 25100 26482 25152
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 22373 24939 22431 24945
rect 22373 24905 22385 24939
rect 22419 24936 22431 24939
rect 22646 24936 22652 24948
rect 22419 24908 22652 24936
rect 22419 24905 22431 24908
rect 22373 24899 22431 24905
rect 22646 24896 22652 24908
rect 22704 24896 22710 24948
rect 25222 24936 25228 24948
rect 25183 24908 25228 24936
rect 25222 24896 25228 24908
rect 25280 24896 25286 24948
rect 46198 24896 46204 24948
rect 46256 24936 46262 24948
rect 46750 24936 46756 24948
rect 46256 24908 46756 24936
rect 46256 24896 46262 24908
rect 46750 24896 46756 24908
rect 46808 24896 46814 24948
rect 14090 24828 14096 24880
rect 14148 24828 14154 24880
rect 23750 24868 23756 24880
rect 23711 24840 23756 24868
rect 23750 24828 23756 24840
rect 23808 24828 23814 24880
rect 45554 24868 45560 24880
rect 45204 24840 45560 24868
rect 9861 24803 9919 24809
rect 9861 24769 9873 24803
rect 9907 24800 9919 24803
rect 11422 24800 11428 24812
rect 9907 24772 11428 24800
rect 9907 24769 9919 24772
rect 9861 24763 9919 24769
rect 11422 24760 11428 24772
rect 11480 24760 11486 24812
rect 17681 24803 17739 24809
rect 17681 24769 17693 24803
rect 17727 24769 17739 24803
rect 17681 24763 17739 24769
rect 17773 24803 17831 24809
rect 17773 24769 17785 24803
rect 17819 24800 17831 24803
rect 17954 24800 17960 24812
rect 17819 24772 17960 24800
rect 17819 24769 17831 24772
rect 17773 24763 17831 24769
rect 9950 24732 9956 24744
rect 9863 24704 9956 24732
rect 9950 24692 9956 24704
rect 10008 24732 10014 24744
rect 10962 24732 10968 24744
rect 10008 24704 10968 24732
rect 10008 24692 10014 24704
rect 10962 24692 10968 24704
rect 11020 24692 11026 24744
rect 13078 24732 13084 24744
rect 13039 24704 13084 24732
rect 13078 24692 13084 24704
rect 13136 24692 13142 24744
rect 13354 24732 13360 24744
rect 13315 24704 13360 24732
rect 13354 24692 13360 24704
rect 13412 24692 13418 24744
rect 17696 24732 17724 24763
rect 17954 24760 17960 24772
rect 18012 24760 18018 24812
rect 18874 24760 18880 24812
rect 18932 24800 18938 24812
rect 19153 24803 19211 24809
rect 19153 24800 19165 24803
rect 18932 24772 19165 24800
rect 18932 24760 18938 24772
rect 19153 24769 19165 24772
rect 19199 24769 19211 24803
rect 19978 24800 19984 24812
rect 19939 24772 19984 24800
rect 19153 24763 19211 24769
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 22186 24800 22192 24812
rect 22147 24772 22192 24800
rect 22186 24760 22192 24772
rect 22244 24760 22250 24812
rect 22462 24760 22468 24812
rect 22520 24800 22526 24812
rect 23474 24800 23480 24812
rect 22520 24772 22565 24800
rect 23435 24772 23480 24800
rect 22520 24760 22526 24772
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 24854 24760 24860 24812
rect 24912 24760 24918 24812
rect 45204 24800 45232 24840
rect 45554 24828 45560 24840
rect 45612 24828 45618 24880
rect 31726 24772 45232 24800
rect 17696 24704 18000 24732
rect 17972 24676 18000 24704
rect 24762 24692 24768 24744
rect 24820 24732 24826 24744
rect 31726 24732 31754 24772
rect 47486 24760 47492 24812
rect 47544 24800 47550 24812
rect 47581 24803 47639 24809
rect 47581 24800 47593 24803
rect 47544 24772 47593 24800
rect 47544 24760 47550 24772
rect 47581 24769 47593 24772
rect 47627 24769 47639 24803
rect 47581 24763 47639 24769
rect 47670 24760 47676 24812
rect 47728 24800 47734 24812
rect 47728 24772 47773 24800
rect 47728 24760 47734 24772
rect 24820 24704 31754 24732
rect 45189 24735 45247 24741
rect 24820 24692 24826 24704
rect 45189 24701 45201 24735
rect 45235 24701 45247 24735
rect 45370 24732 45376 24744
rect 45331 24704 45376 24732
rect 45189 24695 45247 24701
rect 9674 24624 9680 24676
rect 9732 24664 9738 24676
rect 10229 24667 10287 24673
rect 10229 24664 10241 24667
rect 9732 24636 10241 24664
rect 9732 24624 9738 24636
rect 10229 24633 10241 24636
rect 10275 24633 10287 24667
rect 15746 24664 15752 24676
rect 10229 24627 10287 24633
rect 14752 24636 15752 24664
rect 10962 24556 10968 24608
rect 11020 24596 11026 24608
rect 14752 24596 14780 24636
rect 15746 24624 15752 24636
rect 15804 24664 15810 24676
rect 16482 24664 16488 24676
rect 15804 24636 16488 24664
rect 15804 24624 15810 24636
rect 16482 24624 16488 24636
rect 16540 24624 16546 24676
rect 17954 24624 17960 24676
rect 18012 24624 18018 24676
rect 22830 24664 22836 24676
rect 19352 24636 22836 24664
rect 11020 24568 14780 24596
rect 14829 24599 14887 24605
rect 11020 24556 11026 24568
rect 14829 24565 14841 24599
rect 14875 24596 14887 24599
rect 15470 24596 15476 24608
rect 14875 24568 15476 24596
rect 14875 24565 14887 24568
rect 14829 24559 14887 24565
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 19150 24556 19156 24608
rect 19208 24596 19214 24608
rect 19352 24605 19380 24636
rect 22830 24624 22836 24636
rect 22888 24664 22894 24676
rect 23382 24664 23388 24676
rect 22888 24636 23388 24664
rect 22888 24624 22894 24636
rect 23382 24624 23388 24636
rect 23440 24624 23446 24676
rect 19337 24599 19395 24605
rect 19337 24596 19349 24599
rect 19208 24568 19349 24596
rect 19208 24556 19214 24568
rect 19337 24565 19349 24568
rect 19383 24565 19395 24599
rect 19337 24559 19395 24565
rect 20073 24599 20131 24605
rect 20073 24565 20085 24599
rect 20119 24596 20131 24599
rect 20346 24596 20352 24608
rect 20119 24568 20352 24596
rect 20119 24565 20131 24568
rect 20073 24559 20131 24565
rect 20346 24556 20352 24568
rect 20404 24556 20410 24608
rect 22002 24596 22008 24608
rect 21963 24568 22008 24596
rect 22002 24556 22008 24568
rect 22060 24556 22066 24608
rect 45204 24596 45232 24695
rect 45370 24692 45376 24704
rect 45428 24692 45434 24744
rect 46842 24732 46848 24744
rect 46803 24704 46848 24732
rect 46842 24692 46848 24704
rect 46900 24692 46906 24744
rect 46842 24596 46848 24608
rect 45204 24568 46848 24596
rect 46842 24556 46848 24568
rect 46900 24556 46906 24608
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 10410 24352 10416 24404
rect 10468 24392 10474 24404
rect 10505 24395 10563 24401
rect 10505 24392 10517 24395
rect 10468 24364 10517 24392
rect 10468 24352 10474 24364
rect 10505 24361 10517 24364
rect 10551 24361 10563 24395
rect 10505 24355 10563 24361
rect 13173 24395 13231 24401
rect 13173 24361 13185 24395
rect 13219 24392 13231 24395
rect 13354 24392 13360 24404
rect 13219 24364 13360 24392
rect 13219 24361 13231 24364
rect 13173 24355 13231 24361
rect 13354 24352 13360 24364
rect 13412 24352 13418 24404
rect 21361 24395 21419 24401
rect 21361 24361 21373 24395
rect 21407 24392 21419 24395
rect 21910 24392 21916 24404
rect 21407 24364 21916 24392
rect 21407 24361 21419 24364
rect 21361 24355 21419 24361
rect 21910 24352 21916 24364
rect 21968 24352 21974 24404
rect 24946 24352 24952 24404
rect 25004 24392 25010 24404
rect 25130 24392 25136 24404
rect 25004 24364 25136 24392
rect 25004 24352 25010 24364
rect 25130 24352 25136 24364
rect 25188 24352 25194 24404
rect 12986 24324 12992 24336
rect 12084 24296 12992 24324
rect 10410 24188 10416 24200
rect 10371 24160 10416 24188
rect 10410 24148 10416 24160
rect 10468 24148 10474 24200
rect 12084 24197 12112 24296
rect 12986 24284 12992 24296
rect 13044 24284 13050 24336
rect 13078 24284 13084 24336
rect 13136 24324 13142 24336
rect 14093 24327 14151 24333
rect 14093 24324 14105 24327
rect 13136 24296 14105 24324
rect 13136 24284 13142 24296
rect 14093 24293 14105 24296
rect 14139 24293 14151 24327
rect 14093 24287 14151 24293
rect 20990 24284 20996 24336
rect 21048 24324 21054 24336
rect 40770 24324 40776 24336
rect 21048 24296 40776 24324
rect 21048 24284 21054 24296
rect 40770 24284 40776 24296
rect 40828 24284 40834 24336
rect 12802 24256 12808 24268
rect 12763 24228 12808 24256
rect 12802 24216 12808 24228
rect 12860 24216 12866 24268
rect 15470 24256 15476 24268
rect 12912 24228 15476 24256
rect 12912 24197 12940 24228
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 16574 24216 16580 24268
rect 16632 24256 16638 24268
rect 16632 24228 16988 24256
rect 16632 24216 16638 24228
rect 12069 24191 12127 24197
rect 12069 24157 12081 24191
rect 12115 24157 12127 24191
rect 12069 24151 12127 24157
rect 12897 24191 12955 24197
rect 12897 24157 12909 24191
rect 12943 24157 12955 24191
rect 12897 24151 12955 24157
rect 12802 24080 12808 24132
rect 12860 24120 12866 24132
rect 12912 24120 12940 24151
rect 12986 24148 12992 24200
rect 13044 24188 13050 24200
rect 13044 24160 13676 24188
rect 13044 24148 13050 24160
rect 12860 24092 12940 24120
rect 12860 24080 12866 24092
rect 12161 24055 12219 24061
rect 12161 24021 12173 24055
rect 12207 24052 12219 24055
rect 12986 24052 12992 24064
rect 12207 24024 12992 24052
rect 12207 24021 12219 24024
rect 12161 24015 12219 24021
rect 12986 24012 12992 24024
rect 13044 24012 13050 24064
rect 13648 24052 13676 24160
rect 13998 24148 14004 24200
rect 14056 24188 14062 24200
rect 14093 24191 14151 24197
rect 14093 24188 14105 24191
rect 14056 24160 14105 24188
rect 14056 24148 14062 24160
rect 14093 24157 14105 24160
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 15013 24191 15071 24197
rect 15013 24157 15025 24191
rect 15059 24188 15071 24191
rect 15746 24188 15752 24200
rect 15059 24160 15752 24188
rect 15059 24157 15071 24160
rect 15013 24151 15071 24157
rect 15746 24148 15752 24160
rect 15804 24148 15810 24200
rect 16022 24188 16028 24200
rect 15983 24160 16028 24188
rect 16022 24148 16028 24160
rect 16080 24148 16086 24200
rect 16390 24188 16396 24200
rect 16351 24160 16396 24188
rect 16390 24148 16396 24160
rect 16448 24148 16454 24200
rect 16482 24148 16488 24200
rect 16540 24188 16546 24200
rect 16960 24197 16988 24228
rect 19242 24216 19248 24268
rect 19300 24256 19306 24268
rect 19613 24259 19671 24265
rect 19613 24256 19625 24259
rect 19300 24228 19625 24256
rect 19300 24216 19306 24228
rect 19613 24225 19625 24228
rect 19659 24225 19671 24259
rect 19613 24219 19671 24225
rect 19889 24259 19947 24265
rect 19889 24225 19901 24259
rect 19935 24256 19947 24259
rect 22002 24256 22008 24268
rect 19935 24228 22008 24256
rect 19935 24225 19947 24228
rect 19889 24219 19947 24225
rect 22002 24216 22008 24228
rect 22060 24216 22066 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 16945 24191 17003 24197
rect 16540 24160 16585 24188
rect 16540 24148 16546 24160
rect 16945 24157 16957 24191
rect 16991 24157 17003 24191
rect 17954 24188 17960 24200
rect 17915 24160 17960 24188
rect 16945 24151 17003 24157
rect 17954 24148 17960 24160
rect 18012 24148 18018 24200
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 22066 24160 24409 24188
rect 13722 24080 13728 24132
rect 13780 24120 13786 24132
rect 13780 24092 18184 24120
rect 13780 24080 13786 24092
rect 14734 24052 14740 24064
rect 13648 24024 14740 24052
rect 14734 24012 14740 24024
rect 14792 24052 14798 24064
rect 15197 24055 15255 24061
rect 15197 24052 15209 24055
rect 14792 24024 15209 24052
rect 14792 24012 14798 24024
rect 15197 24021 15209 24024
rect 15243 24021 15255 24055
rect 16298 24052 16304 24064
rect 16259 24024 16304 24052
rect 15197 24015 15255 24021
rect 16298 24012 16304 24024
rect 16356 24012 16362 24064
rect 16666 24012 16672 24064
rect 16724 24052 16730 24064
rect 17129 24055 17187 24061
rect 17129 24052 17141 24055
rect 16724 24024 17141 24052
rect 16724 24012 16730 24024
rect 17129 24021 17141 24024
rect 17175 24021 17187 24055
rect 18046 24052 18052 24064
rect 18007 24024 18052 24052
rect 17129 24015 17187 24021
rect 18046 24012 18052 24024
rect 18104 24012 18110 24064
rect 18156 24052 18184 24092
rect 20346 24080 20352 24132
rect 20404 24080 20410 24132
rect 22066 24052 22094 24160
rect 24397 24157 24409 24160
rect 24443 24188 24455 24191
rect 24762 24188 24768 24200
rect 24443 24160 24768 24188
rect 24443 24157 24455 24160
rect 24397 24151 24455 24157
rect 24762 24148 24768 24160
rect 24820 24148 24826 24200
rect 24854 24148 24860 24200
rect 24912 24188 24918 24200
rect 26513 24191 26571 24197
rect 26513 24188 26525 24191
rect 24912 24160 26525 24188
rect 24912 24148 24918 24160
rect 26513 24157 26525 24160
rect 26559 24157 26571 24191
rect 26513 24151 26571 24157
rect 27249 24191 27307 24197
rect 27249 24157 27261 24191
rect 27295 24157 27307 24191
rect 27249 24151 27307 24157
rect 25498 24120 25504 24132
rect 24596 24092 25504 24120
rect 18156 24024 22094 24052
rect 22278 24012 22284 24064
rect 22336 24052 22342 24064
rect 23658 24052 23664 24064
rect 22336 24024 23664 24052
rect 22336 24012 22342 24024
rect 23658 24012 23664 24024
rect 23716 24052 23722 24064
rect 24596 24061 24624 24092
rect 25498 24080 25504 24092
rect 25556 24120 25562 24132
rect 27264 24120 27292 24151
rect 28810 24148 28816 24200
rect 28868 24188 28874 24200
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 28868 24160 29561 24188
rect 28868 24148 28874 24160
rect 29549 24157 29561 24160
rect 29595 24157 29607 24191
rect 29549 24151 29607 24157
rect 45833 24191 45891 24197
rect 45833 24157 45845 24191
rect 45879 24188 45891 24191
rect 46293 24191 46351 24197
rect 46293 24188 46305 24191
rect 45879 24160 46305 24188
rect 45879 24157 45891 24160
rect 45833 24151 45891 24157
rect 46293 24157 46305 24160
rect 46339 24157 46351 24191
rect 46293 24151 46351 24157
rect 29730 24120 29736 24132
rect 25556 24092 27292 24120
rect 29691 24092 29736 24120
rect 25556 24080 25562 24092
rect 29730 24080 29736 24092
rect 29788 24080 29794 24132
rect 31389 24123 31447 24129
rect 31389 24089 31401 24123
rect 31435 24120 31447 24123
rect 40034 24120 40040 24132
rect 31435 24092 40040 24120
rect 31435 24089 31447 24092
rect 31389 24083 31447 24089
rect 40034 24080 40040 24092
rect 40092 24080 40098 24132
rect 46477 24123 46535 24129
rect 46477 24089 46489 24123
rect 46523 24120 46535 24123
rect 47670 24120 47676 24132
rect 46523 24092 47676 24120
rect 46523 24089 46535 24092
rect 46477 24083 46535 24089
rect 47670 24080 47676 24092
rect 47728 24080 47734 24132
rect 24581 24055 24639 24061
rect 24581 24052 24593 24055
rect 23716 24024 24593 24052
rect 23716 24012 23722 24024
rect 24581 24021 24593 24024
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 26697 24055 26755 24061
rect 26697 24021 26709 24055
rect 26743 24052 26755 24055
rect 26970 24052 26976 24064
rect 26743 24024 26976 24052
rect 26743 24021 26755 24024
rect 26697 24015 26755 24021
rect 26970 24012 26976 24024
rect 27028 24012 27034 24064
rect 27338 24052 27344 24064
rect 27299 24024 27344 24052
rect 27338 24012 27344 24024
rect 27396 24012 27402 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 13722 23848 13728 23860
rect 12084 23820 13728 23848
rect 11882 23780 11888 23792
rect 7484 23752 11888 23780
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 7484 23721 7512 23752
rect 11882 23740 11888 23752
rect 11940 23740 11946 23792
rect 7469 23715 7527 23721
rect 7469 23681 7481 23715
rect 7515 23681 7527 23715
rect 10318 23712 10324 23724
rect 10279 23684 10324 23712
rect 7469 23675 7527 23681
rect 10318 23672 10324 23684
rect 10376 23672 10382 23724
rect 12084 23721 12112 23820
rect 13722 23808 13728 23820
rect 13780 23808 13786 23860
rect 15930 23848 15936 23860
rect 15891 23820 15936 23848
rect 15930 23808 15936 23820
rect 15988 23808 15994 23860
rect 16117 23851 16175 23857
rect 16117 23817 16129 23851
rect 16163 23848 16175 23851
rect 16390 23848 16396 23860
rect 16163 23820 16396 23848
rect 16163 23817 16175 23820
rect 16117 23811 16175 23817
rect 16390 23808 16396 23820
rect 16448 23808 16454 23860
rect 17954 23808 17960 23860
rect 18012 23848 18018 23860
rect 22278 23848 22284 23860
rect 18012 23820 22284 23848
rect 18012 23808 18018 23820
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 22388 23820 40724 23848
rect 12986 23780 12992 23792
rect 12947 23752 12992 23780
rect 12986 23740 12992 23752
rect 13044 23740 13050 23792
rect 15470 23740 15476 23792
rect 15528 23780 15534 23792
rect 15841 23783 15899 23789
rect 15841 23780 15853 23783
rect 15528 23752 15853 23780
rect 15528 23740 15534 23752
rect 15841 23749 15853 23752
rect 15887 23749 15899 23783
rect 15841 23743 15899 23749
rect 16298 23740 16304 23792
rect 16356 23780 16362 23792
rect 16945 23783 17003 23789
rect 16945 23780 16957 23783
rect 16356 23752 16957 23780
rect 16356 23740 16362 23752
rect 16945 23749 16957 23752
rect 16991 23749 17003 23783
rect 16945 23743 17003 23749
rect 20993 23783 21051 23789
rect 20993 23749 21005 23783
rect 21039 23780 21051 23783
rect 22388 23780 22416 23820
rect 27246 23780 27252 23792
rect 21039 23752 22416 23780
rect 22940 23752 27252 23780
rect 21039 23749 21051 23752
rect 20993 23743 21051 23749
rect 12069 23715 12127 23721
rect 12069 23681 12081 23715
rect 12115 23681 12127 23715
rect 12802 23712 12808 23724
rect 12763 23684 12808 23712
rect 12069 23675 12127 23681
rect 7650 23644 7656 23656
rect 7611 23616 7656 23644
rect 7650 23604 7656 23616
rect 7708 23604 7714 23656
rect 7926 23644 7932 23656
rect 7887 23616 7932 23644
rect 7926 23604 7932 23616
rect 7984 23604 7990 23656
rect 11882 23604 11888 23656
rect 11940 23644 11946 23656
rect 12084 23644 12112 23675
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 15749 23715 15807 23721
rect 15749 23681 15761 23715
rect 15795 23681 15807 23715
rect 16666 23712 16672 23724
rect 16627 23684 16672 23712
rect 15749 23675 15807 23681
rect 13814 23644 13820 23656
rect 11940 23616 12112 23644
rect 13775 23616 13820 23644
rect 11940 23604 11946 23616
rect 13814 23604 13820 23616
rect 13872 23604 13878 23656
rect 15764 23644 15792 23675
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 18046 23672 18052 23724
rect 18104 23672 18110 23724
rect 22094 23712 22100 23724
rect 22055 23684 22100 23712
rect 22094 23672 22100 23684
rect 22152 23672 22158 23724
rect 16114 23644 16120 23656
rect 15764 23616 16120 23644
rect 16114 23604 16120 23616
rect 16172 23604 16178 23656
rect 19153 23647 19211 23653
rect 19153 23644 19165 23647
rect 18432 23616 19165 23644
rect 15286 23576 15292 23588
rect 6886 23548 15292 23576
rect 1949 23511 2007 23517
rect 1949 23477 1961 23511
rect 1995 23508 2007 23511
rect 6886 23508 6914 23548
rect 15286 23536 15292 23548
rect 15344 23536 15350 23588
rect 15565 23579 15623 23585
rect 15565 23545 15577 23579
rect 15611 23576 15623 23579
rect 16666 23576 16672 23588
rect 15611 23548 16672 23576
rect 15611 23545 15623 23548
rect 15565 23539 15623 23545
rect 16666 23536 16672 23548
rect 16724 23536 16730 23588
rect 10318 23508 10324 23520
rect 1995 23480 6914 23508
rect 10279 23480 10324 23508
rect 1995 23477 2007 23480
rect 1949 23471 2007 23477
rect 10318 23468 10324 23480
rect 10376 23468 10382 23520
rect 12250 23508 12256 23520
rect 12211 23480 12256 23508
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 16684 23508 16712 23536
rect 18432 23517 18460 23616
rect 19153 23613 19165 23616
rect 19199 23613 19211 23647
rect 19334 23644 19340 23656
rect 19295 23616 19340 23644
rect 19153 23607 19211 23613
rect 19334 23604 19340 23616
rect 19392 23604 19398 23656
rect 20806 23604 20812 23656
rect 20864 23644 20870 23656
rect 22189 23647 22247 23653
rect 22189 23644 22201 23647
rect 20864 23616 22201 23644
rect 20864 23604 20870 23616
rect 22189 23613 22201 23616
rect 22235 23644 22247 23647
rect 22940 23644 22968 23752
rect 23109 23715 23167 23721
rect 23109 23681 23121 23715
rect 23155 23681 23167 23715
rect 23658 23712 23664 23724
rect 23619 23684 23664 23712
rect 23109 23675 23167 23681
rect 22235 23616 22968 23644
rect 22235 23613 22247 23616
rect 22189 23607 22247 23613
rect 23014 23604 23020 23656
rect 23072 23644 23078 23656
rect 23124 23644 23152 23675
rect 23658 23672 23664 23684
rect 23716 23672 23722 23724
rect 24673 23715 24731 23721
rect 24673 23681 24685 23715
rect 24719 23712 24731 23715
rect 24854 23712 24860 23724
rect 24719 23684 24860 23712
rect 24719 23681 24731 23684
rect 24673 23675 24731 23681
rect 24688 23644 24716 23675
rect 24854 23672 24860 23684
rect 24912 23672 24918 23724
rect 25501 23715 25559 23721
rect 25501 23681 25513 23715
rect 25547 23681 25559 23715
rect 25682 23712 25688 23724
rect 25643 23684 25688 23712
rect 25501 23675 25559 23681
rect 23072 23616 24716 23644
rect 23072 23604 23078 23616
rect 25516 23576 25544 23675
rect 25682 23672 25688 23684
rect 25740 23672 25746 23724
rect 26142 23712 26148 23724
rect 26103 23684 26148 23712
rect 26142 23672 26148 23684
rect 26200 23672 26206 23724
rect 26234 23672 26240 23724
rect 26292 23712 26298 23724
rect 26436 23721 26464 23752
rect 27246 23740 27252 23752
rect 27304 23740 27310 23792
rect 27338 23740 27344 23792
rect 27396 23780 27402 23792
rect 31573 23783 31631 23789
rect 27396 23752 27738 23780
rect 27396 23740 27402 23752
rect 31573 23749 31585 23783
rect 31619 23780 31631 23783
rect 37274 23780 37280 23792
rect 31619 23752 37280 23780
rect 31619 23749 31631 23752
rect 31573 23743 31631 23749
rect 37274 23740 37280 23752
rect 37332 23740 37338 23792
rect 40696 23780 40724 23820
rect 40770 23808 40776 23860
rect 40828 23848 40834 23860
rect 40828 23820 40873 23848
rect 40828 23808 40834 23820
rect 45370 23808 45376 23860
rect 45428 23848 45434 23860
rect 46937 23851 46995 23857
rect 46937 23848 46949 23851
rect 45428 23820 46949 23848
rect 45428 23808 45434 23820
rect 46937 23817 46949 23820
rect 46983 23817 46995 23851
rect 47670 23848 47676 23860
rect 47631 23820 47676 23848
rect 46937 23811 46995 23817
rect 47670 23808 47676 23820
rect 47728 23808 47734 23860
rect 46566 23780 46572 23792
rect 40696 23752 46572 23780
rect 46566 23740 46572 23752
rect 46624 23740 46630 23792
rect 26329 23715 26387 23721
rect 26329 23712 26341 23715
rect 26292 23684 26341 23712
rect 26292 23672 26298 23684
rect 26329 23681 26341 23684
rect 26375 23681 26387 23715
rect 26329 23675 26387 23681
rect 26421 23715 26479 23721
rect 26421 23681 26433 23715
rect 26467 23681 26479 23715
rect 26970 23712 26976 23724
rect 26931 23684 26976 23712
rect 26421 23675 26479 23681
rect 26970 23672 26976 23684
rect 27028 23672 27034 23724
rect 40770 23672 40776 23724
rect 40828 23712 40834 23724
rect 41141 23715 41199 23721
rect 41141 23712 41153 23715
rect 40828 23684 41153 23712
rect 40828 23672 40834 23684
rect 41141 23681 41153 23684
rect 41187 23712 41199 23715
rect 41187 23684 41368 23712
rect 41187 23681 41199 23684
rect 41141 23675 41199 23681
rect 25593 23647 25651 23653
rect 25593 23613 25605 23647
rect 25639 23644 25651 23647
rect 27249 23647 27307 23653
rect 27249 23644 27261 23647
rect 25639 23616 27261 23644
rect 25639 23613 25651 23616
rect 25593 23607 25651 23613
rect 27249 23613 27261 23616
rect 27295 23613 27307 23647
rect 27249 23607 27307 23613
rect 28721 23647 28779 23653
rect 28721 23613 28733 23647
rect 28767 23644 28779 23647
rect 28810 23644 28816 23656
rect 28767 23616 28816 23644
rect 28767 23613 28779 23616
rect 28721 23607 28779 23613
rect 28810 23604 28816 23616
rect 28868 23604 28874 23656
rect 28994 23604 29000 23656
rect 29052 23644 29058 23656
rect 29733 23647 29791 23653
rect 29733 23644 29745 23647
rect 29052 23616 29745 23644
rect 29052 23604 29058 23616
rect 29733 23613 29745 23616
rect 29779 23613 29791 23647
rect 29914 23644 29920 23656
rect 29875 23616 29920 23644
rect 29733 23607 29791 23613
rect 29914 23604 29920 23616
rect 29972 23604 29978 23656
rect 26145 23579 26203 23585
rect 26145 23576 26157 23579
rect 25516 23548 26157 23576
rect 26145 23545 26157 23548
rect 26191 23545 26203 23579
rect 41340 23576 41368 23684
rect 41414 23672 41420 23724
rect 41472 23712 41478 23724
rect 42429 23715 42487 23721
rect 42429 23712 42441 23715
rect 41472 23684 42441 23712
rect 41472 23672 41478 23684
rect 42429 23681 42441 23684
rect 42475 23681 42487 23715
rect 42429 23675 42487 23681
rect 46750 23672 46756 23724
rect 46808 23712 46814 23724
rect 46845 23715 46903 23721
rect 46845 23712 46857 23715
rect 46808 23684 46857 23712
rect 46808 23672 46814 23684
rect 46845 23681 46857 23684
rect 46891 23681 46903 23715
rect 46845 23675 46903 23681
rect 47118 23672 47124 23724
rect 47176 23712 47182 23724
rect 47578 23712 47584 23724
rect 47176 23684 47584 23712
rect 47176 23672 47182 23684
rect 47578 23672 47584 23684
rect 47636 23672 47642 23724
rect 42705 23647 42763 23653
rect 42705 23613 42717 23647
rect 42751 23644 42763 23647
rect 47136 23644 47164 23672
rect 42751 23616 47164 23644
rect 42751 23613 42763 23616
rect 42705 23607 42763 23613
rect 45738 23576 45744 23588
rect 41340 23548 45744 23576
rect 26145 23539 26203 23545
rect 45738 23536 45744 23548
rect 45796 23536 45802 23588
rect 18417 23511 18475 23517
rect 18417 23508 18429 23511
rect 16684 23480 18429 23508
rect 18417 23477 18429 23480
rect 18463 23477 18475 23511
rect 18417 23471 18475 23477
rect 20806 23468 20812 23520
rect 20864 23508 20870 23520
rect 21174 23508 21180 23520
rect 20864 23480 21180 23508
rect 20864 23468 20870 23480
rect 21174 23468 21180 23480
rect 21232 23468 21238 23520
rect 22278 23468 22284 23520
rect 22336 23508 22342 23520
rect 22465 23511 22523 23517
rect 22465 23508 22477 23511
rect 22336 23480 22477 23508
rect 22336 23468 22342 23480
rect 22465 23477 22477 23480
rect 22511 23477 22523 23511
rect 22922 23508 22928 23520
rect 22883 23480 22928 23508
rect 22465 23471 22523 23477
rect 22922 23468 22928 23480
rect 22980 23468 22986 23520
rect 23566 23468 23572 23520
rect 23624 23508 23630 23520
rect 23753 23511 23811 23517
rect 23753 23508 23765 23511
rect 23624 23480 23765 23508
rect 23624 23468 23630 23480
rect 23753 23477 23765 23480
rect 23799 23477 23811 23511
rect 24486 23508 24492 23520
rect 24447 23480 24492 23508
rect 23753 23471 23811 23477
rect 24486 23468 24492 23480
rect 24544 23468 24550 23520
rect 41322 23468 41328 23520
rect 41380 23508 41386 23520
rect 41417 23511 41475 23517
rect 41417 23508 41429 23511
rect 41380 23480 41429 23508
rect 41380 23468 41386 23480
rect 41417 23477 41429 23480
rect 41463 23477 41475 23511
rect 41417 23471 41475 23477
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 7650 23264 7656 23316
rect 7708 23304 7714 23316
rect 7745 23307 7803 23313
rect 7745 23304 7757 23307
rect 7708 23276 7757 23304
rect 7708 23264 7714 23276
rect 7745 23273 7757 23276
rect 7791 23273 7803 23307
rect 7745 23267 7803 23273
rect 16022 23264 16028 23316
rect 16080 23304 16086 23316
rect 16485 23307 16543 23313
rect 16485 23304 16497 23307
rect 16080 23276 16497 23304
rect 16080 23264 16086 23276
rect 16485 23273 16497 23276
rect 16531 23273 16543 23307
rect 16485 23267 16543 23273
rect 16574 23264 16580 23316
rect 16632 23304 16638 23316
rect 22922 23304 22928 23316
rect 16632 23276 19334 23304
rect 16632 23264 16638 23276
rect 15470 23236 15476 23248
rect 15431 23208 15476 23236
rect 15470 23196 15476 23208
rect 15528 23196 15534 23248
rect 15746 23196 15752 23248
rect 15804 23236 15810 23248
rect 15804 23208 17540 23236
rect 15804 23196 15810 23208
rect 2130 23128 2136 23180
rect 2188 23168 2194 23180
rect 16574 23168 16580 23180
rect 2188 23140 16580 23168
rect 2188 23128 2194 23140
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 7650 23100 7656 23112
rect 7611 23072 7656 23100
rect 7650 23060 7656 23072
rect 7708 23060 7714 23112
rect 8941 23103 8999 23109
rect 8941 23069 8953 23103
rect 8987 23100 8999 23103
rect 9674 23100 9680 23112
rect 8987 23072 9536 23100
rect 9635 23072 9680 23100
rect 8987 23069 8999 23072
rect 8941 23063 8999 23069
rect 8938 22924 8944 22976
rect 8996 22964 9002 22976
rect 9033 22967 9091 22973
rect 9033 22964 9045 22967
rect 8996 22936 9045 22964
rect 8996 22924 9002 22936
rect 9033 22933 9045 22936
rect 9079 22933 9091 22967
rect 9508 22964 9536 23072
rect 9674 23060 9680 23072
rect 9732 23060 9738 23112
rect 9861 23103 9919 23109
rect 9861 23069 9873 23103
rect 9907 23100 9919 23103
rect 9950 23100 9956 23112
rect 9907 23072 9956 23100
rect 9907 23069 9919 23072
rect 9861 23063 9919 23069
rect 9950 23060 9956 23072
rect 10008 23060 10014 23112
rect 10318 23100 10324 23112
rect 10279 23072 10324 23100
rect 10318 23060 10324 23072
rect 10376 23060 10382 23112
rect 11974 23060 11980 23112
rect 12032 23100 12038 23112
rect 12529 23103 12587 23109
rect 12529 23100 12541 23103
rect 12032 23072 12541 23100
rect 12032 23060 12038 23072
rect 12529 23069 12541 23072
rect 12575 23069 12587 23103
rect 13357 23103 13415 23109
rect 13357 23100 13369 23103
rect 12529 23063 12587 23069
rect 13280 23072 13369 23100
rect 9769 23035 9827 23041
rect 9769 23001 9781 23035
rect 9815 23032 9827 23035
rect 10597 23035 10655 23041
rect 10597 23032 10609 23035
rect 9815 23004 10609 23032
rect 9815 23001 9827 23004
rect 9769 22995 9827 23001
rect 10597 23001 10609 23004
rect 10643 23001 10655 23035
rect 12621 23035 12679 23041
rect 12621 23032 12633 23035
rect 11822 23004 12633 23032
rect 10597 22995 10655 23001
rect 12621 23001 12633 23004
rect 12667 23001 12679 23035
rect 12621 22995 12679 23001
rect 10226 22964 10232 22976
rect 9508 22936 10232 22964
rect 9033 22927 9091 22933
rect 10226 22924 10232 22936
rect 10284 22924 10290 22976
rect 11514 22924 11520 22976
rect 11572 22964 11578 22976
rect 12069 22967 12127 22973
rect 12069 22964 12081 22967
rect 11572 22936 12081 22964
rect 11572 22924 11578 22936
rect 12069 22933 12081 22936
rect 12115 22933 12127 22967
rect 12069 22927 12127 22933
rect 12250 22924 12256 22976
rect 12308 22964 12314 22976
rect 13280 22964 13308 23072
rect 13357 23069 13369 23072
rect 13403 23100 13415 23103
rect 13906 23100 13912 23112
rect 13403 23072 13912 23100
rect 13403 23069 13415 23072
rect 13357 23063 13415 23069
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 13998 23060 14004 23112
rect 14056 23100 14062 23112
rect 14461 23103 14519 23109
rect 14461 23100 14473 23103
rect 14056 23072 14473 23100
rect 14056 23060 14062 23072
rect 14461 23069 14473 23072
rect 14507 23069 14519 23103
rect 15838 23100 15844 23112
rect 15799 23072 15844 23100
rect 14461 23063 14519 23069
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 16666 23100 16672 23112
rect 16627 23072 16672 23100
rect 16666 23060 16672 23072
rect 16724 23060 16730 23112
rect 16945 23103 17003 23109
rect 16945 23100 16957 23103
rect 16776 23072 16957 23100
rect 15657 23035 15715 23041
rect 15657 23001 15669 23035
rect 15703 23032 15715 23035
rect 16574 23032 16580 23044
rect 15703 23004 16580 23032
rect 15703 23001 15715 23004
rect 15657 22995 15715 23001
rect 16574 22992 16580 23004
rect 16632 22992 16638 23044
rect 13446 22964 13452 22976
rect 12308 22936 13308 22964
rect 13407 22936 13452 22964
rect 12308 22924 12314 22936
rect 13446 22924 13452 22936
rect 13504 22924 13510 22976
rect 14366 22924 14372 22976
rect 14424 22964 14430 22976
rect 14645 22967 14703 22973
rect 14645 22964 14657 22967
rect 14424 22936 14657 22964
rect 14424 22924 14430 22936
rect 14645 22933 14657 22936
rect 14691 22933 14703 22967
rect 14645 22927 14703 22933
rect 15749 22967 15807 22973
rect 15749 22933 15761 22967
rect 15795 22964 15807 22967
rect 15838 22964 15844 22976
rect 15795 22936 15844 22964
rect 15795 22933 15807 22936
rect 15749 22927 15807 22933
rect 15838 22924 15844 22936
rect 15896 22924 15902 22976
rect 16022 22964 16028 22976
rect 15983 22936 16028 22964
rect 16022 22924 16028 22936
rect 16080 22964 16086 22976
rect 16776 22964 16804 23072
rect 16945 23069 16957 23072
rect 16991 23069 17003 23103
rect 17512 23100 17540 23208
rect 19306 23168 19334 23276
rect 22020 23276 22928 23304
rect 21358 23168 21364 23180
rect 19306 23140 21364 23168
rect 21358 23128 21364 23140
rect 21416 23128 21422 23180
rect 22020 23177 22048 23276
rect 22922 23264 22928 23276
rect 22980 23264 22986 23316
rect 28077 23307 28135 23313
rect 28077 23273 28089 23307
rect 28123 23273 28135 23307
rect 28077 23267 28135 23273
rect 28905 23307 28963 23313
rect 28905 23273 28917 23307
rect 28951 23304 28963 23307
rect 29730 23304 29736 23316
rect 28951 23276 29736 23304
rect 28951 23273 28963 23276
rect 28905 23267 28963 23273
rect 28092 23236 28120 23267
rect 29730 23264 29736 23276
rect 29788 23264 29794 23316
rect 38286 23236 38292 23248
rect 27172 23208 28120 23236
rect 28966 23208 38292 23236
rect 22005 23171 22063 23177
rect 22005 23137 22017 23171
rect 22051 23137 22063 23171
rect 22278 23168 22284 23180
rect 22239 23140 22284 23168
rect 22005 23131 22063 23137
rect 22278 23128 22284 23140
rect 22336 23128 22342 23180
rect 24486 23128 24492 23180
rect 24544 23168 24550 23180
rect 24581 23171 24639 23177
rect 24581 23168 24593 23171
rect 24544 23140 24593 23168
rect 24544 23128 24550 23140
rect 24581 23137 24593 23140
rect 24627 23137 24639 23171
rect 24581 23131 24639 23137
rect 26234 23128 26240 23180
rect 26292 23168 26298 23180
rect 27172 23168 27200 23208
rect 26292 23140 27200 23168
rect 26292 23128 26298 23140
rect 18049 23103 18107 23109
rect 18049 23100 18061 23103
rect 17512 23072 18061 23100
rect 16945 23063 17003 23069
rect 18049 23069 18061 23072
rect 18095 23100 18107 23103
rect 19337 23103 19395 23109
rect 19337 23100 19349 23103
rect 18095 23072 19349 23100
rect 18095 23069 18107 23072
rect 18049 23063 18107 23069
rect 19337 23069 19349 23072
rect 19383 23100 19395 23103
rect 20530 23100 20536 23112
rect 19383 23072 20536 23100
rect 19383 23069 19395 23072
rect 19337 23063 19395 23069
rect 20530 23060 20536 23072
rect 20588 23060 20594 23112
rect 20714 23100 20720 23112
rect 20675 23072 20720 23100
rect 20714 23060 20720 23072
rect 20772 23060 20778 23112
rect 26142 23060 26148 23112
rect 26200 23100 26206 23112
rect 27172 23100 27200 23140
rect 27338 23128 27344 23180
rect 27396 23168 27402 23180
rect 28966 23168 28994 23208
rect 38286 23196 38292 23208
rect 38344 23196 38350 23248
rect 47302 23168 47308 23180
rect 27396 23140 28994 23168
rect 47263 23140 47308 23168
rect 27396 23128 27402 23140
rect 47302 23128 47308 23140
rect 47360 23128 47366 23180
rect 27249 23103 27307 23109
rect 27249 23100 27261 23103
rect 26200 23072 27108 23100
rect 27172 23072 27261 23100
rect 26200 23060 26206 23072
rect 18598 23032 18604 23044
rect 18559 23004 18604 23032
rect 18598 22992 18604 23004
rect 18656 22992 18662 23044
rect 18966 22992 18972 23044
rect 19024 23032 19030 23044
rect 19426 23032 19432 23044
rect 19024 23004 19432 23032
rect 19024 22992 19030 23004
rect 19426 22992 19432 23004
rect 19484 23032 19490 23044
rect 19705 23035 19763 23041
rect 19705 23032 19717 23035
rect 19484 23004 19717 23032
rect 19484 22992 19490 23004
rect 19705 23001 19717 23004
rect 19751 23001 19763 23035
rect 19705 22995 19763 23001
rect 22186 22992 22192 23044
rect 22244 23032 22250 23044
rect 23566 23032 23572 23044
rect 22244 23004 22692 23032
rect 23506 23004 23572 23032
rect 22244 22992 22250 23004
rect 16080 22936 16804 22964
rect 16080 22924 16086 22936
rect 16850 22924 16856 22976
rect 16908 22964 16914 22976
rect 22664 22964 22692 23004
rect 23566 22992 23572 23004
rect 23624 22992 23630 23044
rect 24854 23032 24860 23044
rect 24815 23004 24860 23032
rect 24854 22992 24860 23004
rect 24912 22992 24918 23044
rect 25590 22992 25596 23044
rect 25648 22992 25654 23044
rect 26234 23032 26240 23044
rect 26160 23004 26240 23032
rect 23753 22967 23811 22973
rect 23753 22964 23765 22967
rect 16908 22936 16953 22964
rect 22664 22936 23765 22964
rect 16908 22924 16914 22936
rect 23753 22933 23765 22936
rect 23799 22964 23811 22967
rect 26160 22964 26188 23004
rect 26234 22992 26240 23004
rect 26292 22992 26298 23044
rect 26881 23035 26939 23041
rect 26881 23001 26893 23035
rect 26927 23032 26939 23035
rect 26970 23032 26976 23044
rect 26927 23004 26976 23032
rect 26927 23001 26939 23004
rect 26881 22995 26939 23001
rect 26970 22992 26976 23004
rect 27028 22992 27034 23044
rect 27080 23032 27108 23072
rect 27249 23069 27261 23072
rect 27295 23069 27307 23103
rect 27249 23063 27307 23069
rect 28626 23060 28632 23112
rect 28684 23100 28690 23112
rect 28813 23103 28871 23109
rect 28813 23102 28825 23103
rect 28736 23100 28825 23102
rect 28684 23074 28825 23100
rect 28684 23072 28764 23074
rect 28684 23060 28690 23072
rect 28813 23069 28825 23074
rect 28859 23069 28871 23103
rect 28813 23063 28871 23069
rect 28902 23060 28908 23112
rect 28960 23100 28966 23112
rect 41322 23100 41328 23112
rect 28960 23060 28994 23100
rect 27157 23035 27215 23041
rect 27157 23032 27169 23035
rect 27080 23004 27169 23032
rect 27157 23001 27169 23004
rect 27203 23032 27215 23035
rect 27893 23035 27951 23041
rect 27893 23032 27905 23035
rect 27203 23004 27905 23032
rect 27203 23001 27215 23004
rect 27157 22995 27215 23001
rect 27893 23001 27905 23004
rect 27939 23032 27951 23035
rect 28966 23032 28994 23060
rect 38626 23072 41328 23100
rect 30009 23035 30067 23041
rect 30009 23032 30021 23035
rect 27939 23004 28856 23032
rect 28966 23004 30021 23032
rect 27939 23001 27951 23004
rect 27893 22995 27951 23001
rect 28828 22976 28856 23004
rect 30009 23001 30021 23004
rect 30055 23032 30067 23035
rect 38626 23032 38654 23072
rect 41322 23060 41328 23072
rect 41380 23060 41386 23112
rect 46934 23060 46940 23112
rect 46992 23100 46998 23112
rect 47581 23103 47639 23109
rect 47581 23100 47593 23103
rect 46992 23072 47593 23100
rect 46992 23060 46998 23072
rect 47581 23069 47593 23072
rect 47627 23069 47639 23103
rect 47581 23063 47639 23069
rect 30055 23004 38654 23032
rect 30055 23001 30067 23004
rect 30009 22995 30067 23001
rect 26326 22964 26332 22976
rect 23799 22936 26188 22964
rect 26287 22936 26332 22964
rect 23799 22933 23811 22936
rect 23753 22927 23811 22933
rect 26326 22924 26332 22936
rect 26384 22964 26390 22976
rect 27065 22967 27123 22973
rect 27065 22964 27077 22967
rect 26384 22936 27077 22964
rect 26384 22924 26390 22936
rect 27065 22933 27077 22936
rect 27111 22933 27123 22967
rect 27430 22964 27436 22976
rect 27391 22936 27436 22964
rect 27065 22927 27123 22933
rect 27430 22924 27436 22936
rect 27488 22924 27494 22976
rect 27522 22924 27528 22976
rect 27580 22964 27586 22976
rect 28093 22967 28151 22973
rect 28093 22964 28105 22967
rect 27580 22936 28105 22964
rect 27580 22924 27586 22936
rect 28093 22933 28105 22936
rect 28139 22933 28151 22967
rect 28258 22964 28264 22976
rect 28219 22936 28264 22964
rect 28093 22927 28151 22933
rect 28258 22924 28264 22936
rect 28316 22924 28322 22976
rect 28810 22924 28816 22976
rect 28868 22924 28874 22976
rect 29546 22924 29552 22976
rect 29604 22964 29610 22976
rect 30101 22967 30159 22973
rect 30101 22964 30113 22967
rect 29604 22936 30113 22964
rect 29604 22924 29610 22936
rect 30101 22933 30113 22936
rect 30147 22933 30159 22967
rect 30101 22927 30159 22933
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 3694 22720 3700 22772
rect 3752 22760 3758 22772
rect 3752 22732 10180 22760
rect 3752 22720 3758 22732
rect 7009 22695 7067 22701
rect 7009 22661 7021 22695
rect 7055 22692 7067 22695
rect 7745 22695 7803 22701
rect 7745 22692 7757 22695
rect 7055 22664 7757 22692
rect 7055 22661 7067 22664
rect 7009 22655 7067 22661
rect 7745 22661 7757 22664
rect 7791 22661 7803 22695
rect 7745 22655 7803 22661
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22624 6975 22627
rect 7466 22624 7472 22636
rect 6963 22596 7472 22624
rect 6963 22593 6975 22596
rect 6917 22587 6975 22593
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 9401 22627 9459 22633
rect 9401 22593 9413 22627
rect 9447 22624 9459 22627
rect 9861 22627 9919 22633
rect 9447 22596 9536 22624
rect 9447 22593 9459 22596
rect 9401 22587 9459 22593
rect 7561 22559 7619 22565
rect 7561 22525 7573 22559
rect 7607 22556 7619 22559
rect 9306 22556 9312 22568
rect 7607 22528 9312 22556
rect 7607 22525 7619 22528
rect 7561 22519 7619 22525
rect 9306 22516 9312 22528
rect 9364 22516 9370 22568
rect 3510 22448 3516 22500
rect 3568 22488 3574 22500
rect 9508 22488 9536 22596
rect 9861 22593 9873 22627
rect 9907 22624 9919 22627
rect 9907 22596 10088 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 3568 22460 9536 22488
rect 3568 22448 3574 22460
rect 9950 22420 9956 22432
rect 9911 22392 9956 22420
rect 9950 22380 9956 22392
rect 10008 22380 10014 22432
rect 10060 22420 10088 22596
rect 10152 22488 10180 22732
rect 10226 22720 10232 22772
rect 10284 22760 10290 22772
rect 10873 22763 10931 22769
rect 10873 22760 10885 22763
rect 10284 22732 10885 22760
rect 10284 22720 10290 22732
rect 10873 22729 10885 22732
rect 10919 22729 10931 22763
rect 16114 22760 16120 22772
rect 16075 22732 16120 22760
rect 10873 22723 10931 22729
rect 16114 22720 16120 22732
rect 16172 22760 16178 22772
rect 16850 22760 16856 22772
rect 16172 22732 16856 22760
rect 16172 22720 16178 22732
rect 16850 22720 16856 22732
rect 16908 22720 16914 22772
rect 19334 22720 19340 22772
rect 19392 22760 19398 22772
rect 19797 22763 19855 22769
rect 19797 22760 19809 22763
rect 19392 22732 19809 22760
rect 19392 22720 19398 22732
rect 19797 22729 19809 22732
rect 19843 22729 19855 22763
rect 46750 22760 46756 22772
rect 19797 22723 19855 22729
rect 22066 22732 46756 22760
rect 13446 22652 13452 22704
rect 13504 22692 13510 22704
rect 13504 22664 15134 22692
rect 13504 22652 13510 22664
rect 10689 22627 10747 22633
rect 10689 22593 10701 22627
rect 10735 22624 10747 22627
rect 11422 22624 11428 22636
rect 10735 22596 11428 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 11422 22584 11428 22596
rect 11480 22584 11486 22636
rect 14366 22624 14372 22636
rect 14327 22596 14372 22624
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 16868 22624 16896 22720
rect 18598 22652 18604 22704
rect 18656 22692 18662 22704
rect 22066 22692 22094 22732
rect 46750 22720 46756 22732
rect 46808 22720 46814 22772
rect 47762 22720 47768 22772
rect 47820 22720 47826 22772
rect 25590 22692 25596 22704
rect 18656 22664 22094 22692
rect 25551 22664 25596 22692
rect 18656 22652 18662 22664
rect 25590 22652 25596 22664
rect 25648 22652 25654 22704
rect 25682 22652 25688 22704
rect 25740 22692 25746 22704
rect 27430 22692 27436 22704
rect 25740 22664 26464 22692
rect 25740 22652 25746 22664
rect 17405 22627 17463 22633
rect 17405 22624 17417 22627
rect 16868 22596 17417 22624
rect 17405 22593 17417 22596
rect 17451 22593 17463 22627
rect 17405 22587 17463 22593
rect 19610 22584 19616 22636
rect 19668 22624 19674 22636
rect 19705 22627 19763 22633
rect 19705 22624 19717 22627
rect 19668 22596 19717 22624
rect 19668 22584 19674 22596
rect 19705 22593 19717 22596
rect 19751 22593 19763 22627
rect 19705 22587 19763 22593
rect 19978 22584 19984 22636
rect 20036 22624 20042 22636
rect 20165 22627 20223 22633
rect 20165 22624 20177 22627
rect 20036 22596 20177 22624
rect 20036 22584 20042 22596
rect 20165 22593 20177 22596
rect 20211 22593 20223 22627
rect 20165 22587 20223 22593
rect 20717 22627 20775 22633
rect 20717 22593 20729 22627
rect 20763 22624 20775 22627
rect 20990 22624 20996 22636
rect 20763 22596 20996 22624
rect 20763 22593 20775 22596
rect 20717 22587 20775 22593
rect 20990 22584 20996 22596
rect 21048 22584 21054 22636
rect 21913 22627 21971 22633
rect 21913 22624 21925 22627
rect 21192 22596 21925 22624
rect 11514 22556 11520 22568
rect 11475 22528 11520 22556
rect 11514 22516 11520 22528
rect 11572 22516 11578 22568
rect 11698 22556 11704 22568
rect 11659 22528 11704 22556
rect 11698 22516 11704 22528
rect 11756 22516 11762 22568
rect 11977 22559 12035 22565
rect 11977 22525 11989 22559
rect 12023 22525 12035 22559
rect 11977 22519 12035 22525
rect 14645 22559 14703 22565
rect 14645 22525 14657 22559
rect 14691 22556 14703 22559
rect 15930 22556 15936 22568
rect 14691 22528 15936 22556
rect 14691 22525 14703 22528
rect 14645 22519 14703 22525
rect 11992 22488 12020 22519
rect 15930 22516 15936 22528
rect 15988 22516 15994 22568
rect 17586 22556 17592 22568
rect 17547 22528 17592 22556
rect 17586 22516 17592 22528
rect 17644 22516 17650 22568
rect 19150 22556 19156 22568
rect 19111 22528 19156 22556
rect 19150 22516 19156 22528
rect 19208 22516 19214 22568
rect 10152 22460 12020 22488
rect 10410 22420 10416 22432
rect 10060 22392 10416 22420
rect 10410 22380 10416 22392
rect 10468 22420 10474 22432
rect 11974 22420 11980 22432
rect 10468 22392 11980 22420
rect 10468 22380 10474 22392
rect 11974 22380 11980 22392
rect 12032 22380 12038 22432
rect 20254 22420 20260 22432
rect 20215 22392 20260 22420
rect 20254 22380 20260 22392
rect 20312 22380 20318 22432
rect 20714 22380 20720 22432
rect 20772 22420 20778 22432
rect 21192 22429 21220 22596
rect 21913 22593 21925 22596
rect 21959 22593 21971 22627
rect 21913 22587 21971 22593
rect 22830 22584 22836 22636
rect 22888 22624 22894 22636
rect 23017 22627 23075 22633
rect 23017 22624 23029 22627
rect 22888 22596 23029 22624
rect 22888 22584 22894 22596
rect 23017 22593 23029 22596
rect 23063 22593 23075 22627
rect 23017 22587 23075 22593
rect 24210 22584 24216 22636
rect 24268 22624 24274 22636
rect 24673 22627 24731 22633
rect 24673 22624 24685 22627
rect 24268 22596 24685 22624
rect 24268 22584 24274 22596
rect 24673 22593 24685 22596
rect 24719 22624 24731 22627
rect 24719 22596 25452 22624
rect 24719 22593 24731 22596
rect 24673 22587 24731 22593
rect 22465 22559 22523 22565
rect 22465 22525 22477 22559
rect 22511 22556 22523 22559
rect 22554 22556 22560 22568
rect 22511 22528 22560 22556
rect 22511 22525 22523 22528
rect 22465 22519 22523 22525
rect 22554 22516 22560 22528
rect 22612 22516 22618 22568
rect 24765 22559 24823 22565
rect 24765 22525 24777 22559
rect 24811 22525 24823 22559
rect 24765 22519 24823 22525
rect 24780 22488 24808 22519
rect 24854 22516 24860 22568
rect 24912 22556 24918 22568
rect 25041 22559 25099 22565
rect 25041 22556 25053 22559
rect 24912 22528 25053 22556
rect 24912 22516 24918 22528
rect 25041 22525 25053 22528
rect 25087 22525 25099 22559
rect 25424 22556 25452 22596
rect 25498 22584 25504 22636
rect 25556 22624 25562 22636
rect 25556 22596 25601 22624
rect 25556 22584 25562 22596
rect 26142 22584 26148 22636
rect 26200 22624 26206 22636
rect 26436 22633 26464 22664
rect 27172 22664 27436 22692
rect 27172 22633 27200 22664
rect 27430 22652 27436 22664
rect 27488 22652 27494 22704
rect 27706 22652 27712 22704
rect 27764 22692 27770 22704
rect 28350 22692 28356 22704
rect 27764 22664 28356 22692
rect 27764 22652 27770 22664
rect 28350 22652 28356 22664
rect 28408 22652 28414 22704
rect 29641 22695 29699 22701
rect 29641 22661 29653 22695
rect 29687 22692 29699 22695
rect 29914 22692 29920 22704
rect 29687 22664 29920 22692
rect 29687 22661 29699 22664
rect 29641 22655 29699 22661
rect 29914 22652 29920 22664
rect 29972 22652 29978 22704
rect 47780 22692 47808 22720
rect 35866 22664 47808 22692
rect 26329 22627 26387 22633
rect 26200 22596 26245 22624
rect 26200 22584 26206 22596
rect 26329 22593 26341 22627
rect 26375 22593 26387 22627
rect 26329 22587 26387 22593
rect 26421 22627 26479 22633
rect 26421 22593 26433 22627
rect 26467 22593 26479 22627
rect 26421 22587 26479 22593
rect 27157 22627 27215 22633
rect 27157 22593 27169 22627
rect 27203 22593 27215 22627
rect 27157 22587 27215 22593
rect 26234 22556 26240 22568
rect 25424 22528 26240 22556
rect 25041 22519 25099 22525
rect 26234 22516 26240 22528
rect 26292 22556 26298 22568
rect 26344 22556 26372 22587
rect 26436 22556 26464 22587
rect 27246 22584 27252 22636
rect 27304 22624 27310 22636
rect 27304 22596 27349 22624
rect 27304 22584 27310 22596
rect 27614 22584 27620 22636
rect 27672 22624 27678 22636
rect 28442 22624 28448 22636
rect 27672 22596 28448 22624
rect 27672 22584 27678 22596
rect 28442 22584 28448 22596
rect 28500 22624 28506 22636
rect 28626 22624 28632 22636
rect 28500 22596 28632 22624
rect 28500 22584 28506 22596
rect 28626 22584 28632 22596
rect 28684 22624 28690 22636
rect 29546 22624 29552 22636
rect 28684 22596 29552 22624
rect 28684 22584 28690 22596
rect 29546 22584 29552 22596
rect 29604 22584 29610 22636
rect 28258 22556 28264 22568
rect 26292 22528 26385 22556
rect 26436 22528 28264 22556
rect 26292 22516 26298 22528
rect 28258 22516 28264 22528
rect 28316 22516 28322 22568
rect 25682 22488 25688 22500
rect 24780 22460 25688 22488
rect 25682 22448 25688 22460
rect 25740 22448 25746 22500
rect 26050 22448 26056 22500
rect 26108 22488 26114 22500
rect 26970 22488 26976 22500
rect 26108 22460 26976 22488
rect 26108 22448 26114 22460
rect 26970 22448 26976 22460
rect 27028 22488 27034 22500
rect 28994 22488 29000 22500
rect 27028 22460 29000 22488
rect 27028 22448 27034 22460
rect 28994 22448 29000 22460
rect 29052 22448 29058 22500
rect 35866 22488 35894 22664
rect 45830 22584 45836 22636
rect 45888 22624 45894 22636
rect 46477 22627 46535 22633
rect 46477 22624 46489 22627
rect 45888 22596 46489 22624
rect 45888 22584 45894 22596
rect 46477 22593 46489 22596
rect 46523 22593 46535 22627
rect 46477 22587 46535 22593
rect 46842 22584 46848 22636
rect 46900 22624 46906 22636
rect 47765 22627 47823 22633
rect 47765 22624 47777 22627
rect 46900 22596 47777 22624
rect 46900 22584 46906 22596
rect 47765 22593 47777 22596
rect 47811 22593 47823 22627
rect 47765 22587 47823 22593
rect 46201 22559 46259 22565
rect 46201 22525 46213 22559
rect 46247 22556 46259 22559
rect 46566 22556 46572 22568
rect 46247 22528 46572 22556
rect 46247 22525 46259 22528
rect 46201 22519 46259 22525
rect 46566 22516 46572 22528
rect 46624 22516 46630 22568
rect 31726 22460 35894 22488
rect 21177 22423 21235 22429
rect 21177 22420 21189 22423
rect 20772 22392 21189 22420
rect 20772 22380 20778 22392
rect 21177 22389 21189 22392
rect 21223 22389 21235 22423
rect 23198 22420 23204 22432
rect 23159 22392 23204 22420
rect 21177 22383 21235 22389
rect 23198 22380 23204 22392
rect 23256 22380 23262 22432
rect 26145 22423 26203 22429
rect 26145 22389 26157 22423
rect 26191 22420 26203 22423
rect 26602 22420 26608 22432
rect 26191 22392 26608 22420
rect 26191 22389 26203 22392
rect 26145 22383 26203 22389
rect 26602 22380 26608 22392
rect 26660 22380 26666 22432
rect 26878 22380 26884 22432
rect 26936 22420 26942 22432
rect 27433 22423 27491 22429
rect 27433 22420 27445 22423
rect 26936 22392 27445 22420
rect 26936 22380 26942 22392
rect 27433 22389 27445 22392
rect 27479 22389 27491 22423
rect 27433 22383 27491 22389
rect 27522 22380 27528 22432
rect 27580 22420 27586 22432
rect 31726 22420 31754 22460
rect 27580 22392 31754 22420
rect 27580 22380 27586 22392
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 11241 22219 11299 22225
rect 11241 22185 11253 22219
rect 11287 22216 11299 22219
rect 11698 22216 11704 22228
rect 11287 22188 11704 22216
rect 11287 22185 11299 22188
rect 11241 22179 11299 22185
rect 11698 22176 11704 22188
rect 11756 22176 11762 22228
rect 11790 22176 11796 22228
rect 11848 22216 11854 22228
rect 13265 22219 13323 22225
rect 13265 22216 13277 22219
rect 11848 22188 13277 22216
rect 11848 22176 11854 22188
rect 13265 22185 13277 22188
rect 13311 22185 13323 22219
rect 13265 22179 13323 22185
rect 13998 22176 14004 22228
rect 14056 22216 14062 22228
rect 14277 22219 14335 22225
rect 14277 22216 14289 22219
rect 14056 22188 14289 22216
rect 14056 22176 14062 22188
rect 14277 22185 14289 22188
rect 14323 22185 14335 22219
rect 17586 22216 17592 22228
rect 17547 22188 17592 22216
rect 14277 22179 14335 22185
rect 17586 22176 17592 22188
rect 17644 22176 17650 22228
rect 22830 22216 22836 22228
rect 22743 22188 22836 22216
rect 22830 22176 22836 22188
rect 22888 22216 22894 22228
rect 43162 22216 43168 22228
rect 22888 22188 43168 22216
rect 22888 22176 22894 22188
rect 43162 22176 43168 22188
rect 43220 22176 43226 22228
rect 16022 22148 16028 22160
rect 15672 22120 16028 22148
rect 8938 22080 8944 22092
rect 8899 22052 8944 22080
rect 8938 22040 8944 22052
rect 8996 22040 9002 22092
rect 11422 22040 11428 22092
rect 11480 22080 11486 22092
rect 12250 22080 12256 22092
rect 11480 22052 12256 22080
rect 11480 22040 11486 22052
rect 12250 22040 12256 22052
rect 12308 22080 12314 22092
rect 15473 22083 15531 22089
rect 12308 22052 14136 22080
rect 12308 22040 12314 22052
rect 7558 22012 7564 22024
rect 7519 21984 7564 22012
rect 7558 21972 7564 21984
rect 7616 21972 7622 22024
rect 11146 22012 11152 22024
rect 11107 21984 11152 22012
rect 11146 21972 11152 21984
rect 11204 21972 11210 22024
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 22012 11851 22015
rect 11882 22012 11888 22024
rect 11839 21984 11888 22012
rect 11839 21981 11851 21984
rect 11793 21975 11851 21981
rect 11882 21972 11888 21984
rect 11940 21972 11946 22024
rect 14108 22021 14136 22052
rect 15473 22049 15485 22083
rect 15519 22080 15531 22083
rect 15672 22080 15700 22120
rect 16022 22108 16028 22120
rect 16080 22108 16086 22160
rect 22554 22108 22560 22160
rect 22612 22148 22618 22160
rect 27246 22148 27252 22160
rect 22612 22120 27252 22148
rect 22612 22108 22618 22120
rect 27246 22108 27252 22120
rect 27304 22108 27310 22160
rect 15930 22080 15936 22092
rect 15519 22052 15700 22080
rect 15891 22052 15936 22080
rect 15519 22049 15531 22052
rect 15473 22043 15531 22049
rect 15930 22040 15936 22052
rect 15988 22040 15994 22092
rect 16666 22040 16672 22092
rect 16724 22080 16730 22092
rect 20806 22080 20812 22092
rect 16724 22052 20812 22080
rect 16724 22040 16730 22052
rect 20806 22040 20812 22052
rect 20864 22040 20870 22092
rect 23934 22040 23940 22092
rect 23992 22080 23998 22092
rect 27614 22080 27620 22092
rect 23992 22052 27620 22080
rect 23992 22040 23998 22052
rect 27614 22040 27620 22052
rect 27672 22040 27678 22092
rect 28994 22080 29000 22092
rect 28955 22052 29000 22080
rect 28994 22040 29000 22052
rect 29052 22040 29058 22092
rect 46477 22083 46535 22089
rect 46477 22049 46489 22083
rect 46523 22080 46535 22083
rect 46934 22080 46940 22092
rect 46523 22052 46940 22080
rect 46523 22049 46535 22052
rect 46477 22043 46535 22049
rect 46934 22040 46940 22052
rect 46992 22040 46998 22092
rect 47118 22080 47124 22092
rect 47079 22052 47124 22080
rect 47118 22040 47124 22052
rect 47176 22080 47182 22092
rect 47762 22080 47768 22092
rect 47176 22052 47768 22080
rect 47176 22040 47182 22052
rect 47762 22040 47768 22052
rect 47820 22040 47826 22092
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 15565 22015 15623 22021
rect 15565 21981 15577 22015
rect 15611 22012 15623 22015
rect 16114 22012 16120 22024
rect 15611 21984 16120 22012
rect 15611 21981 15623 21984
rect 15565 21975 15623 21981
rect 16114 21972 16120 21984
rect 16172 21972 16178 22024
rect 17494 22012 17500 22024
rect 17455 21984 17500 22012
rect 17494 21972 17500 21984
rect 17552 22012 17558 22024
rect 19610 22012 19616 22024
rect 17552 21984 19616 22012
rect 17552 21972 17558 21984
rect 19610 21972 19616 21984
rect 19668 21972 19674 22024
rect 19705 22015 19763 22021
rect 19705 21981 19717 22015
rect 19751 22012 19763 22015
rect 20162 22012 20168 22024
rect 19751 21984 20168 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 20162 21972 20168 21984
rect 20220 21972 20226 22024
rect 20441 22015 20499 22021
rect 20441 21981 20453 22015
rect 20487 22012 20499 22015
rect 24762 22012 24768 22024
rect 20487 21984 20852 22012
rect 24723 21984 24768 22012
rect 20487 21981 20499 21984
rect 20441 21975 20499 21981
rect 9214 21944 9220 21956
rect 9175 21916 9220 21944
rect 9214 21904 9220 21916
rect 9272 21904 9278 21956
rect 9950 21904 9956 21956
rect 10008 21904 10014 21956
rect 11514 21904 11520 21956
rect 11572 21944 11578 21956
rect 13081 21947 13139 21953
rect 13081 21944 13093 21947
rect 11572 21916 13093 21944
rect 11572 21904 11578 21916
rect 13081 21913 13093 21916
rect 13127 21913 13139 21947
rect 13081 21907 13139 21913
rect 13297 21947 13355 21953
rect 13297 21913 13309 21947
rect 13343 21944 13355 21947
rect 14918 21944 14924 21956
rect 13343 21916 14924 21944
rect 13343 21913 13355 21916
rect 13297 21907 13355 21913
rect 14918 21904 14924 21916
rect 14976 21904 14982 21956
rect 7466 21836 7472 21888
rect 7524 21876 7530 21888
rect 7653 21879 7711 21885
rect 7653 21876 7665 21879
rect 7524 21848 7665 21876
rect 7524 21836 7530 21848
rect 7653 21845 7665 21848
rect 7699 21845 7711 21879
rect 7653 21839 7711 21845
rect 9306 21836 9312 21888
rect 9364 21876 9370 21888
rect 10689 21879 10747 21885
rect 10689 21876 10701 21879
rect 9364 21848 10701 21876
rect 9364 21836 9370 21848
rect 10689 21845 10701 21848
rect 10735 21845 10747 21879
rect 10689 21839 10747 21845
rect 11698 21836 11704 21888
rect 11756 21876 11762 21888
rect 11974 21876 11980 21888
rect 11756 21848 11980 21876
rect 11756 21836 11762 21848
rect 11974 21836 11980 21848
rect 12032 21836 12038 21888
rect 13449 21879 13507 21885
rect 13449 21845 13461 21879
rect 13495 21876 13507 21879
rect 13630 21876 13636 21888
rect 13495 21848 13636 21876
rect 13495 21845 13507 21848
rect 13449 21839 13507 21845
rect 13630 21836 13636 21848
rect 13688 21836 13694 21888
rect 19628 21876 19656 21972
rect 20824 21956 20852 21984
rect 24762 21972 24768 21984
rect 24820 21972 24826 22024
rect 26602 22012 26608 22024
rect 26563 21984 26608 22012
rect 26602 21972 26608 21984
rect 26660 21972 26666 22024
rect 26789 22015 26847 22021
rect 26789 21981 26801 22015
rect 26835 22012 26847 22015
rect 26878 22012 26884 22024
rect 26835 21984 26884 22012
rect 26835 21981 26847 21984
rect 26789 21975 26847 21981
rect 26878 21972 26884 21984
rect 26936 21972 26942 22024
rect 27246 22012 27252 22024
rect 27207 21984 27252 22012
rect 27246 21972 27252 21984
rect 27304 21972 27310 22024
rect 46293 22015 46351 22021
rect 46293 21981 46305 22015
rect 46339 21981 46351 22015
rect 46293 21975 46351 21981
rect 20717 21947 20775 21953
rect 20717 21913 20729 21947
rect 20763 21913 20775 21947
rect 20717 21907 20775 21913
rect 19889 21879 19947 21885
rect 19889 21876 19901 21879
rect 19628 21848 19901 21876
rect 19889 21845 19901 21848
rect 19935 21845 19947 21879
rect 20732 21876 20760 21907
rect 20806 21904 20812 21956
rect 20864 21944 20870 21956
rect 21082 21944 21088 21956
rect 20864 21916 21088 21944
rect 20864 21904 20870 21916
rect 21082 21904 21088 21916
rect 21140 21944 21146 21956
rect 21361 21947 21419 21953
rect 21361 21944 21373 21947
rect 21140 21916 21373 21944
rect 21140 21904 21146 21916
rect 21361 21913 21373 21916
rect 21407 21913 21419 21947
rect 21361 21907 21419 21913
rect 26697 21947 26755 21953
rect 26697 21913 26709 21947
rect 26743 21944 26755 21947
rect 27525 21947 27583 21953
rect 27525 21944 27537 21947
rect 26743 21916 27537 21944
rect 26743 21913 26755 21916
rect 26697 21907 26755 21913
rect 27525 21913 27537 21916
rect 27571 21913 27583 21947
rect 27525 21907 27583 21913
rect 28534 21904 28540 21956
rect 28592 21904 28598 21956
rect 46308 21944 46336 21975
rect 46750 21944 46756 21956
rect 46308 21916 46756 21944
rect 46750 21904 46756 21916
rect 46808 21904 46814 21956
rect 21542 21876 21548 21888
rect 20732 21848 21548 21876
rect 19889 21839 19947 21845
rect 21542 21836 21548 21848
rect 21600 21836 21606 21888
rect 24949 21879 25007 21885
rect 24949 21845 24961 21879
rect 24995 21876 25007 21879
rect 26970 21876 26976 21888
rect 24995 21848 26976 21876
rect 24995 21845 25007 21848
rect 24949 21839 25007 21845
rect 26970 21836 26976 21848
rect 27028 21836 27034 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 9122 21672 9128 21684
rect 7300 21644 9128 21672
rect 7300 21545 7328 21644
rect 9122 21632 9128 21644
rect 9180 21632 9186 21684
rect 9214 21632 9220 21684
rect 9272 21672 9278 21684
rect 9585 21675 9643 21681
rect 9585 21672 9597 21675
rect 9272 21644 9597 21672
rect 9272 21632 9278 21644
rect 9585 21641 9597 21644
rect 9631 21641 9643 21675
rect 9766 21672 9772 21684
rect 9727 21644 9772 21672
rect 9585 21635 9643 21641
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 17494 21672 17500 21684
rect 9876 21644 17500 21672
rect 7466 21604 7472 21616
rect 7427 21576 7472 21604
rect 7466 21564 7472 21576
rect 7524 21564 7530 21616
rect 7558 21564 7564 21616
rect 7616 21604 7622 21616
rect 9876 21604 9904 21644
rect 17494 21632 17500 21644
rect 17552 21632 17558 21684
rect 20162 21632 20168 21684
rect 20220 21672 20226 21684
rect 21177 21675 21235 21681
rect 21177 21672 21189 21675
rect 20220 21644 21189 21672
rect 20220 21632 20226 21644
rect 21177 21641 21189 21644
rect 21223 21641 21235 21675
rect 21177 21635 21235 21641
rect 7616 21576 9904 21604
rect 10689 21607 10747 21613
rect 7616 21564 7622 21576
rect 10689 21573 10701 21607
rect 10735 21604 10747 21607
rect 11514 21604 11520 21616
rect 10735 21576 11520 21604
rect 10735 21573 10747 21576
rect 10689 21567 10747 21573
rect 11514 21564 11520 21576
rect 11572 21564 11578 21616
rect 18966 21604 18972 21616
rect 18616 21576 18972 21604
rect 7285 21539 7343 21545
rect 7285 21505 7297 21539
rect 7331 21505 7343 21539
rect 7285 21499 7343 21505
rect 9766 21539 9824 21545
rect 9766 21505 9778 21539
rect 9812 21536 9824 21539
rect 10873 21539 10931 21545
rect 10873 21536 10885 21539
rect 9812 21508 10885 21536
rect 9812 21505 9824 21508
rect 9766 21499 9824 21505
rect 10873 21505 10885 21508
rect 10919 21505 10931 21539
rect 10873 21499 10931 21505
rect 7745 21471 7803 21477
rect 7745 21437 7757 21471
rect 7791 21437 7803 21471
rect 7745 21431 7803 21437
rect 14 21360 20 21412
rect 72 21400 78 21412
rect 7760 21400 7788 21431
rect 9306 21428 9312 21480
rect 9364 21468 9370 21480
rect 10137 21471 10195 21477
rect 10137 21468 10149 21471
rect 9364 21440 10149 21468
rect 9364 21428 9370 21440
rect 10137 21437 10149 21440
rect 10183 21437 10195 21471
rect 10137 21431 10195 21437
rect 10226 21428 10232 21480
rect 10284 21468 10290 21480
rect 10888 21468 10916 21499
rect 10962 21496 10968 21548
rect 11020 21536 11026 21548
rect 11020 21508 11065 21536
rect 11020 21496 11026 21508
rect 11882 21496 11888 21548
rect 11940 21536 11946 21548
rect 12342 21536 12348 21548
rect 11940 21508 12348 21536
rect 11940 21496 11946 21508
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 14734 21496 14740 21548
rect 14792 21536 14798 21548
rect 16666 21536 16672 21548
rect 14792 21508 16672 21536
rect 14792 21496 14798 21508
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 18616 21545 18644 21576
rect 18966 21564 18972 21576
rect 19024 21564 19030 21616
rect 20254 21604 20260 21616
rect 20102 21576 20260 21604
rect 20254 21564 20260 21576
rect 20312 21564 20318 21616
rect 20990 21564 20996 21616
rect 21048 21604 21054 21616
rect 21085 21607 21143 21613
rect 21085 21604 21097 21607
rect 21048 21576 21097 21604
rect 21048 21564 21054 21576
rect 21085 21573 21097 21576
rect 21131 21573 21143 21607
rect 21085 21567 21143 21573
rect 18601 21539 18659 21545
rect 18601 21505 18613 21539
rect 18647 21505 18659 21539
rect 21192 21536 21220 21635
rect 26970 21632 26976 21684
rect 27028 21672 27034 21684
rect 27028 21644 27200 21672
rect 27028 21632 27034 21644
rect 27172 21604 27200 21644
rect 27246 21632 27252 21684
rect 27304 21672 27310 21684
rect 27525 21675 27583 21681
rect 27525 21672 27537 21675
rect 27304 21644 27537 21672
rect 27304 21632 27310 21644
rect 27525 21641 27537 21644
rect 27571 21641 27583 21675
rect 28534 21672 28540 21684
rect 28495 21644 28540 21672
rect 27525 21635 27583 21641
rect 28534 21632 28540 21644
rect 28592 21632 28598 21684
rect 47946 21604 47952 21616
rect 27172 21576 28488 21604
rect 47907 21576 47952 21604
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21192 21508 21833 21536
rect 18601 21499 18659 21505
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 23934 21536 23940 21548
rect 23895 21508 23940 21536
rect 21821 21499 21879 21505
rect 23934 21496 23940 21508
rect 23992 21496 23998 21548
rect 24854 21496 24860 21548
rect 24912 21536 24918 21548
rect 24949 21539 25007 21545
rect 24949 21536 24961 21539
rect 24912 21508 24961 21536
rect 24912 21496 24918 21508
rect 24949 21505 24961 21508
rect 24995 21505 25007 21539
rect 24949 21499 25007 21505
rect 26694 21496 26700 21548
rect 26752 21536 26758 21548
rect 28460 21545 28488 21576
rect 47946 21564 47952 21576
rect 48004 21564 48010 21616
rect 27341 21539 27399 21545
rect 27341 21536 27353 21539
rect 26752 21508 27353 21536
rect 26752 21496 26758 21508
rect 27341 21505 27353 21508
rect 27387 21505 27399 21539
rect 27341 21499 27399 21505
rect 28445 21539 28503 21545
rect 28445 21505 28457 21539
rect 28491 21505 28503 21539
rect 28445 21499 28503 21505
rect 11054 21468 11060 21480
rect 10284 21440 10329 21468
rect 10888 21440 11060 21468
rect 10284 21428 10290 21440
rect 11054 21428 11060 21440
rect 11112 21468 11118 21480
rect 11790 21468 11796 21480
rect 11112 21440 11796 21468
rect 11112 21428 11118 21440
rect 11790 21428 11796 21440
rect 11848 21428 11854 21480
rect 16574 21428 16580 21480
rect 16632 21468 16638 21480
rect 16945 21471 17003 21477
rect 16945 21468 16957 21471
rect 16632 21440 16957 21468
rect 16632 21428 16638 21440
rect 16945 21437 16957 21440
rect 16991 21468 17003 21471
rect 17402 21468 17408 21480
rect 16991 21440 17408 21468
rect 16991 21437 17003 21440
rect 16945 21431 17003 21437
rect 17402 21428 17408 21440
rect 17460 21428 17466 21480
rect 18874 21468 18880 21480
rect 18835 21440 18880 21468
rect 18874 21428 18880 21440
rect 18932 21428 18938 21480
rect 18966 21428 18972 21480
rect 19024 21468 19030 21480
rect 22370 21468 22376 21480
rect 19024 21440 22376 21468
rect 19024 21428 19030 21440
rect 22370 21428 22376 21440
rect 22428 21428 22434 21480
rect 22554 21468 22560 21480
rect 22515 21440 22560 21468
rect 22554 21428 22560 21440
rect 22612 21428 22618 21480
rect 25041 21471 25099 21477
rect 25041 21437 25053 21471
rect 25087 21468 25099 21471
rect 27522 21468 27528 21480
rect 25087 21440 27528 21468
rect 25087 21437 25099 21440
rect 25041 21431 25099 21437
rect 27522 21428 27528 21440
rect 27580 21428 27586 21480
rect 72 21372 7788 21400
rect 72 21360 78 21372
rect 9674 21360 9680 21412
rect 9732 21400 9738 21412
rect 10689 21403 10747 21409
rect 10689 21400 10701 21403
rect 9732 21372 10701 21400
rect 9732 21360 9738 21372
rect 10689 21369 10701 21372
rect 10735 21369 10747 21403
rect 22572 21400 22600 21428
rect 46474 21400 46480 21412
rect 22572 21372 46480 21400
rect 10689 21363 10747 21369
rect 46474 21360 46480 21372
rect 46532 21360 46538 21412
rect 9766 21292 9772 21344
rect 9824 21332 9830 21344
rect 10318 21332 10324 21344
rect 9824 21304 10324 21332
rect 9824 21292 9830 21304
rect 10318 21292 10324 21304
rect 10376 21332 10382 21344
rect 10962 21332 10968 21344
rect 10376 21304 10968 21332
rect 10376 21292 10382 21304
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 11974 21292 11980 21344
rect 12032 21332 12038 21344
rect 12250 21332 12256 21344
rect 12032 21304 12256 21332
rect 12032 21292 12038 21304
rect 12250 21292 12256 21304
rect 12308 21332 12314 21344
rect 20349 21335 20407 21341
rect 20349 21332 20361 21335
rect 12308 21304 20361 21332
rect 12308 21292 12314 21304
rect 20349 21301 20361 21304
rect 20395 21332 20407 21335
rect 20438 21332 20444 21344
rect 20395 21304 20444 21332
rect 20395 21301 20407 21304
rect 20349 21295 20407 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 24029 21335 24087 21341
rect 24029 21301 24041 21335
rect 24075 21332 24087 21335
rect 24762 21332 24768 21344
rect 24075 21304 24768 21332
rect 24075 21301 24087 21304
rect 24029 21295 24087 21301
rect 24762 21292 24768 21304
rect 24820 21292 24826 21344
rect 25314 21332 25320 21344
rect 25275 21304 25320 21332
rect 25314 21292 25320 21304
rect 25372 21292 25378 21344
rect 25958 21292 25964 21344
rect 26016 21332 26022 21344
rect 48041 21335 48099 21341
rect 48041 21332 48053 21335
rect 26016 21304 48053 21332
rect 26016 21292 26022 21304
rect 48041 21301 48053 21304
rect 48087 21301 48099 21335
rect 48041 21295 48099 21301
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 9953 21131 10011 21137
rect 9953 21097 9965 21131
rect 9999 21128 10011 21131
rect 10594 21128 10600 21140
rect 9999 21100 10600 21128
rect 9999 21097 10011 21100
rect 9953 21091 10011 21097
rect 10594 21088 10600 21100
rect 10652 21088 10658 21140
rect 10778 21128 10784 21140
rect 10739 21100 10784 21128
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 10962 21088 10968 21140
rect 11020 21128 11026 21140
rect 11609 21131 11667 21137
rect 11609 21128 11621 21131
rect 11020 21100 11621 21128
rect 11020 21088 11026 21100
rect 11609 21097 11621 21100
rect 11655 21097 11667 21131
rect 14918 21128 14924 21140
rect 14879 21100 14924 21128
rect 11609 21091 11667 21097
rect 14918 21088 14924 21100
rect 14976 21088 14982 21140
rect 18601 21131 18659 21137
rect 18601 21097 18613 21131
rect 18647 21128 18659 21131
rect 18874 21128 18880 21140
rect 18647 21100 18880 21128
rect 18647 21097 18659 21100
rect 18601 21091 18659 21097
rect 18874 21088 18880 21100
rect 18932 21088 18938 21140
rect 22925 21131 22983 21137
rect 22066 21100 22876 21128
rect 10137 21063 10195 21069
rect 10137 21029 10149 21063
rect 10183 21060 10195 21063
rect 11054 21060 11060 21072
rect 10183 21032 11060 21060
rect 10183 21029 10195 21032
rect 10137 21023 10195 21029
rect 11054 21020 11060 21032
rect 11112 21020 11118 21072
rect 11146 21020 11152 21072
rect 11204 21060 11210 21072
rect 20346 21060 20352 21072
rect 11204 21032 20352 21060
rect 11204 21020 11210 21032
rect 20346 21020 20352 21032
rect 20404 21060 20410 21072
rect 20441 21063 20499 21069
rect 20441 21060 20453 21063
rect 20404 21032 20453 21060
rect 20404 21020 20410 21032
rect 20441 21029 20453 21032
rect 20487 21029 20499 21063
rect 22066 21060 22094 21100
rect 20441 21023 20499 21029
rect 20548 21032 22094 21060
rect 3602 20952 3608 21004
rect 3660 20992 3666 21004
rect 20548 20992 20576 21032
rect 22848 20992 22876 21100
rect 22925 21097 22937 21131
rect 22971 21128 22983 21131
rect 23014 21128 23020 21140
rect 22971 21100 23020 21128
rect 22971 21097 22983 21100
rect 22925 21091 22983 21097
rect 23014 21088 23020 21100
rect 23072 21128 23078 21140
rect 26694 21128 26700 21140
rect 23072 21100 26700 21128
rect 23072 21088 23078 21100
rect 26694 21088 26700 21100
rect 26752 21088 26758 21140
rect 24857 20995 24915 21001
rect 24857 20992 24869 20995
rect 3660 20964 20576 20992
rect 20824 20964 22094 20992
rect 22848 20964 24869 20992
rect 3660 20952 3666 20964
rect 14090 20924 14096 20936
rect 14051 20896 14096 20924
rect 14090 20884 14096 20896
rect 14148 20884 14154 20936
rect 18414 20884 18420 20936
rect 18472 20924 18478 20936
rect 18509 20927 18567 20933
rect 18509 20924 18521 20927
rect 18472 20896 18521 20924
rect 18472 20884 18478 20896
rect 18509 20893 18521 20896
rect 18555 20893 18567 20927
rect 19242 20924 19248 20936
rect 19203 20896 19248 20924
rect 18509 20887 18567 20893
rect 19242 20884 19248 20896
rect 19300 20884 19306 20936
rect 20162 20884 20168 20936
rect 20220 20924 20226 20936
rect 20257 20927 20315 20933
rect 20257 20924 20269 20927
rect 20220 20896 20269 20924
rect 20220 20884 20226 20896
rect 20257 20893 20269 20896
rect 20303 20893 20315 20927
rect 20257 20887 20315 20893
rect 9306 20816 9312 20868
rect 9364 20856 9370 20868
rect 9769 20859 9827 20865
rect 9769 20856 9781 20859
rect 9364 20828 9781 20856
rect 9364 20816 9370 20828
rect 9769 20825 9781 20828
rect 9815 20825 9827 20859
rect 10594 20856 10600 20868
rect 10555 20828 10600 20856
rect 9769 20819 9827 20825
rect 10594 20816 10600 20828
rect 10652 20816 10658 20868
rect 10813 20859 10871 20865
rect 10813 20825 10825 20859
rect 10859 20856 10871 20859
rect 11517 20859 11575 20865
rect 11517 20856 11529 20859
rect 10859 20828 11529 20856
rect 10859 20825 10871 20828
rect 10813 20819 10871 20825
rect 11517 20825 11529 20828
rect 11563 20856 11575 20859
rect 14734 20856 14740 20868
rect 11563 20828 14320 20856
rect 14695 20828 14740 20856
rect 11563 20825 11575 20828
rect 11517 20819 11575 20825
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 9969 20791 10027 20797
rect 9969 20788 9981 20791
rect 9732 20760 9981 20788
rect 9732 20748 9738 20760
rect 9969 20757 9981 20760
rect 10015 20757 10027 20791
rect 9969 20751 10027 20757
rect 10226 20748 10232 20800
rect 10284 20788 10290 20800
rect 10965 20791 11023 20797
rect 10965 20788 10977 20791
rect 10284 20760 10977 20788
rect 10284 20748 10290 20760
rect 10965 20757 10977 20760
rect 11011 20757 11023 20791
rect 14182 20788 14188 20800
rect 14143 20760 14188 20788
rect 10965 20751 11023 20757
rect 14182 20748 14188 20760
rect 14240 20748 14246 20800
rect 14292 20788 14320 20828
rect 14734 20816 14740 20828
rect 14792 20816 14798 20868
rect 14953 20859 15011 20865
rect 14953 20825 14965 20859
rect 14999 20856 15011 20859
rect 15654 20856 15660 20868
rect 14999 20828 15660 20856
rect 14999 20825 15011 20828
rect 14953 20819 15011 20825
rect 15654 20816 15660 20828
rect 15712 20816 15718 20868
rect 20272 20856 20300 20887
rect 20438 20884 20444 20936
rect 20496 20924 20502 20936
rect 20824 20924 20852 20964
rect 21082 20924 21088 20936
rect 20496 20896 20852 20924
rect 21043 20896 21088 20924
rect 20496 20884 20502 20896
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 22066 20924 22094 20964
rect 24857 20961 24869 20964
rect 24903 20961 24915 20995
rect 24857 20955 24915 20961
rect 26878 20952 26884 21004
rect 26936 20992 26942 21004
rect 27430 20992 27436 21004
rect 26936 20964 27436 20992
rect 26936 20952 26942 20964
rect 27430 20952 27436 20964
rect 27488 20952 27494 21004
rect 27893 20995 27951 21001
rect 27893 20961 27905 20995
rect 27939 20992 27951 20995
rect 28074 20992 28080 21004
rect 27939 20964 28080 20992
rect 27939 20961 27951 20964
rect 27893 20955 27951 20961
rect 28074 20952 28080 20964
rect 28132 20952 28138 21004
rect 32214 20992 32220 21004
rect 32175 20964 32220 20992
rect 32214 20952 32220 20964
rect 32272 20952 32278 21004
rect 46293 20995 46351 21001
rect 46293 20961 46305 20995
rect 46339 20992 46351 20995
rect 47762 20992 47768 21004
rect 46339 20964 47768 20992
rect 46339 20961 46351 20964
rect 46293 20955 46351 20961
rect 47762 20952 47768 20964
rect 47820 20952 47826 21004
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 22741 20927 22799 20933
rect 22741 20924 22753 20927
rect 22066 20896 22753 20924
rect 22741 20893 22753 20896
rect 22787 20893 22799 20927
rect 22741 20887 22799 20893
rect 23382 20884 23388 20936
rect 23440 20924 23446 20936
rect 23477 20927 23535 20933
rect 23477 20924 23489 20927
rect 23440 20896 23489 20924
rect 23440 20884 23446 20896
rect 23477 20893 23489 20896
rect 23523 20893 23535 20927
rect 23477 20887 23535 20893
rect 24397 20927 24455 20933
rect 24397 20893 24409 20927
rect 24443 20893 24455 20927
rect 26694 20924 26700 20936
rect 26655 20896 26700 20924
rect 24397 20887 24455 20893
rect 21913 20859 21971 20865
rect 21913 20856 21925 20859
rect 20272 20828 21925 20856
rect 21913 20825 21925 20828
rect 21959 20825 21971 20859
rect 21913 20819 21971 20825
rect 22186 20816 22192 20868
rect 22244 20856 22250 20868
rect 22281 20859 22339 20865
rect 22281 20856 22293 20859
rect 22244 20828 22293 20856
rect 22244 20816 22250 20828
rect 22281 20825 22293 20828
rect 22327 20856 22339 20859
rect 23400 20856 23428 20884
rect 22327 20828 23428 20856
rect 24412 20856 24440 20887
rect 26694 20884 26700 20896
rect 26752 20884 26758 20936
rect 27246 20884 27252 20936
rect 27304 20924 27310 20936
rect 27525 20927 27583 20933
rect 27525 20924 27537 20927
rect 27304 20896 27537 20924
rect 27304 20884 27310 20896
rect 27525 20893 27537 20896
rect 27571 20924 27583 20927
rect 29546 20924 29552 20936
rect 27571 20896 29552 20924
rect 27571 20893 27583 20896
rect 27525 20887 27583 20893
rect 29546 20884 29552 20896
rect 29604 20924 29610 20936
rect 30377 20927 30435 20933
rect 30377 20924 30389 20927
rect 29604 20896 30389 20924
rect 29604 20884 29610 20896
rect 30377 20893 30389 20896
rect 30423 20893 30435 20927
rect 30377 20887 30435 20893
rect 24581 20859 24639 20865
rect 24412 20828 24532 20856
rect 22327 20825 22339 20828
rect 22281 20819 22339 20825
rect 15105 20791 15163 20797
rect 15105 20788 15117 20791
rect 14292 20760 15117 20788
rect 15105 20757 15117 20760
rect 15151 20757 15163 20791
rect 15105 20751 15163 20757
rect 18598 20748 18604 20800
rect 18656 20788 18662 20800
rect 19429 20791 19487 20797
rect 19429 20788 19441 20791
rect 18656 20760 19441 20788
rect 18656 20748 18662 20760
rect 19429 20757 19441 20760
rect 19475 20757 19487 20791
rect 19429 20751 19487 20757
rect 21174 20748 21180 20800
rect 21232 20788 21238 20800
rect 21269 20791 21327 20797
rect 21269 20788 21281 20791
rect 21232 20760 21281 20788
rect 21232 20748 21238 20760
rect 21269 20757 21281 20760
rect 21315 20757 21327 20791
rect 21269 20751 21327 20757
rect 23569 20791 23627 20797
rect 23569 20757 23581 20791
rect 23615 20788 23627 20791
rect 24394 20788 24400 20800
rect 23615 20760 24400 20788
rect 23615 20757 23627 20760
rect 23569 20751 23627 20757
rect 24394 20748 24400 20760
rect 24452 20748 24458 20800
rect 24504 20788 24532 20828
rect 24581 20825 24593 20859
rect 24627 20856 24639 20859
rect 24762 20856 24768 20868
rect 24627 20828 24768 20856
rect 24627 20825 24639 20828
rect 24581 20819 24639 20825
rect 24762 20816 24768 20828
rect 24820 20816 24826 20868
rect 30558 20856 30564 20868
rect 30519 20828 30564 20856
rect 30558 20816 30564 20828
rect 30616 20816 30622 20868
rect 46474 20856 46480 20868
rect 46435 20828 46480 20856
rect 46474 20816 46480 20828
rect 46532 20816 46538 20868
rect 24854 20788 24860 20800
rect 24504 20760 24860 20788
rect 24854 20748 24860 20760
rect 24912 20788 24918 20800
rect 26142 20788 26148 20800
rect 24912 20760 26148 20788
rect 24912 20748 24918 20760
rect 26142 20748 26148 20760
rect 26200 20748 26206 20800
rect 26789 20791 26847 20797
rect 26789 20757 26801 20791
rect 26835 20788 26847 20791
rect 27798 20788 27804 20800
rect 26835 20760 27804 20788
rect 26835 20757 26847 20760
rect 26789 20751 26847 20757
rect 27798 20748 27804 20760
rect 27856 20748 27862 20800
rect 46290 20748 46296 20800
rect 46348 20788 46354 20800
rect 47302 20788 47308 20800
rect 46348 20760 47308 20788
rect 46348 20748 46354 20760
rect 47302 20748 47308 20760
rect 47360 20748 47366 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 10594 20584 10600 20596
rect 10060 20556 10600 20584
rect 10060 20457 10088 20556
rect 10594 20544 10600 20556
rect 10652 20584 10658 20596
rect 13078 20584 13084 20596
rect 10652 20556 13084 20584
rect 10652 20544 10658 20556
rect 13078 20544 13084 20556
rect 13136 20544 13142 20596
rect 21358 20544 21364 20596
rect 21416 20584 21422 20596
rect 29546 20584 29552 20596
rect 21416 20556 29408 20584
rect 29507 20556 29552 20584
rect 21416 20544 21422 20556
rect 14182 20516 14188 20528
rect 13570 20488 14188 20516
rect 14182 20476 14188 20488
rect 14240 20476 14246 20528
rect 21174 20516 21180 20528
rect 15948 20488 21180 20516
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 10229 20451 10287 20457
rect 10229 20417 10241 20451
rect 10275 20417 10287 20451
rect 10229 20411 10287 20417
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 10244 20380 10272 20411
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 14277 20451 14335 20457
rect 10376 20420 10421 20448
rect 10376 20408 10382 20420
rect 14277 20417 14289 20451
rect 14323 20417 14335 20451
rect 14277 20411 14335 20417
rect 10778 20380 10784 20392
rect 9732 20352 10784 20380
rect 9732 20340 9738 20352
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 11606 20340 11612 20392
rect 11664 20380 11670 20392
rect 12069 20383 12127 20389
rect 12069 20380 12081 20383
rect 11664 20352 12081 20380
rect 11664 20340 11670 20352
rect 12069 20349 12081 20352
rect 12115 20349 12127 20383
rect 12342 20380 12348 20392
rect 12303 20352 12348 20380
rect 12069 20343 12127 20349
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 14292 20380 14320 20411
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 15948 20457 15976 20488
rect 21174 20476 21180 20488
rect 21232 20476 21238 20528
rect 22094 20516 22100 20528
rect 21928 20488 22100 20516
rect 15933 20451 15991 20457
rect 15933 20448 15945 20451
rect 15896 20420 15945 20448
rect 15896 20408 15902 20420
rect 15933 20417 15945 20420
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20417 17463 20451
rect 17405 20411 17463 20417
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20448 18107 20451
rect 18414 20448 18420 20460
rect 18095 20420 18420 20448
rect 18095 20417 18107 20420
rect 18049 20411 18107 20417
rect 12492 20352 14320 20380
rect 17420 20380 17448 20411
rect 18414 20408 18420 20420
rect 18472 20408 18478 20460
rect 18598 20448 18604 20460
rect 18559 20420 18604 20448
rect 18598 20408 18604 20420
rect 18656 20408 18662 20460
rect 20162 20408 20168 20460
rect 20220 20448 20226 20460
rect 21928 20457 21956 20488
rect 22094 20476 22100 20488
rect 22152 20476 22158 20528
rect 24394 20516 24400 20528
rect 24355 20488 24400 20516
rect 24394 20476 24400 20488
rect 24452 20476 24458 20528
rect 28074 20516 28080 20528
rect 28035 20488 28080 20516
rect 28074 20476 28080 20488
rect 28132 20476 28138 20528
rect 28626 20476 28632 20528
rect 28684 20476 28690 20528
rect 29380 20516 29408 20556
rect 29546 20544 29552 20556
rect 29604 20544 29610 20596
rect 30558 20584 30564 20596
rect 30519 20556 30564 20584
rect 30558 20544 30564 20556
rect 30616 20544 30622 20596
rect 46382 20584 46388 20596
rect 35866 20556 46388 20584
rect 30098 20516 30104 20528
rect 29380 20488 30104 20516
rect 30098 20476 30104 20488
rect 30156 20476 30162 20528
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 20220 20420 20637 20448
rect 20220 20408 20226 20420
rect 20625 20417 20637 20420
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 21913 20451 21971 20457
rect 21913 20417 21925 20451
rect 21959 20417 21971 20451
rect 24210 20448 24216 20460
rect 24171 20420 24216 20448
rect 21913 20411 21971 20417
rect 24210 20408 24216 20420
rect 24268 20408 24274 20460
rect 26970 20448 26976 20460
rect 26931 20420 26976 20448
rect 26970 20408 26976 20420
rect 27028 20448 27034 20460
rect 27614 20448 27620 20460
rect 27028 20420 27620 20448
rect 27028 20408 27034 20420
rect 27614 20408 27620 20420
rect 27672 20408 27678 20460
rect 27798 20448 27804 20460
rect 27759 20420 27804 20448
rect 27798 20408 27804 20420
rect 27856 20408 27862 20460
rect 30466 20448 30472 20460
rect 30379 20420 30472 20448
rect 30466 20408 30472 20420
rect 30524 20448 30530 20460
rect 35866 20448 35894 20556
rect 46382 20544 46388 20556
rect 46440 20544 46446 20596
rect 46474 20544 46480 20596
rect 46532 20584 46538 20596
rect 46845 20587 46903 20593
rect 46845 20584 46857 20587
rect 46532 20556 46857 20584
rect 46532 20544 46538 20556
rect 46845 20553 46857 20556
rect 46891 20553 46903 20587
rect 46845 20547 46903 20553
rect 46290 20516 46296 20528
rect 45112 20488 46296 20516
rect 45112 20457 45140 20488
rect 45756 20457 45784 20488
rect 46290 20476 46296 20488
rect 46348 20476 46354 20528
rect 30524 20420 35894 20448
rect 45097 20451 45155 20457
rect 30524 20408 30530 20420
rect 45097 20417 45109 20451
rect 45143 20417 45155 20451
rect 45097 20411 45155 20417
rect 45281 20451 45339 20457
rect 45281 20417 45293 20451
rect 45327 20417 45339 20451
rect 45281 20411 45339 20417
rect 45741 20451 45799 20457
rect 45741 20417 45753 20451
rect 45787 20417 45799 20451
rect 45922 20448 45928 20460
rect 45883 20420 45928 20448
rect 45741 20411 45799 20417
rect 18506 20380 18512 20392
rect 17420 20352 18512 20380
rect 12492 20340 12498 20352
rect 18506 20340 18512 20352
rect 18564 20340 18570 20392
rect 21177 20383 21235 20389
rect 21177 20349 21189 20383
rect 21223 20380 21235 20383
rect 21358 20380 21364 20392
rect 21223 20352 21364 20380
rect 21223 20349 21235 20352
rect 21177 20343 21235 20349
rect 21358 20340 21364 20352
rect 21416 20340 21422 20392
rect 22097 20383 22155 20389
rect 22097 20349 22109 20383
rect 22143 20380 22155 20383
rect 22278 20380 22284 20392
rect 22143 20352 22284 20380
rect 22143 20349 22155 20352
rect 22097 20343 22155 20349
rect 22278 20340 22284 20352
rect 22336 20340 22342 20392
rect 22373 20383 22431 20389
rect 22373 20349 22385 20383
rect 22419 20349 22431 20383
rect 26050 20380 26056 20392
rect 26011 20352 26056 20380
rect 22373 20343 22431 20349
rect 13906 20272 13912 20324
rect 13964 20312 13970 20324
rect 22388 20312 22416 20343
rect 26050 20340 26056 20352
rect 26108 20340 26114 20392
rect 45296 20380 45324 20411
rect 45922 20408 45928 20420
rect 45980 20408 45986 20460
rect 46474 20408 46480 20460
rect 46532 20448 46538 20460
rect 46753 20451 46811 20457
rect 46753 20448 46765 20451
rect 46532 20420 46765 20448
rect 46532 20408 46538 20420
rect 46753 20417 46765 20420
rect 46799 20417 46811 20451
rect 47762 20448 47768 20460
rect 47723 20420 47768 20448
rect 46753 20411 46811 20417
rect 47762 20408 47768 20420
rect 47820 20408 47826 20460
rect 45940 20380 45968 20408
rect 45296 20352 45968 20380
rect 13964 20284 22416 20312
rect 13964 20272 13970 20284
rect 9861 20247 9919 20253
rect 9861 20213 9873 20247
rect 9907 20244 9919 20247
rect 9950 20244 9956 20256
rect 9907 20216 9956 20244
rect 9907 20213 9919 20216
rect 9861 20207 9919 20213
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 13817 20247 13875 20253
rect 13817 20213 13829 20247
rect 13863 20244 13875 20247
rect 14090 20244 14096 20256
rect 13863 20216 14096 20244
rect 13863 20213 13875 20216
rect 13817 20207 13875 20213
rect 14090 20204 14096 20216
rect 14148 20204 14154 20256
rect 14182 20204 14188 20256
rect 14240 20244 14246 20256
rect 14458 20244 14464 20256
rect 14240 20216 14464 20244
rect 14240 20204 14246 20216
rect 14458 20204 14464 20216
rect 14516 20204 14522 20256
rect 15930 20204 15936 20256
rect 15988 20244 15994 20256
rect 16025 20247 16083 20253
rect 16025 20244 16037 20247
rect 15988 20216 16037 20244
rect 15988 20204 15994 20216
rect 16025 20213 16037 20216
rect 16071 20213 16083 20247
rect 17218 20244 17224 20256
rect 17179 20216 17224 20244
rect 16025 20207 16083 20213
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 17494 20204 17500 20256
rect 17552 20244 17558 20256
rect 17865 20247 17923 20253
rect 17865 20244 17877 20247
rect 17552 20216 17877 20244
rect 17552 20204 17558 20216
rect 17865 20213 17877 20216
rect 17911 20213 17923 20247
rect 17865 20207 17923 20213
rect 18693 20247 18751 20253
rect 18693 20213 18705 20247
rect 18739 20244 18751 20247
rect 18782 20244 18788 20256
rect 18739 20216 18788 20244
rect 18739 20213 18751 20216
rect 18693 20207 18751 20213
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 23382 20204 23388 20256
rect 23440 20244 23446 20256
rect 25774 20244 25780 20256
rect 23440 20216 25780 20244
rect 23440 20204 23446 20216
rect 25774 20204 25780 20216
rect 25832 20204 25838 20256
rect 27062 20244 27068 20256
rect 27023 20216 27068 20244
rect 27062 20204 27068 20216
rect 27120 20204 27126 20256
rect 45186 20244 45192 20256
rect 45147 20216 45192 20244
rect 45186 20204 45192 20216
rect 45244 20204 45250 20256
rect 45738 20244 45744 20256
rect 45699 20216 45744 20244
rect 45738 20204 45744 20216
rect 45796 20204 45802 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 11606 20040 11612 20052
rect 11567 20012 11612 20040
rect 11606 20000 11612 20012
rect 11664 20000 11670 20052
rect 12161 20043 12219 20049
rect 12161 20009 12173 20043
rect 12207 20040 12219 20043
rect 12342 20040 12348 20052
rect 12207 20012 12348 20040
rect 12207 20009 12219 20012
rect 12161 20003 12219 20009
rect 12342 20000 12348 20012
rect 12400 20000 12406 20052
rect 14645 20043 14703 20049
rect 14645 20009 14657 20043
rect 14691 20040 14703 20043
rect 14918 20040 14924 20052
rect 14691 20012 14924 20040
rect 14691 20009 14703 20012
rect 14645 20003 14703 20009
rect 14918 20000 14924 20012
rect 14976 20000 14982 20052
rect 26142 20040 26148 20052
rect 17604 20012 22094 20040
rect 9950 19972 9956 19984
rect 9911 19944 9956 19972
rect 9950 19932 9956 19944
rect 10008 19932 10014 19984
rect 13906 19972 13912 19984
rect 10060 19944 13912 19972
rect 3970 19864 3976 19916
rect 4028 19904 4034 19916
rect 10060 19904 10088 19944
rect 13906 19932 13912 19944
rect 13964 19932 13970 19984
rect 14090 19972 14096 19984
rect 14051 19944 14096 19972
rect 14090 19932 14096 19944
rect 14148 19932 14154 19984
rect 4028 19876 10088 19904
rect 4028 19864 4034 19876
rect 10318 19864 10324 19916
rect 10376 19904 10382 19916
rect 13998 19904 14004 19916
rect 10376 19876 12204 19904
rect 10376 19864 10382 19876
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 9677 19839 9735 19845
rect 9677 19805 9689 19839
rect 9723 19836 9735 19839
rect 10226 19836 10232 19848
rect 9723 19808 10232 19836
rect 9723 19805 9735 19808
rect 9677 19799 9735 19805
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 10594 19796 10600 19848
rect 10652 19836 10658 19848
rect 11425 19839 11483 19845
rect 10652 19830 11376 19836
rect 11425 19830 11437 19839
rect 10652 19808 11437 19830
rect 10652 19796 10658 19808
rect 11348 19805 11437 19808
rect 11471 19805 11483 19839
rect 11348 19802 11483 19805
rect 12176 19830 12204 19876
rect 12636 19876 14004 19904
rect 12636 19845 12664 19876
rect 13998 19864 14004 19876
rect 14056 19864 14062 19916
rect 12345 19839 12403 19845
rect 12345 19836 12357 19839
rect 12268 19830 12357 19836
rect 12176 19808 12357 19830
rect 12176 19802 12296 19808
rect 12345 19805 12357 19808
rect 12391 19805 12403 19839
rect 11425 19799 11483 19802
rect 12345 19799 12403 19805
rect 12621 19839 12679 19845
rect 12621 19805 12633 19839
rect 12667 19805 12679 19839
rect 12621 19799 12679 19805
rect 12805 19839 12863 19845
rect 12805 19805 12817 19839
rect 12851 19836 12863 19839
rect 14108 19836 14136 19932
rect 15930 19904 15936 19916
rect 15891 19876 15936 19904
rect 15930 19864 15936 19876
rect 15988 19864 15994 19916
rect 17604 19913 17632 20012
rect 18414 19932 18420 19984
rect 18472 19972 18478 19984
rect 19889 19975 19947 19981
rect 19889 19972 19901 19975
rect 18472 19944 19901 19972
rect 18472 19932 18478 19944
rect 19889 19941 19901 19944
rect 19935 19972 19947 19975
rect 20254 19972 20260 19984
rect 19935 19944 20260 19972
rect 19935 19941 19947 19944
rect 19889 19935 19947 19941
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 17589 19907 17647 19913
rect 17589 19873 17601 19907
rect 17635 19873 17647 19907
rect 18322 19904 18328 19916
rect 18283 19876 18328 19904
rect 17589 19867 17647 19873
rect 18322 19864 18328 19876
rect 18380 19864 18386 19916
rect 22066 19904 22094 20012
rect 23216 20012 25728 20040
rect 26103 20012 26148 20040
rect 23216 19904 23244 20012
rect 23382 19904 23388 19916
rect 18432 19876 21864 19904
rect 22066 19876 23244 19904
rect 23343 19876 23388 19904
rect 18432 19848 18460 19876
rect 21836 19848 21864 19876
rect 23382 19864 23388 19876
rect 23440 19864 23446 19916
rect 24673 19907 24731 19913
rect 24673 19873 24685 19907
rect 24719 19904 24731 19907
rect 25314 19904 25320 19916
rect 24719 19876 25320 19904
rect 24719 19873 24731 19876
rect 24673 19867 24731 19873
rect 25314 19864 25320 19876
rect 25372 19864 25378 19916
rect 25700 19904 25728 20012
rect 26142 20000 26148 20012
rect 26200 20000 26206 20052
rect 27522 20040 27528 20052
rect 27483 20012 27528 20040
rect 27522 20000 27528 20012
rect 27580 20000 27586 20052
rect 28626 20040 28632 20052
rect 28587 20012 28632 20040
rect 28626 20000 28632 20012
rect 28684 20000 28690 20052
rect 46198 20040 46204 20052
rect 35866 20012 46204 20040
rect 25774 19932 25780 19984
rect 25832 19972 25838 19984
rect 30466 19972 30472 19984
rect 25832 19944 30472 19972
rect 25832 19932 25838 19944
rect 30466 19932 30472 19944
rect 30524 19932 30530 19984
rect 35866 19904 35894 20012
rect 46198 20000 46204 20012
rect 46256 20000 46262 20052
rect 45186 19932 45192 19984
rect 45244 19972 45250 19984
rect 45649 19975 45707 19981
rect 45649 19972 45661 19975
rect 45244 19944 45661 19972
rect 45244 19932 45250 19944
rect 45649 19941 45661 19944
rect 45695 19941 45707 19975
rect 45649 19935 45707 19941
rect 25700 19876 35894 19904
rect 45373 19907 45431 19913
rect 45373 19873 45385 19907
rect 45419 19904 45431 19907
rect 45554 19904 45560 19916
rect 45419 19876 45560 19904
rect 45419 19873 45431 19876
rect 45373 19867 45431 19873
rect 45554 19864 45560 19876
rect 45612 19904 45618 19916
rect 45738 19904 45744 19916
rect 45612 19876 45744 19904
rect 45612 19864 45618 19876
rect 45738 19864 45744 19876
rect 45796 19864 45802 19916
rect 46293 19907 46351 19913
rect 46293 19873 46305 19907
rect 46339 19904 46351 19907
rect 47026 19904 47032 19916
rect 46339 19876 47032 19904
rect 46339 19873 46351 19876
rect 46293 19867 46351 19873
rect 47026 19864 47032 19876
rect 47084 19864 47090 19916
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 12851 19808 14136 19836
rect 14292 19808 15761 19836
rect 12851 19805 12863 19808
rect 12805 19799 12863 19805
rect 9122 19728 9128 19780
rect 9180 19768 9186 19780
rect 11440 19768 11468 19799
rect 12066 19768 12072 19780
rect 9180 19740 10916 19768
rect 11440 19740 12072 19768
rect 9180 19728 9186 19740
rect 10137 19703 10195 19709
rect 10137 19669 10149 19703
rect 10183 19700 10195 19703
rect 10778 19700 10784 19712
rect 10183 19672 10784 19700
rect 10183 19669 10195 19672
rect 10137 19663 10195 19669
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 10888 19700 10916 19740
rect 12066 19728 12072 19740
rect 12124 19728 12130 19780
rect 12820 19768 12848 19799
rect 12406 19740 12848 19768
rect 12406 19700 12434 19740
rect 10888 19672 12434 19700
rect 13446 19660 13452 19712
rect 13504 19700 13510 19712
rect 14292 19709 14320 19808
rect 15749 19805 15761 19808
rect 15795 19805 15807 19839
rect 18230 19836 18236 19848
rect 18191 19808 18236 19836
rect 15749 19799 15807 19805
rect 18230 19796 18236 19808
rect 18288 19796 18294 19848
rect 18414 19836 18420 19848
rect 18375 19808 18420 19836
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 18509 19839 18567 19845
rect 18509 19805 18521 19839
rect 18555 19805 18567 19839
rect 18509 19799 18567 19805
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19836 19763 19839
rect 19978 19836 19984 19848
rect 19751 19808 19984 19836
rect 19751 19805 19763 19808
rect 19705 19799 19763 19805
rect 14369 19771 14427 19777
rect 14369 19737 14381 19771
rect 14415 19768 14427 19771
rect 14734 19768 14740 19780
rect 14415 19740 14740 19768
rect 14415 19737 14427 19740
rect 14369 19731 14427 19737
rect 14734 19728 14740 19740
rect 14792 19728 14798 19780
rect 17126 19728 17132 19780
rect 17184 19768 17190 19780
rect 17184 19740 18276 19768
rect 17184 19728 17190 19740
rect 18248 19739 18276 19740
rect 18524 19739 18552 19799
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 20438 19836 20444 19848
rect 20399 19808 20444 19836
rect 20438 19796 20444 19808
rect 20496 19796 20502 19848
rect 21174 19836 21180 19848
rect 21135 19808 21180 19836
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21818 19836 21824 19848
rect 21731 19808 21824 19836
rect 21818 19796 21824 19808
rect 21876 19796 21882 19848
rect 24394 19836 24400 19848
rect 24355 19808 24400 19836
rect 24394 19796 24400 19808
rect 24452 19796 24458 19848
rect 27062 19836 27068 19848
rect 25806 19808 27068 19836
rect 27062 19796 27068 19808
rect 27120 19796 27126 19848
rect 27246 19836 27252 19848
rect 27207 19808 27252 19836
rect 27246 19796 27252 19808
rect 27304 19796 27310 19848
rect 27338 19796 27344 19848
rect 27396 19796 27402 19848
rect 27614 19796 27620 19848
rect 27672 19836 27678 19848
rect 28537 19839 28595 19845
rect 28537 19836 28549 19839
rect 27672 19808 28549 19836
rect 27672 19796 27678 19808
rect 28537 19805 28549 19808
rect 28583 19805 28595 19839
rect 28537 19799 28595 19805
rect 14277 19703 14335 19709
rect 14277 19700 14289 19703
rect 13504 19672 14289 19700
rect 13504 19660 13510 19672
rect 14277 19669 14289 19672
rect 14323 19669 14335 19703
rect 14277 19663 14335 19669
rect 14461 19703 14519 19709
rect 14461 19669 14473 19703
rect 14507 19700 14519 19703
rect 14550 19700 14556 19712
rect 14507 19672 14556 19700
rect 14507 19669 14519 19672
rect 14461 19663 14519 19669
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 18046 19700 18052 19712
rect 18007 19672 18052 19700
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 18248 19711 18552 19739
rect 21269 19771 21327 19777
rect 21269 19737 21281 19771
rect 21315 19768 21327 19771
rect 22005 19771 22063 19777
rect 22005 19768 22017 19771
rect 21315 19740 22017 19768
rect 21315 19737 21327 19740
rect 21269 19731 21327 19737
rect 22005 19737 22017 19740
rect 22051 19737 22063 19771
rect 22005 19731 22063 19737
rect 22370 19728 22376 19780
rect 22428 19768 22434 19780
rect 22646 19768 22652 19780
rect 22428 19740 22652 19768
rect 22428 19728 22434 19740
rect 22646 19728 22652 19740
rect 22704 19728 22710 19780
rect 26878 19728 26884 19780
rect 26936 19768 26942 19780
rect 26973 19771 27031 19777
rect 26973 19768 26985 19771
rect 26936 19740 26985 19768
rect 26936 19728 26942 19740
rect 26973 19737 26985 19740
rect 27019 19737 27031 19771
rect 26973 19731 27031 19737
rect 27157 19771 27215 19777
rect 27157 19737 27169 19771
rect 27203 19768 27215 19771
rect 27356 19768 27384 19796
rect 27203 19740 27384 19768
rect 46477 19771 46535 19777
rect 27203 19737 27215 19740
rect 27157 19731 27215 19737
rect 46477 19737 46489 19771
rect 46523 19768 46535 19771
rect 47670 19768 47676 19780
rect 46523 19740 47676 19768
rect 46523 19737 46535 19740
rect 46477 19731 46535 19737
rect 47670 19728 47676 19740
rect 47728 19728 47734 19780
rect 48130 19768 48136 19780
rect 48091 19740 48136 19768
rect 48130 19728 48136 19740
rect 48188 19728 48194 19780
rect 18524 19700 18552 19711
rect 19242 19700 19248 19712
rect 18524 19672 19248 19700
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 19978 19660 19984 19712
rect 20036 19700 20042 19712
rect 20625 19703 20683 19709
rect 20625 19700 20637 19703
rect 20036 19672 20637 19700
rect 20036 19660 20042 19672
rect 20625 19669 20637 19672
rect 20671 19669 20683 19703
rect 20625 19663 20683 19669
rect 27341 19703 27399 19709
rect 27341 19669 27353 19703
rect 27387 19700 27399 19703
rect 27430 19700 27436 19712
rect 27387 19672 27436 19700
rect 27387 19669 27399 19672
rect 27341 19663 27399 19669
rect 27430 19660 27436 19672
rect 27488 19660 27494 19712
rect 45833 19703 45891 19709
rect 45833 19669 45845 19703
rect 45879 19700 45891 19703
rect 46290 19700 46296 19712
rect 45879 19672 46296 19700
rect 45879 19669 45891 19672
rect 45833 19663 45891 19669
rect 46290 19660 46296 19672
rect 46348 19660 46354 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 10597 19499 10655 19505
rect 10597 19465 10609 19499
rect 10643 19496 10655 19499
rect 11606 19496 11612 19508
rect 10643 19468 11612 19496
rect 10643 19465 10655 19468
rect 10597 19459 10655 19465
rect 11606 19456 11612 19468
rect 11664 19456 11670 19508
rect 11716 19468 11928 19496
rect 3510 19388 3516 19440
rect 3568 19428 3574 19440
rect 11716 19428 11744 19468
rect 3568 19400 11744 19428
rect 11900 19428 11928 19468
rect 12066 19456 12072 19508
rect 12124 19496 12130 19508
rect 12161 19499 12219 19505
rect 12161 19496 12173 19499
rect 12124 19468 12173 19496
rect 12124 19456 12130 19468
rect 12161 19465 12173 19468
rect 12207 19465 12219 19499
rect 22278 19496 22284 19508
rect 12161 19459 12219 19465
rect 12406 19468 22094 19496
rect 22239 19468 22284 19496
rect 12406 19428 12434 19468
rect 11900 19400 12434 19428
rect 13633 19431 13691 19437
rect 3568 19388 3574 19400
rect 13633 19397 13645 19431
rect 13679 19428 13691 19431
rect 14734 19428 14740 19440
rect 13679 19400 14740 19428
rect 13679 19397 13691 19400
rect 13633 19391 13691 19397
rect 14734 19388 14740 19400
rect 14792 19388 14798 19440
rect 17218 19388 17224 19440
rect 17276 19428 17282 19440
rect 17773 19431 17831 19437
rect 17773 19428 17785 19431
rect 17276 19400 17785 19428
rect 17276 19388 17282 19400
rect 17773 19397 17785 19400
rect 17819 19397 17831 19431
rect 17773 19391 17831 19397
rect 18782 19388 18788 19440
rect 18840 19388 18846 19440
rect 22066 19428 22094 19468
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 26878 19496 26884 19508
rect 22848 19468 26884 19496
rect 22066 19400 22324 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 9033 19363 9091 19369
rect 9033 19329 9045 19363
rect 9079 19360 9091 19363
rect 9674 19360 9680 19372
rect 9079 19332 9680 19360
rect 9079 19329 9091 19332
rect 9033 19323 9091 19329
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 9858 19360 9864 19372
rect 9819 19332 9864 19360
rect 9858 19320 9864 19332
rect 9916 19360 9922 19372
rect 10594 19360 10600 19372
rect 9916 19332 10600 19360
rect 9916 19320 9922 19332
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 10778 19360 10784 19372
rect 10739 19332 10784 19360
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 11974 19360 11980 19372
rect 11935 19332 11980 19360
rect 11974 19320 11980 19332
rect 12032 19320 12038 19372
rect 12066 19320 12072 19372
rect 12124 19360 12130 19372
rect 12434 19360 12440 19372
rect 12124 19332 12440 19360
rect 12124 19320 12130 19332
rect 12434 19320 12440 19332
rect 12492 19360 12498 19372
rect 12713 19363 12771 19369
rect 12713 19360 12725 19363
rect 12492 19332 12725 19360
rect 12492 19320 12498 19332
rect 12713 19329 12725 19332
rect 12759 19329 12771 19363
rect 12713 19323 12771 19329
rect 13725 19363 13783 19369
rect 13725 19329 13737 19363
rect 13771 19329 13783 19363
rect 13725 19323 13783 19329
rect 13817 19363 13875 19369
rect 13817 19329 13829 19363
rect 13863 19360 13875 19363
rect 14274 19360 14280 19372
rect 13863 19332 14280 19360
rect 13863 19329 13875 19332
rect 13817 19323 13875 19329
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19292 9183 19295
rect 10318 19292 10324 19304
rect 9171 19264 10324 19292
rect 9171 19261 9183 19264
rect 9125 19255 9183 19261
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 13446 19224 13452 19236
rect 13407 19196 13452 19224
rect 13446 19184 13452 19196
rect 13504 19184 13510 19236
rect 13740 19224 13768 19323
rect 14274 19320 14280 19332
rect 14332 19320 14338 19372
rect 17494 19360 17500 19372
rect 17455 19332 17500 19360
rect 17494 19320 17500 19332
rect 17552 19320 17558 19372
rect 20530 19360 20536 19372
rect 20491 19332 20536 19360
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 22186 19360 22192 19372
rect 22147 19332 22192 19360
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22296 19360 22324 19400
rect 22848 19369 22876 19468
rect 26878 19456 26884 19468
rect 26936 19456 26942 19508
rect 27246 19456 27252 19508
rect 27304 19496 27310 19508
rect 27617 19499 27675 19505
rect 27617 19496 27629 19499
rect 27304 19468 27629 19496
rect 27304 19456 27310 19468
rect 27617 19465 27629 19468
rect 27663 19465 27675 19499
rect 27617 19459 27675 19465
rect 45186 19388 45192 19440
rect 45244 19428 45250 19440
rect 47673 19431 47731 19437
rect 47673 19428 47685 19431
rect 45244 19400 46244 19428
rect 45244 19388 45250 19400
rect 22833 19363 22891 19369
rect 22296 19332 22784 19360
rect 13998 19292 14004 19304
rect 13959 19264 14004 19292
rect 13998 19252 14004 19264
rect 14056 19252 14062 19304
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 18414 19292 18420 19304
rect 17276 19264 18420 19292
rect 17276 19252 17282 19264
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 22278 19252 22284 19304
rect 22336 19292 22342 19304
rect 22554 19292 22560 19304
rect 22336 19264 22560 19292
rect 22336 19252 22342 19264
rect 22554 19252 22560 19264
rect 22612 19252 22618 19304
rect 13906 19224 13912 19236
rect 13740 19196 13912 19224
rect 13906 19184 13912 19196
rect 13964 19224 13970 19236
rect 14550 19224 14556 19236
rect 13964 19196 14556 19224
rect 13964 19184 13970 19196
rect 14550 19184 14556 19196
rect 14608 19184 14614 19236
rect 16850 19184 16856 19236
rect 16908 19224 16914 19236
rect 17310 19224 17316 19236
rect 16908 19196 17316 19224
rect 16908 19184 16914 19196
rect 17310 19184 17316 19196
rect 17368 19184 17374 19236
rect 22756 19224 22784 19332
rect 22833 19329 22845 19363
rect 22879 19329 22891 19363
rect 22833 19323 22891 19329
rect 27338 19320 27344 19372
rect 27396 19360 27402 19372
rect 27433 19363 27491 19369
rect 27433 19360 27445 19363
rect 27396 19332 27445 19360
rect 27396 19320 27402 19332
rect 27433 19329 27445 19332
rect 27479 19329 27491 19363
rect 27433 19323 27491 19329
rect 27522 19320 27528 19372
rect 27580 19360 27586 19372
rect 27709 19363 27767 19369
rect 27709 19360 27721 19363
rect 27580 19332 27721 19360
rect 27580 19320 27586 19332
rect 27709 19329 27721 19332
rect 27755 19329 27767 19363
rect 45554 19360 45560 19372
rect 45515 19332 45560 19360
rect 27709 19323 27767 19329
rect 45554 19320 45560 19332
rect 45612 19320 45618 19372
rect 45738 19360 45744 19372
rect 45699 19332 45744 19360
rect 45738 19320 45744 19332
rect 45796 19320 45802 19372
rect 46216 19369 46244 19400
rect 46308 19400 47685 19428
rect 46201 19363 46259 19369
rect 46201 19329 46213 19363
rect 46247 19329 46259 19363
rect 46201 19323 46259 19329
rect 23014 19292 23020 19304
rect 22975 19264 23020 19292
rect 23014 19252 23020 19264
rect 23072 19252 23078 19304
rect 23293 19295 23351 19301
rect 23293 19261 23305 19295
rect 23339 19261 23351 19295
rect 23293 19255 23351 19261
rect 23308 19224 23336 19255
rect 18800 19196 22094 19224
rect 22756 19196 23336 19224
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 9401 19159 9459 19165
rect 9401 19156 9413 19159
rect 9364 19128 9413 19156
rect 9364 19116 9370 19128
rect 9401 19125 9413 19128
rect 9447 19125 9459 19159
rect 9401 19119 9459 19125
rect 10045 19159 10103 19165
rect 10045 19125 10057 19159
rect 10091 19156 10103 19159
rect 11330 19156 11336 19168
rect 10091 19128 11336 19156
rect 10091 19125 10103 19128
rect 10045 19119 10103 19125
rect 11330 19116 11336 19128
rect 11388 19116 11394 19168
rect 12894 19156 12900 19168
rect 12855 19128 12900 19156
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 18800 19156 18828 19196
rect 19242 19156 19248 19168
rect 13044 19128 18828 19156
rect 19203 19128 19248 19156
rect 13044 19116 13050 19128
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 20349 19159 20407 19165
rect 20349 19125 20361 19159
rect 20395 19156 20407 19159
rect 20806 19156 20812 19168
rect 20395 19128 20812 19156
rect 20395 19125 20407 19128
rect 20349 19119 20407 19125
rect 20806 19116 20812 19128
rect 20864 19116 20870 19168
rect 22066 19156 22094 19196
rect 46106 19184 46112 19236
rect 46164 19224 46170 19236
rect 46201 19227 46259 19233
rect 46201 19224 46213 19227
rect 46164 19196 46213 19224
rect 46164 19184 46170 19196
rect 46201 19193 46213 19196
rect 46247 19193 46259 19227
rect 46308 19224 46336 19400
rect 47673 19397 47685 19400
rect 47719 19397 47731 19431
rect 47673 19391 47731 19397
rect 46382 19320 46388 19372
rect 46440 19360 46446 19372
rect 47581 19363 47639 19369
rect 47581 19360 47593 19363
rect 46440 19332 47593 19360
rect 46440 19320 46446 19332
rect 47581 19329 47593 19332
rect 47627 19329 47639 19363
rect 47581 19323 47639 19329
rect 46382 19224 46388 19236
rect 46308 19196 46388 19224
rect 46201 19187 46259 19193
rect 46382 19184 46388 19196
rect 46440 19184 46446 19236
rect 22830 19156 22836 19168
rect 22066 19128 22836 19156
rect 22830 19116 22836 19128
rect 22888 19116 22894 19168
rect 27433 19159 27491 19165
rect 27433 19125 27445 19159
rect 27479 19156 27491 19159
rect 28166 19156 28172 19168
rect 27479 19128 28172 19156
rect 27479 19125 27491 19128
rect 27433 19119 27491 19125
rect 28166 19116 28172 19128
rect 28224 19116 28230 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 2225 18915 2283 18921
rect 3970 18912 3976 18964
rect 4028 18952 4034 18964
rect 4028 18924 17264 18952
rect 4028 18912 4034 18924
rect 9306 18816 9312 18828
rect 9267 18788 9312 18816
rect 9306 18776 9312 18788
rect 9364 18776 9370 18828
rect 9398 18776 9404 18828
rect 9456 18816 9462 18828
rect 11330 18816 11336 18828
rect 9456 18788 10916 18816
rect 11291 18788 11336 18816
rect 9456 18776 9462 18788
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18748 2194 18760
rect 9030 18748 9036 18760
rect 2188 18720 2774 18748
rect 8991 18720 9036 18748
rect 2188 18708 2194 18720
rect 2746 18680 2774 18720
rect 9030 18708 9036 18720
rect 9088 18708 9094 18760
rect 6638 18680 6644 18692
rect 2746 18652 6644 18680
rect 6638 18640 6644 18652
rect 6696 18680 6702 18692
rect 9398 18680 9404 18692
rect 6696 18652 9404 18680
rect 6696 18640 6702 18652
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 10318 18640 10324 18692
rect 10376 18640 10382 18692
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 10781 18615 10839 18621
rect 10781 18612 10793 18615
rect 9732 18584 10793 18612
rect 9732 18572 9738 18584
rect 10781 18581 10793 18584
rect 10827 18581 10839 18615
rect 10888 18612 10916 18788
rect 11330 18776 11336 18788
rect 11388 18776 11394 18828
rect 11606 18816 11612 18828
rect 11567 18788 11612 18816
rect 11606 18776 11612 18788
rect 11664 18776 11670 18828
rect 12894 18776 12900 18828
rect 12952 18816 12958 18828
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 12952 18788 14105 18816
rect 12952 18776 12958 18788
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 17126 18816 17132 18828
rect 17087 18788 17132 18816
rect 14093 18779 14151 18785
rect 17126 18776 17132 18788
rect 17184 18776 17190 18828
rect 17236 18816 17264 18924
rect 18506 18912 18512 18964
rect 18564 18952 18570 18964
rect 18601 18955 18659 18961
rect 18601 18952 18613 18955
rect 18564 18924 18613 18952
rect 18564 18912 18570 18924
rect 18601 18921 18613 18924
rect 18647 18921 18659 18955
rect 18601 18915 18659 18921
rect 19705 18955 19763 18961
rect 19705 18921 19717 18955
rect 19751 18952 19763 18955
rect 20530 18952 20536 18964
rect 19751 18924 20536 18952
rect 19751 18921 19763 18924
rect 19705 18915 19763 18921
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 21818 18912 21824 18964
rect 21876 18952 21882 18964
rect 22281 18955 22339 18961
rect 22281 18952 22293 18955
rect 21876 18924 22293 18952
rect 21876 18912 21882 18924
rect 22281 18921 22293 18924
rect 22327 18921 22339 18955
rect 22281 18915 22339 18921
rect 22925 18955 22983 18961
rect 22925 18921 22937 18955
rect 22971 18952 22983 18955
rect 23014 18952 23020 18964
rect 22971 18924 23020 18952
rect 22971 18921 22983 18924
rect 22925 18915 22983 18921
rect 23014 18912 23020 18924
rect 23072 18912 23078 18964
rect 24394 18952 24400 18964
rect 24355 18924 24400 18952
rect 24394 18912 24400 18924
rect 24452 18912 24458 18964
rect 27246 18912 27252 18964
rect 27304 18952 27310 18964
rect 27525 18955 27583 18961
rect 27525 18952 27537 18955
rect 27304 18924 27537 18952
rect 27304 18912 27310 18924
rect 27525 18921 27537 18924
rect 27571 18921 27583 18955
rect 27525 18915 27583 18921
rect 18046 18844 18052 18896
rect 18104 18884 18110 18896
rect 18417 18887 18475 18893
rect 18417 18884 18429 18887
rect 18104 18856 18429 18884
rect 18104 18844 18110 18856
rect 18417 18853 18429 18856
rect 18463 18853 18475 18887
rect 47394 18884 47400 18896
rect 18417 18847 18475 18853
rect 23676 18856 47400 18884
rect 17236 18788 23520 18816
rect 16666 18748 16672 18760
rect 16627 18720 16672 18748
rect 16666 18708 16672 18720
rect 16724 18708 16730 18760
rect 17402 18708 17408 18760
rect 17460 18748 17466 18760
rect 17681 18751 17739 18757
rect 17681 18748 17693 18751
rect 17460 18720 17693 18748
rect 17460 18708 17466 18720
rect 17681 18717 17693 18720
rect 17727 18748 17739 18751
rect 18141 18751 18199 18757
rect 18141 18748 18153 18751
rect 17727 18720 18153 18748
rect 17727 18717 17739 18720
rect 17681 18711 17739 18717
rect 18141 18717 18153 18720
rect 18187 18717 18199 18751
rect 19334 18748 19340 18760
rect 19295 18720 19340 18748
rect 18141 18711 18199 18717
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 19426 18708 19432 18760
rect 19484 18748 19490 18760
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 19484 18720 19533 18748
rect 19484 18708 19490 18720
rect 19521 18717 19533 18720
rect 19567 18717 19579 18751
rect 20530 18748 20536 18760
rect 20491 18720 20536 18748
rect 19521 18711 19579 18717
rect 20530 18708 20536 18720
rect 20588 18708 20594 18760
rect 22186 18708 22192 18760
rect 22244 18748 22250 18760
rect 22833 18751 22891 18757
rect 22833 18748 22845 18751
rect 22244 18720 22845 18748
rect 22244 18708 22250 18720
rect 22833 18717 22845 18720
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 12066 18640 12072 18692
rect 12124 18640 12130 18692
rect 13630 18640 13636 18692
rect 13688 18680 13694 18692
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 13688 18652 14381 18680
rect 13688 18640 13694 18652
rect 14369 18649 14381 18652
rect 14415 18649 14427 18683
rect 14369 18643 14427 18649
rect 14826 18640 14832 18692
rect 14884 18640 14890 18692
rect 16574 18640 16580 18692
rect 16632 18680 16638 18692
rect 17218 18680 17224 18692
rect 16632 18652 17224 18680
rect 16632 18640 16638 18652
rect 17218 18640 17224 18652
rect 17276 18680 17282 18692
rect 17313 18683 17371 18689
rect 17313 18680 17325 18683
rect 17276 18652 17325 18680
rect 17276 18640 17282 18652
rect 17313 18649 17325 18652
rect 17359 18649 17371 18683
rect 18414 18680 18420 18692
rect 17313 18643 17371 18649
rect 17420 18652 18420 18680
rect 12986 18612 12992 18624
rect 10888 18584 12992 18612
rect 10781 18575 10839 18581
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 13078 18572 13084 18624
rect 13136 18612 13142 18624
rect 13136 18584 13181 18612
rect 13136 18572 13142 18584
rect 13446 18572 13452 18624
rect 13504 18612 13510 18624
rect 17420 18621 17448 18652
rect 18414 18640 18420 18652
rect 18472 18640 18478 18692
rect 20070 18640 20076 18692
rect 20128 18680 20134 18692
rect 20809 18683 20867 18689
rect 20809 18680 20821 18683
rect 20128 18652 20821 18680
rect 20128 18640 20134 18652
rect 20809 18649 20821 18652
rect 20855 18649 20867 18683
rect 22646 18680 22652 18692
rect 22034 18652 22652 18680
rect 20809 18643 20867 18649
rect 22646 18640 22652 18652
rect 22704 18640 22710 18692
rect 23492 18680 23520 18788
rect 23676 18757 23704 18856
rect 47394 18844 47400 18856
rect 47452 18844 47458 18896
rect 25317 18819 25375 18825
rect 25317 18785 25329 18819
rect 25363 18785 25375 18819
rect 25317 18779 25375 18785
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18717 23719 18751
rect 24394 18748 24400 18760
rect 24355 18720 24400 18748
rect 23661 18711 23719 18717
rect 24394 18708 24400 18720
rect 24452 18708 24458 18760
rect 24854 18680 24860 18692
rect 23492 18652 24860 18680
rect 24854 18640 24860 18652
rect 24912 18640 24918 18692
rect 25332 18680 25360 18779
rect 25590 18776 25596 18828
rect 25648 18816 25654 18828
rect 25777 18819 25835 18825
rect 25777 18816 25789 18819
rect 25648 18788 25789 18816
rect 25648 18776 25654 18788
rect 25777 18785 25789 18788
rect 25823 18785 25835 18819
rect 26878 18816 26884 18828
rect 25777 18779 25835 18785
rect 25884 18788 26884 18816
rect 25409 18751 25467 18757
rect 25409 18717 25421 18751
rect 25455 18748 25467 18751
rect 25884 18748 25912 18788
rect 26878 18776 26884 18788
rect 26936 18776 26942 18828
rect 47302 18776 47308 18828
rect 47360 18816 47366 18828
rect 47489 18819 47547 18825
rect 47489 18816 47501 18819
rect 47360 18788 47501 18816
rect 47360 18776 47366 18788
rect 47489 18785 47501 18788
rect 47535 18785 47547 18819
rect 47489 18779 47547 18785
rect 25455 18720 25912 18748
rect 26237 18751 26295 18757
rect 25455 18717 25467 18720
rect 25409 18711 25467 18717
rect 26237 18717 26249 18751
rect 26283 18748 26295 18751
rect 26970 18748 26976 18760
rect 26283 18720 26976 18748
rect 26283 18717 26295 18720
rect 26237 18711 26295 18717
rect 26970 18708 26976 18720
rect 27028 18708 27034 18760
rect 28166 18748 28172 18760
rect 27264 18720 27568 18748
rect 28127 18720 28172 18748
rect 27264 18680 27292 18720
rect 25332 18652 27292 18680
rect 27338 18640 27344 18692
rect 27396 18680 27402 18692
rect 27540 18680 27568 18720
rect 28166 18708 28172 18720
rect 28224 18708 28230 18760
rect 28353 18751 28411 18757
rect 28353 18717 28365 18751
rect 28399 18717 28411 18751
rect 28353 18711 28411 18717
rect 28368 18680 28396 18711
rect 45738 18708 45744 18760
rect 45796 18748 45802 18760
rect 45925 18751 45983 18757
rect 45925 18748 45937 18751
rect 45796 18720 45937 18748
rect 45796 18708 45802 18720
rect 45925 18717 45937 18720
rect 45971 18717 45983 18751
rect 46290 18748 46296 18760
rect 46251 18720 46296 18748
rect 45925 18711 45983 18717
rect 46290 18708 46296 18720
rect 46348 18708 46354 18760
rect 27396 18652 27441 18680
rect 27540 18652 28396 18680
rect 27396 18640 27402 18652
rect 15841 18615 15899 18621
rect 15841 18612 15853 18615
rect 13504 18584 15853 18612
rect 13504 18572 13510 18584
rect 15841 18581 15853 18584
rect 15887 18581 15899 18615
rect 15841 18575 15899 18581
rect 16485 18615 16543 18621
rect 16485 18581 16497 18615
rect 16531 18612 16543 18615
rect 17405 18615 17463 18621
rect 17405 18612 17417 18615
rect 16531 18584 17417 18612
rect 16531 18581 16543 18584
rect 16485 18575 16543 18581
rect 17405 18581 17417 18584
rect 17451 18581 17463 18615
rect 17405 18575 17463 18581
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 23753 18615 23811 18621
rect 17552 18584 17597 18612
rect 17552 18572 17558 18584
rect 23753 18581 23765 18615
rect 23799 18612 23811 18615
rect 24210 18612 24216 18624
rect 23799 18584 24216 18612
rect 23799 18581 23811 18584
rect 23753 18575 23811 18581
rect 24210 18572 24216 18584
rect 24268 18572 24274 18624
rect 26234 18572 26240 18624
rect 26292 18612 26298 18624
rect 26329 18615 26387 18621
rect 26329 18612 26341 18615
rect 26292 18584 26341 18612
rect 26292 18572 26298 18584
rect 26329 18581 26341 18584
rect 26375 18581 26387 18615
rect 26329 18575 26387 18581
rect 27522 18572 27528 18624
rect 27580 18621 27586 18624
rect 27724 18621 27752 18652
rect 27580 18615 27599 18621
rect 27587 18581 27599 18615
rect 27580 18575 27599 18581
rect 27709 18615 27767 18621
rect 27709 18581 27721 18615
rect 27755 18581 27767 18615
rect 28258 18612 28264 18624
rect 28219 18584 28264 18612
rect 27709 18575 27767 18581
rect 27580 18572 27586 18575
rect 28258 18572 28264 18584
rect 28316 18572 28322 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 9030 18368 9036 18420
rect 9088 18408 9094 18420
rect 9585 18411 9643 18417
rect 9585 18408 9597 18411
rect 9088 18380 9597 18408
rect 9088 18368 9094 18380
rect 9585 18377 9597 18380
rect 9631 18377 9643 18411
rect 9585 18371 9643 18377
rect 10229 18411 10287 18417
rect 10229 18377 10241 18411
rect 10275 18408 10287 18411
rect 10318 18408 10324 18420
rect 10275 18380 10324 18408
rect 10275 18377 10287 18380
rect 10229 18371 10287 18377
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 11609 18411 11667 18417
rect 11609 18377 11621 18411
rect 11655 18408 11667 18411
rect 12066 18408 12072 18420
rect 11655 18380 12072 18408
rect 11655 18377 11667 18380
rect 11609 18371 11667 18377
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 14369 18411 14427 18417
rect 14369 18377 14381 18411
rect 14415 18408 14427 18411
rect 14826 18408 14832 18420
rect 14415 18380 14832 18408
rect 14415 18377 14427 18380
rect 14369 18371 14427 18377
rect 14826 18368 14832 18380
rect 14884 18368 14890 18420
rect 16666 18368 16672 18420
rect 16724 18408 16730 18420
rect 16853 18411 16911 18417
rect 16853 18408 16865 18411
rect 16724 18380 16865 18408
rect 16724 18368 16730 18380
rect 16853 18377 16865 18380
rect 16899 18408 16911 18411
rect 18509 18411 18567 18417
rect 16899 18380 18460 18408
rect 16899 18377 16911 18380
rect 16853 18371 16911 18377
rect 2041 18343 2099 18349
rect 2041 18309 2053 18343
rect 2087 18340 2099 18343
rect 2087 18312 15608 18340
rect 2087 18309 2099 18312
rect 2041 18303 2099 18309
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18272 9643 18275
rect 9858 18272 9864 18284
rect 9631 18244 9864 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 10137 18275 10195 18281
rect 10137 18241 10149 18275
rect 10183 18272 10195 18275
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 10183 18244 11529 18272
rect 10183 18241 10195 18244
rect 10137 18235 10195 18241
rect 11517 18241 11529 18244
rect 11563 18272 11575 18275
rect 11698 18272 11704 18284
rect 11563 18244 11704 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 13265 18275 13323 18281
rect 13265 18241 13277 18275
rect 13311 18272 13323 18275
rect 13446 18272 13452 18284
rect 13311 18244 13452 18272
rect 13311 18241 13323 18244
rect 13265 18235 13323 18241
rect 13446 18232 13452 18244
rect 13504 18232 13510 18284
rect 14277 18275 14335 18281
rect 14277 18241 14289 18275
rect 14323 18272 14335 18275
rect 14458 18272 14464 18284
rect 14323 18244 14464 18272
rect 14323 18241 14335 18244
rect 14277 18235 14335 18241
rect 14458 18232 14464 18244
rect 14516 18272 14522 18284
rect 14826 18272 14832 18284
rect 14516 18244 14832 18272
rect 14516 18232 14522 18244
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18241 15531 18275
rect 15580 18272 15608 18312
rect 16390 18300 16396 18352
rect 16448 18340 16454 18352
rect 17037 18343 17095 18349
rect 17037 18340 17049 18343
rect 16448 18312 17049 18340
rect 16448 18300 16454 18312
rect 17037 18309 17049 18312
rect 17083 18309 17095 18343
rect 17037 18303 17095 18309
rect 17494 18300 17500 18352
rect 17552 18340 17558 18352
rect 18141 18343 18199 18349
rect 18141 18340 18153 18343
rect 17552 18312 18153 18340
rect 17552 18300 17558 18312
rect 18141 18309 18153 18312
rect 18187 18309 18199 18343
rect 18432 18340 18460 18380
rect 18509 18377 18521 18411
rect 18555 18408 18567 18411
rect 19426 18408 19432 18420
rect 18555 18380 19432 18408
rect 18555 18377 18567 18380
rect 18509 18371 18567 18377
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 20070 18408 20076 18420
rect 20031 18380 20076 18408
rect 20070 18368 20076 18380
rect 20128 18368 20134 18420
rect 20530 18368 20536 18420
rect 20588 18408 20594 18420
rect 22005 18411 22063 18417
rect 22005 18408 22017 18411
rect 20588 18380 22017 18408
rect 20588 18368 20594 18380
rect 22005 18377 22017 18380
rect 22051 18377 22063 18411
rect 22646 18408 22652 18420
rect 22607 18380 22652 18408
rect 22005 18371 22063 18377
rect 22646 18368 22652 18380
rect 22704 18368 22710 18420
rect 28258 18408 28264 18420
rect 27264 18380 28264 18408
rect 22922 18340 22928 18352
rect 18432 18312 22928 18340
rect 18141 18303 18199 18309
rect 22922 18300 22928 18312
rect 22980 18300 22986 18352
rect 24210 18340 24216 18352
rect 24171 18312 24216 18340
rect 24210 18300 24216 18312
rect 24268 18300 24274 18352
rect 27264 18349 27292 18380
rect 28258 18368 28264 18380
rect 28316 18368 28322 18420
rect 47670 18408 47676 18420
rect 47631 18380 47676 18408
rect 47670 18368 47676 18380
rect 47728 18368 47734 18420
rect 27249 18343 27307 18349
rect 27249 18309 27261 18343
rect 27295 18309 27307 18343
rect 27249 18303 27307 18309
rect 27982 18300 27988 18352
rect 28040 18300 28046 18352
rect 16850 18272 16856 18284
rect 15580 18244 16856 18272
rect 15473 18235 15531 18241
rect 13354 18204 13360 18216
rect 13315 18176 13360 18204
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 13630 18204 13636 18216
rect 13591 18176 13636 18204
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 15289 18207 15347 18213
rect 15289 18173 15301 18207
rect 15335 18173 15347 18207
rect 15488 18204 15516 18235
rect 16850 18232 16856 18244
rect 16908 18232 16914 18284
rect 16942 18232 16948 18284
rect 17000 18272 17006 18284
rect 18325 18275 18383 18281
rect 17000 18244 17045 18272
rect 17000 18232 17006 18244
rect 18325 18241 18337 18275
rect 18371 18272 18383 18275
rect 18414 18272 18420 18284
rect 18371 18244 18420 18272
rect 18371 18241 18383 18244
rect 18325 18235 18383 18241
rect 18414 18232 18420 18244
rect 18472 18232 18478 18284
rect 18506 18232 18512 18284
rect 18564 18272 18570 18284
rect 19705 18275 19763 18281
rect 19705 18272 19717 18275
rect 18564 18244 19717 18272
rect 18564 18232 18570 18244
rect 19705 18241 19717 18244
rect 19751 18241 19763 18275
rect 19705 18235 19763 18241
rect 20254 18232 20260 18284
rect 20312 18272 20318 18284
rect 20717 18275 20775 18281
rect 20717 18272 20729 18275
rect 20312 18244 20729 18272
rect 20312 18232 20318 18244
rect 20717 18241 20729 18244
rect 20763 18272 20775 18275
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 20763 18244 21833 18272
rect 20763 18241 20775 18244
rect 20717 18235 20775 18241
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 22557 18275 22615 18281
rect 22557 18241 22569 18275
rect 22603 18272 22615 18275
rect 23198 18272 23204 18284
rect 22603 18244 23204 18272
rect 22603 18241 22615 18244
rect 22557 18235 22615 18241
rect 23198 18232 23204 18244
rect 23256 18232 23262 18284
rect 46382 18272 46388 18284
rect 46343 18244 46388 18272
rect 46382 18232 46388 18244
rect 46440 18232 46446 18284
rect 47026 18272 47032 18284
rect 46987 18244 47032 18272
rect 47026 18232 47032 18244
rect 47084 18232 47090 18284
rect 47578 18272 47584 18284
rect 47539 18244 47584 18272
rect 47578 18232 47584 18244
rect 47636 18232 47642 18284
rect 15654 18204 15660 18216
rect 15488 18176 15660 18204
rect 15289 18167 15347 18173
rect 15304 18136 15332 18167
rect 15654 18164 15660 18176
rect 15712 18204 15718 18216
rect 17221 18207 17279 18213
rect 17221 18204 17233 18207
rect 15712 18176 17233 18204
rect 15712 18164 15718 18176
rect 17221 18173 17233 18176
rect 17267 18173 17279 18207
rect 17221 18167 17279 18173
rect 19334 18164 19340 18216
rect 19392 18204 19398 18216
rect 19613 18207 19671 18213
rect 19613 18204 19625 18207
rect 19392 18176 19625 18204
rect 19392 18164 19398 18176
rect 19613 18173 19625 18176
rect 19659 18173 19671 18207
rect 19613 18167 19671 18173
rect 24029 18207 24087 18213
rect 24029 18173 24041 18207
rect 24075 18204 24087 18207
rect 24578 18204 24584 18216
rect 24075 18176 24584 18204
rect 24075 18173 24087 18176
rect 24029 18167 24087 18173
rect 24578 18164 24584 18176
rect 24636 18164 24642 18216
rect 24854 18204 24860 18216
rect 24815 18176 24860 18204
rect 24854 18164 24860 18176
rect 24912 18164 24918 18216
rect 26970 18204 26976 18216
rect 26931 18176 26976 18204
rect 26970 18164 26976 18176
rect 27028 18164 27034 18216
rect 16666 18136 16672 18148
rect 15304 18108 15792 18136
rect 16627 18108 16672 18136
rect 14274 18028 14280 18080
rect 14332 18068 14338 18080
rect 15657 18071 15715 18077
rect 15657 18068 15669 18071
rect 14332 18040 15669 18068
rect 14332 18028 14338 18040
rect 15657 18037 15669 18040
rect 15703 18037 15715 18071
rect 15764 18068 15792 18108
rect 16666 18096 16672 18108
rect 16724 18136 16730 18148
rect 17126 18136 17132 18148
rect 16724 18108 17132 18136
rect 16724 18096 16730 18108
rect 17126 18096 17132 18108
rect 17184 18096 17190 18148
rect 17494 18068 17500 18080
rect 15764 18040 17500 18068
rect 15657 18031 15715 18037
rect 17494 18028 17500 18040
rect 17552 18028 17558 18080
rect 20714 18068 20720 18080
rect 20675 18040 20720 18068
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 22738 18028 22744 18080
rect 22796 18068 22802 18080
rect 23293 18071 23351 18077
rect 23293 18068 23305 18071
rect 22796 18040 23305 18068
rect 22796 18028 22802 18040
rect 23293 18037 23305 18040
rect 23339 18037 23351 18071
rect 23293 18031 23351 18037
rect 27338 18028 27344 18080
rect 27396 18068 27402 18080
rect 28721 18071 28779 18077
rect 28721 18068 28733 18071
rect 27396 18040 28733 18068
rect 27396 18028 27402 18040
rect 28721 18037 28733 18040
rect 28767 18068 28779 18071
rect 29086 18068 29092 18080
rect 28767 18040 29092 18068
rect 28767 18037 28779 18040
rect 28721 18031 28779 18037
rect 29086 18028 29092 18040
rect 29144 18028 29150 18080
rect 46198 18068 46204 18080
rect 46159 18040 46204 18068
rect 46198 18028 46204 18040
rect 46256 18028 46262 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 13998 17824 14004 17876
rect 14056 17864 14062 17876
rect 14277 17867 14335 17873
rect 14277 17864 14289 17867
rect 14056 17836 14289 17864
rect 14056 17824 14062 17836
rect 14277 17833 14289 17836
rect 14323 17833 14335 17867
rect 14277 17827 14335 17833
rect 16117 17867 16175 17873
rect 16117 17833 16129 17867
rect 16163 17864 16175 17867
rect 17310 17864 17316 17876
rect 16163 17836 17316 17864
rect 16163 17833 16175 17836
rect 16117 17827 16175 17833
rect 17310 17824 17316 17836
rect 17368 17824 17374 17876
rect 19334 17864 19340 17876
rect 19295 17836 19340 17864
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 19978 17824 19984 17876
rect 20036 17864 20042 17876
rect 24394 17864 24400 17876
rect 20036 17836 24400 17864
rect 20036 17824 20042 17836
rect 24394 17824 24400 17836
rect 24452 17824 24458 17876
rect 26878 17824 26884 17876
rect 26936 17864 26942 17876
rect 26973 17867 27031 17873
rect 26973 17864 26985 17867
rect 26936 17836 26985 17864
rect 26936 17824 26942 17836
rect 26973 17833 26985 17836
rect 27019 17833 27031 17867
rect 26973 17827 27031 17833
rect 27982 17824 27988 17876
rect 28040 17864 28046 17876
rect 28077 17867 28135 17873
rect 28077 17864 28089 17867
rect 28040 17836 28089 17864
rect 28040 17824 28046 17836
rect 28077 17833 28089 17836
rect 28123 17833 28135 17867
rect 28077 17827 28135 17833
rect 14461 17799 14519 17805
rect 14461 17765 14473 17799
rect 14507 17765 14519 17799
rect 14461 17759 14519 17765
rect 16301 17799 16359 17805
rect 16301 17765 16313 17799
rect 16347 17796 16359 17799
rect 16942 17796 16948 17808
rect 16347 17768 16948 17796
rect 16347 17765 16359 17768
rect 16301 17759 16359 17765
rect 12434 17620 12440 17672
rect 12492 17660 12498 17672
rect 13265 17663 13323 17669
rect 12492 17632 12537 17660
rect 12492 17620 12498 17632
rect 13265 17629 13277 17663
rect 13311 17629 13323 17663
rect 13265 17623 13323 17629
rect 13280 17592 13308 17623
rect 13354 17620 13360 17672
rect 13412 17660 13418 17672
rect 13449 17663 13507 17669
rect 13449 17660 13461 17663
rect 13412 17632 13461 17660
rect 13412 17620 13418 17632
rect 13449 17629 13461 17632
rect 13495 17660 13507 17663
rect 14476 17660 14504 17759
rect 16942 17756 16948 17768
rect 17000 17756 17006 17808
rect 16666 17688 16672 17740
rect 16724 17728 16730 17740
rect 16761 17731 16819 17737
rect 16761 17728 16773 17731
rect 16724 17700 16773 17728
rect 16724 17688 16730 17700
rect 16761 17697 16773 17700
rect 16807 17697 16819 17731
rect 18414 17728 18420 17740
rect 16761 17691 16819 17697
rect 16868 17700 18420 17728
rect 13495 17632 14504 17660
rect 13495 17629 13507 17632
rect 13449 17623 13507 17629
rect 16206 17620 16212 17672
rect 16264 17620 16270 17672
rect 16868 17660 16896 17700
rect 18414 17688 18420 17700
rect 18472 17728 18478 17740
rect 18472 17700 19472 17728
rect 18472 17688 18478 17700
rect 16776 17632 16896 17660
rect 13814 17592 13820 17604
rect 13280 17564 13820 17592
rect 13814 17552 13820 17564
rect 13872 17552 13878 17604
rect 14093 17595 14151 17601
rect 14093 17561 14105 17595
rect 14139 17561 14151 17595
rect 14093 17555 14151 17561
rect 12529 17527 12587 17533
rect 12529 17493 12541 17527
rect 12575 17524 12587 17527
rect 12710 17524 12716 17536
rect 12575 17496 12716 17524
rect 12575 17493 12587 17496
rect 12529 17487 12587 17493
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 12986 17484 12992 17536
rect 13044 17524 13050 17536
rect 13357 17527 13415 17533
rect 13357 17524 13369 17527
rect 13044 17496 13369 17524
rect 13044 17484 13050 17496
rect 13357 17493 13369 17496
rect 13403 17493 13415 17527
rect 14108 17524 14136 17555
rect 14274 17552 14280 17604
rect 14332 17601 14338 17604
rect 14332 17595 14351 17601
rect 14339 17561 14351 17595
rect 14332 17555 14351 17561
rect 15933 17595 15991 17601
rect 15933 17561 15945 17595
rect 15979 17592 15991 17595
rect 16224 17592 16252 17620
rect 15979 17564 16252 17592
rect 15979 17561 15991 17564
rect 15933 17555 15991 17561
rect 14332 17552 14338 17555
rect 14734 17524 14740 17536
rect 14108 17496 14740 17524
rect 13357 17487 13415 17493
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 16143 17527 16201 17533
rect 16143 17493 16155 17527
rect 16189 17524 16201 17527
rect 16574 17524 16580 17536
rect 16189 17496 16580 17524
rect 16189 17493 16201 17496
rect 16143 17487 16201 17493
rect 16574 17484 16580 17496
rect 16632 17484 16638 17536
rect 16776 17524 16804 17632
rect 16942 17620 16948 17672
rect 17000 17660 17006 17672
rect 17129 17663 17187 17669
rect 17129 17660 17141 17663
rect 17000 17632 17141 17660
rect 17000 17620 17006 17632
rect 17129 17629 17141 17632
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 16850 17552 16856 17604
rect 16908 17592 16914 17604
rect 17313 17595 17371 17601
rect 17313 17592 17325 17595
rect 16908 17564 17325 17592
rect 16908 17552 16914 17564
rect 17313 17561 17325 17564
rect 17359 17561 17371 17595
rect 18340 17592 18368 17623
rect 18506 17620 18512 17672
rect 18564 17660 18570 17672
rect 19444 17669 19472 17700
rect 20714 17688 20720 17740
rect 20772 17728 20778 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 20772 17700 20913 17728
rect 20772 17688 20778 17700
rect 20901 17697 20913 17700
rect 20947 17697 20959 17731
rect 20901 17691 20959 17697
rect 25501 17731 25559 17737
rect 25501 17697 25513 17731
rect 25547 17728 25559 17731
rect 25590 17728 25596 17740
rect 25547 17700 25596 17728
rect 25547 17697 25559 17700
rect 25501 17691 25559 17697
rect 25590 17688 25596 17700
rect 25648 17688 25654 17740
rect 46014 17728 46020 17740
rect 26804 17700 46020 17728
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 18564 17632 19257 17660
rect 18564 17620 18570 17632
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 25222 17660 25228 17672
rect 25183 17632 25228 17660
rect 19429 17623 19487 17629
rect 25222 17620 25228 17632
rect 25280 17620 25286 17672
rect 20254 17592 20260 17604
rect 18340 17564 20260 17592
rect 17313 17555 17371 17561
rect 20254 17552 20260 17564
rect 20312 17552 20318 17604
rect 20806 17552 20812 17604
rect 20864 17592 20870 17604
rect 21177 17595 21235 17601
rect 21177 17592 21189 17595
rect 20864 17564 21189 17592
rect 20864 17552 20870 17564
rect 21177 17561 21189 17564
rect 21223 17561 21235 17595
rect 22738 17592 22744 17604
rect 22402 17564 22744 17592
rect 21177 17555 21235 17561
rect 22738 17552 22744 17564
rect 22796 17552 22802 17604
rect 22922 17552 22928 17604
rect 22980 17592 22986 17604
rect 22980 17564 23073 17592
rect 22980 17552 22986 17564
rect 26234 17552 26240 17604
rect 26292 17552 26298 17604
rect 16945 17527 17003 17533
rect 16945 17524 16957 17527
rect 16776 17496 16957 17524
rect 16945 17493 16957 17496
rect 16991 17493 17003 17527
rect 16945 17487 17003 17493
rect 17037 17527 17095 17533
rect 17037 17493 17049 17527
rect 17083 17524 17095 17527
rect 17494 17524 17500 17536
rect 17083 17496 17500 17524
rect 17083 17493 17095 17496
rect 17037 17487 17095 17493
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 18138 17484 18144 17536
rect 18196 17524 18202 17536
rect 18417 17527 18475 17533
rect 18417 17524 18429 17527
rect 18196 17496 18429 17524
rect 18196 17484 18202 17496
rect 18417 17493 18429 17496
rect 18463 17493 18475 17527
rect 22940 17524 22968 17552
rect 26804 17524 26832 17700
rect 46014 17688 46020 17700
rect 46072 17688 46078 17740
rect 27062 17620 27068 17672
rect 27120 17660 27126 17672
rect 27985 17663 28043 17669
rect 27985 17660 27997 17663
rect 27120 17632 27997 17660
rect 27120 17620 27126 17632
rect 27985 17629 27997 17632
rect 28031 17629 28043 17663
rect 45833 17663 45891 17669
rect 27985 17623 28043 17629
rect 30668 17632 35894 17660
rect 30668 17604 30696 17632
rect 29638 17592 29644 17604
rect 29599 17564 29644 17592
rect 29638 17552 29644 17564
rect 29696 17552 29702 17604
rect 29733 17595 29791 17601
rect 29733 17561 29745 17595
rect 29779 17592 29791 17595
rect 30006 17592 30012 17604
rect 29779 17564 30012 17592
rect 29779 17561 29791 17564
rect 29733 17555 29791 17561
rect 30006 17552 30012 17564
rect 30064 17552 30070 17604
rect 30650 17592 30656 17604
rect 30563 17564 30656 17592
rect 30650 17552 30656 17564
rect 30708 17552 30714 17604
rect 22940 17496 26832 17524
rect 35866 17524 35894 17632
rect 45833 17629 45845 17663
rect 45879 17660 45891 17663
rect 46293 17663 46351 17669
rect 46293 17660 46305 17663
rect 45879 17632 46305 17660
rect 45879 17629 45891 17632
rect 45833 17623 45891 17629
rect 46293 17629 46305 17632
rect 46339 17629 46351 17663
rect 46293 17623 46351 17629
rect 46477 17595 46535 17601
rect 46477 17561 46489 17595
rect 46523 17592 46535 17595
rect 47670 17592 47676 17604
rect 46523 17564 47676 17592
rect 46523 17561 46535 17564
rect 46477 17555 46535 17561
rect 47670 17552 47676 17564
rect 47728 17552 47734 17604
rect 48130 17592 48136 17604
rect 48091 17564 48136 17592
rect 48130 17552 48136 17564
rect 48188 17552 48194 17604
rect 40218 17524 40224 17536
rect 35866 17496 40224 17524
rect 18417 17487 18475 17493
rect 40218 17484 40224 17496
rect 40276 17484 40282 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 4982 17280 4988 17332
rect 5040 17320 5046 17332
rect 5040 17292 22094 17320
rect 5040 17280 5046 17292
rect 12986 17252 12992 17264
rect 12947 17224 12992 17252
rect 12986 17212 12992 17224
rect 13044 17212 13050 17264
rect 15289 17255 15347 17261
rect 15289 17252 15301 17255
rect 14214 17224 15301 17252
rect 15289 17221 15301 17224
rect 15335 17221 15347 17255
rect 15289 17215 15347 17221
rect 19426 17212 19432 17264
rect 19484 17212 19490 17264
rect 22066 17252 22094 17292
rect 25222 17280 25228 17332
rect 25280 17320 25286 17332
rect 25317 17323 25375 17329
rect 25317 17320 25329 17323
rect 25280 17292 25329 17320
rect 25280 17280 25286 17292
rect 25317 17289 25329 17292
rect 25363 17289 25375 17323
rect 25317 17283 25375 17289
rect 25961 17323 26019 17329
rect 25961 17289 25973 17323
rect 26007 17320 26019 17323
rect 26970 17320 26976 17332
rect 26007 17292 26976 17320
rect 26007 17289 26019 17292
rect 25961 17283 26019 17289
rect 26970 17280 26976 17292
rect 27028 17280 27034 17332
rect 47670 17320 47676 17332
rect 47631 17292 47676 17320
rect 47670 17280 47676 17292
rect 47728 17280 47734 17332
rect 23658 17252 23664 17264
rect 22066 17224 23664 17252
rect 23658 17212 23664 17224
rect 23716 17212 23722 17264
rect 24394 17212 24400 17264
rect 24452 17252 24458 17264
rect 28537 17255 28595 17261
rect 24452 17224 25176 17252
rect 24452 17212 24458 17224
rect 12710 17184 12716 17196
rect 12671 17156 12716 17184
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 14826 17144 14832 17196
rect 14884 17184 14890 17196
rect 15197 17187 15255 17193
rect 15197 17184 15209 17187
rect 14884 17156 15209 17184
rect 14884 17144 14890 17156
rect 15197 17153 15209 17156
rect 15243 17153 15255 17187
rect 15838 17184 15844 17196
rect 15799 17156 15844 17184
rect 15197 17147 15255 17153
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 17310 17184 17316 17196
rect 17271 17156 17316 17184
rect 17310 17144 17316 17156
rect 17368 17144 17374 17196
rect 18138 17184 18144 17196
rect 18099 17156 18144 17184
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 25148 17193 25176 17224
rect 28537 17221 28549 17255
rect 28583 17252 28595 17255
rect 29273 17255 29331 17261
rect 29273 17252 29285 17255
rect 28583 17224 29285 17252
rect 28583 17221 28595 17224
rect 28537 17215 28595 17221
rect 29273 17221 29285 17224
rect 29319 17221 29331 17255
rect 29273 17215 29331 17221
rect 45094 17212 45100 17264
rect 45152 17252 45158 17264
rect 45373 17255 45431 17261
rect 45373 17252 45385 17255
rect 45152 17224 45385 17252
rect 45152 17212 45158 17224
rect 45373 17221 45385 17224
rect 45419 17221 45431 17255
rect 45373 17215 45431 17221
rect 47029 17255 47087 17261
rect 47029 17221 47041 17255
rect 47075 17252 47087 17255
rect 47118 17252 47124 17264
rect 47075 17224 47124 17252
rect 47075 17221 47087 17224
rect 47029 17215 47087 17221
rect 47118 17212 47124 17224
rect 47176 17212 47182 17264
rect 23477 17187 23535 17193
rect 23477 17153 23489 17187
rect 23523 17153 23535 17187
rect 23477 17147 23535 17153
rect 23845 17187 23903 17193
rect 23845 17153 23857 17187
rect 23891 17184 23903 17187
rect 24489 17187 24547 17193
rect 24489 17184 24501 17187
rect 23891 17156 24501 17184
rect 23891 17153 23903 17156
rect 23845 17147 23903 17153
rect 24489 17153 24501 17156
rect 24535 17153 24547 17187
rect 24489 17147 24547 17153
rect 25133 17187 25191 17193
rect 25133 17153 25145 17187
rect 25179 17184 25191 17187
rect 25869 17187 25927 17193
rect 25869 17184 25881 17187
rect 25179 17156 25881 17184
rect 25179 17153 25191 17156
rect 25133 17147 25191 17153
rect 25869 17153 25881 17156
rect 25915 17153 25927 17187
rect 28442 17184 28448 17196
rect 28403 17156 28448 17184
rect 25869 17147 25927 17153
rect 3326 17076 3332 17128
rect 3384 17116 3390 17128
rect 7926 17116 7932 17128
rect 3384 17088 7932 17116
rect 3384 17076 3390 17088
rect 7926 17076 7932 17088
rect 7984 17076 7990 17128
rect 14734 17116 14740 17128
rect 14695 17088 14740 17116
rect 14734 17076 14740 17088
rect 14792 17076 14798 17128
rect 17402 17116 17408 17128
rect 17363 17088 17408 17116
rect 17402 17076 17408 17088
rect 17460 17076 17466 17128
rect 18417 17119 18475 17125
rect 18417 17116 18429 17119
rect 18248 17088 18429 17116
rect 16666 17048 16672 17060
rect 15764 17020 16672 17048
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 1452 16952 2053 16980
rect 1452 16940 1458 16952
rect 2041 16949 2053 16952
rect 2087 16949 2099 16983
rect 2041 16943 2099 16949
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 15764 16980 15792 17020
rect 16666 17008 16672 17020
rect 16724 17008 16730 17060
rect 17681 17051 17739 17057
rect 17681 17017 17693 17051
rect 17727 17048 17739 17051
rect 18248 17048 18276 17088
rect 18417 17085 18429 17088
rect 18463 17085 18475 17119
rect 18417 17079 18475 17085
rect 23492 17060 23520 17147
rect 28442 17144 28448 17156
rect 28500 17144 28506 17196
rect 29086 17184 29092 17196
rect 29047 17156 29092 17184
rect 29086 17144 29092 17156
rect 29144 17144 29150 17196
rect 46842 17144 46848 17196
rect 46900 17184 46906 17196
rect 47394 17184 47400 17196
rect 46900 17156 47400 17184
rect 46900 17144 46906 17156
rect 47394 17144 47400 17156
rect 47452 17184 47458 17196
rect 47581 17187 47639 17193
rect 47581 17184 47593 17187
rect 47452 17156 47593 17184
rect 47452 17144 47458 17156
rect 47581 17153 47593 17156
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 23750 17076 23756 17128
rect 23808 17116 23814 17128
rect 24305 17119 24363 17125
rect 24305 17116 24317 17119
rect 23808 17088 24317 17116
rect 23808 17076 23814 17088
rect 24305 17085 24317 17088
rect 24351 17085 24363 17119
rect 30926 17116 30932 17128
rect 30887 17088 30932 17116
rect 24305 17079 24363 17085
rect 30926 17076 30932 17088
rect 30984 17076 30990 17128
rect 45186 17116 45192 17128
rect 45147 17088 45192 17116
rect 45186 17076 45192 17088
rect 45244 17076 45250 17128
rect 23474 17048 23480 17060
rect 17727 17020 18276 17048
rect 23387 17020 23480 17048
rect 17727 17017 17739 17020
rect 17681 17011 17739 17017
rect 23474 17008 23480 17020
rect 23532 17048 23538 17060
rect 30650 17048 30656 17060
rect 23532 17020 30656 17048
rect 23532 17008 23538 17020
rect 30650 17008 30656 17020
rect 30708 17008 30714 17060
rect 10744 16952 15792 16980
rect 10744 16940 10750 16952
rect 15838 16940 15844 16992
rect 15896 16980 15902 16992
rect 15933 16983 15991 16989
rect 15933 16980 15945 16983
rect 15896 16952 15945 16980
rect 15896 16940 15902 16952
rect 15933 16949 15945 16952
rect 15979 16949 15991 16983
rect 15933 16943 15991 16949
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 19889 16983 19947 16989
rect 19889 16980 19901 16983
rect 17368 16952 19901 16980
rect 17368 16940 17374 16952
rect 19889 16949 19901 16952
rect 19935 16949 19947 16983
rect 19889 16943 19947 16949
rect 24673 16983 24731 16989
rect 24673 16949 24685 16983
rect 24719 16980 24731 16983
rect 24854 16980 24860 16992
rect 24719 16952 24860 16980
rect 24719 16949 24731 16952
rect 24673 16943 24731 16949
rect 24854 16940 24860 16952
rect 24912 16940 24918 16992
rect 39758 16940 39764 16992
rect 39816 16980 39822 16992
rect 45462 16980 45468 16992
rect 39816 16952 45468 16980
rect 39816 16940 39822 16952
rect 45462 16940 45468 16952
rect 45520 16940 45526 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 10704 16748 12434 16776
rect 10704 16708 10732 16748
rect 2746 16680 10732 16708
rect 12406 16708 12434 16748
rect 13814 16736 13820 16788
rect 13872 16776 13878 16788
rect 14093 16779 14151 16785
rect 14093 16776 14105 16779
rect 13872 16748 14105 16776
rect 13872 16736 13878 16748
rect 14093 16745 14105 16748
rect 14139 16745 14151 16779
rect 20990 16776 20996 16788
rect 14093 16739 14151 16745
rect 14660 16748 20996 16776
rect 14660 16708 14688 16748
rect 20990 16736 20996 16748
rect 21048 16776 21054 16788
rect 29638 16776 29644 16788
rect 21048 16748 29644 16776
rect 21048 16736 21054 16748
rect 29638 16736 29644 16748
rect 29696 16736 29702 16788
rect 45922 16776 45928 16788
rect 39868 16748 45928 16776
rect 12406 16680 14688 16708
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 2314 16600 2320 16652
rect 2372 16640 2378 16652
rect 2746 16640 2774 16680
rect 14734 16668 14740 16720
rect 14792 16708 14798 16720
rect 14792 16680 26234 16708
rect 14792 16668 14798 16680
rect 2372 16612 2774 16640
rect 2372 16600 2378 16612
rect 3418 16600 3424 16652
rect 3476 16640 3482 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 3476 16612 11161 16640
rect 3476 16600 3482 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 13078 16600 13084 16652
rect 13136 16640 13142 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 13136 16612 15669 16640
rect 13136 16600 13142 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15838 16640 15844 16652
rect 15799 16612 15844 16640
rect 15657 16603 15715 16609
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 20990 16640 20996 16652
rect 20951 16612 20996 16640
rect 20990 16600 20996 16612
rect 21048 16600 21054 16652
rect 24486 16600 24492 16652
rect 24544 16640 24550 16652
rect 25133 16643 25191 16649
rect 25133 16640 25145 16643
rect 24544 16612 25145 16640
rect 24544 16600 24550 16612
rect 25133 16609 25145 16612
rect 25179 16640 25191 16643
rect 25406 16640 25412 16652
rect 25179 16612 25412 16640
rect 25179 16609 25191 16612
rect 25133 16603 25191 16609
rect 25406 16600 25412 16612
rect 25464 16600 25470 16652
rect 26206 16640 26234 16680
rect 30009 16643 30067 16649
rect 30009 16640 30021 16643
rect 26206 16612 30021 16640
rect 30009 16609 30021 16612
rect 30055 16609 30067 16643
rect 30009 16603 30067 16609
rect 31849 16643 31907 16649
rect 31849 16609 31861 16643
rect 31895 16640 31907 16643
rect 39758 16640 39764 16652
rect 31895 16612 39764 16640
rect 31895 16609 31907 16612
rect 31849 16603 31907 16609
rect 39758 16600 39764 16612
rect 39816 16600 39822 16652
rect 39868 16640 39896 16748
rect 45922 16736 45928 16748
rect 45980 16736 45986 16788
rect 39945 16643 40003 16649
rect 39945 16640 39957 16643
rect 39868 16612 39957 16640
rect 39945 16609 39957 16612
rect 39991 16609 40003 16643
rect 40218 16640 40224 16652
rect 40179 16612 40224 16640
rect 39945 16603 40003 16609
rect 40218 16600 40224 16612
rect 40276 16600 40282 16652
rect 46293 16643 46351 16649
rect 46293 16609 46305 16643
rect 46339 16640 46351 16643
rect 47026 16640 47032 16652
rect 46339 16612 47032 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47026 16600 47032 16612
rect 47084 16600 47090 16652
rect 10686 16572 10692 16584
rect 10647 16544 10692 16572
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 14274 16532 14280 16584
rect 14332 16572 14338 16584
rect 14369 16575 14427 16581
rect 14369 16572 14381 16575
rect 14332 16544 14381 16572
rect 14332 16532 14338 16544
rect 14369 16541 14381 16544
rect 14415 16541 14427 16575
rect 19334 16572 19340 16584
rect 14369 16535 14427 16541
rect 17052 16544 19340 16572
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 2130 16504 2136 16516
rect 1627 16476 2136 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 10870 16504 10876 16516
rect 10831 16476 10876 16504
rect 10870 16464 10876 16476
rect 10928 16464 10934 16516
rect 14093 16507 14151 16513
rect 14093 16473 14105 16507
rect 14139 16504 14151 16507
rect 14734 16504 14740 16516
rect 14139 16476 14740 16504
rect 14139 16473 14151 16476
rect 14093 16467 14151 16473
rect 14734 16464 14740 16476
rect 14792 16464 14798 16516
rect 15838 16464 15844 16516
rect 15896 16504 15902 16516
rect 17052 16504 17080 16544
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16572 19763 16575
rect 19978 16572 19984 16584
rect 19751 16544 19984 16572
rect 19751 16541 19763 16544
rect 19705 16535 19763 16541
rect 19978 16532 19984 16544
rect 20036 16532 20042 16584
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16572 23443 16575
rect 23474 16572 23480 16584
rect 23431 16544 23480 16572
rect 23431 16541 23443 16544
rect 23385 16535 23443 16541
rect 23474 16532 23480 16544
rect 23532 16532 23538 16584
rect 23658 16572 23664 16584
rect 23619 16544 23664 16572
rect 23658 16532 23664 16544
rect 23716 16532 23722 16584
rect 24854 16572 24860 16584
rect 24815 16544 24860 16572
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 45646 16532 45652 16584
rect 45704 16572 45710 16584
rect 46014 16572 46020 16584
rect 45704 16544 46020 16572
rect 45704 16532 45710 16544
rect 46014 16532 46020 16544
rect 46072 16532 46078 16584
rect 17494 16504 17500 16516
rect 15896 16476 17080 16504
rect 17455 16476 17500 16504
rect 15896 16464 15902 16476
rect 17494 16464 17500 16476
rect 17552 16464 17558 16516
rect 21085 16507 21143 16513
rect 21085 16473 21097 16507
rect 21131 16473 21143 16507
rect 22002 16504 22008 16516
rect 21963 16476 22008 16504
rect 21085 16467 21143 16473
rect 13998 16396 14004 16448
rect 14056 16436 14062 16448
rect 14277 16439 14335 16445
rect 14277 16436 14289 16439
rect 14056 16408 14289 16436
rect 14056 16396 14062 16408
rect 14277 16405 14289 16408
rect 14323 16436 14335 16439
rect 15102 16436 15108 16448
rect 14323 16408 15108 16436
rect 14323 16405 14335 16408
rect 14277 16399 14335 16405
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 19797 16439 19855 16445
rect 19797 16436 19809 16439
rect 19392 16408 19809 16436
rect 19392 16396 19398 16408
rect 19797 16405 19809 16408
rect 19843 16405 19855 16439
rect 19797 16399 19855 16405
rect 20162 16396 20168 16448
rect 20220 16436 20226 16448
rect 21100 16436 21128 16467
rect 22002 16464 22008 16476
rect 22060 16464 22066 16516
rect 23750 16504 23756 16516
rect 23711 16476 23756 16504
rect 23750 16464 23756 16476
rect 23808 16464 23814 16516
rect 30190 16504 30196 16516
rect 30151 16476 30196 16504
rect 30190 16464 30196 16476
rect 30248 16464 30254 16516
rect 40037 16507 40095 16513
rect 40037 16473 40049 16507
rect 40083 16504 40095 16507
rect 40402 16504 40408 16516
rect 40083 16476 40408 16504
rect 40083 16473 40095 16476
rect 40037 16467 40095 16473
rect 40402 16464 40408 16476
rect 40460 16464 40466 16516
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 47670 16504 47676 16516
rect 46523 16476 47676 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 47670 16464 47676 16476
rect 47728 16464 47734 16516
rect 48130 16504 48136 16516
rect 48091 16476 48136 16504
rect 48130 16464 48136 16476
rect 48188 16464 48194 16516
rect 20220 16408 21128 16436
rect 20220 16396 20226 16408
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 10870 16232 10876 16244
rect 10831 16204 10876 16232
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 16574 16192 16580 16244
rect 16632 16232 16638 16244
rect 17221 16235 17279 16241
rect 17221 16232 17233 16235
rect 16632 16204 17233 16232
rect 16632 16192 16638 16204
rect 17221 16201 17233 16204
rect 17267 16232 17279 16235
rect 17310 16232 17316 16244
rect 17267 16204 17316 16232
rect 17267 16201 17279 16204
rect 17221 16195 17279 16201
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 19245 16235 19303 16241
rect 19245 16201 19257 16235
rect 19291 16232 19303 16235
rect 19426 16232 19432 16244
rect 19291 16204 19432 16232
rect 19291 16201 19303 16204
rect 19245 16195 19303 16201
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 30190 16232 30196 16244
rect 30151 16204 30196 16232
rect 30190 16192 30196 16204
rect 30248 16192 30254 16244
rect 46474 16232 46480 16244
rect 35866 16204 46480 16232
rect 15838 16164 15844 16176
rect 2746 16136 15844 16164
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 2004 16068 2053 16096
rect 2004 16056 2010 16068
rect 2041 16065 2053 16068
rect 2087 16096 2099 16099
rect 2746 16096 2774 16136
rect 15838 16124 15844 16136
rect 15896 16124 15902 16176
rect 16206 16124 16212 16176
rect 16264 16164 16270 16176
rect 17037 16167 17095 16173
rect 17037 16164 17049 16167
rect 16264 16136 17049 16164
rect 16264 16124 16270 16136
rect 17037 16133 17049 16136
rect 17083 16164 17095 16167
rect 18046 16164 18052 16176
rect 17083 16136 18052 16164
rect 17083 16133 17095 16136
rect 17037 16127 17095 16133
rect 18046 16124 18052 16136
rect 18104 16124 18110 16176
rect 24578 16124 24584 16176
rect 24636 16124 24642 16176
rect 2087 16068 2774 16096
rect 10781 16099 10839 16105
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 10781 16065 10793 16099
rect 10827 16096 10839 16099
rect 11054 16096 11060 16108
rect 10827 16068 11060 16096
rect 10827 16065 10839 16068
rect 10781 16059 10839 16065
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16666 16096 16672 16108
rect 16163 16068 16672 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 15948 16028 15976 16059
rect 16666 16056 16672 16068
rect 16724 16096 16730 16108
rect 16850 16096 16856 16108
rect 16724 16068 16856 16096
rect 16724 16056 16730 16068
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16096 17371 16099
rect 17402 16096 17408 16108
rect 17359 16068 17408 16096
rect 17359 16065 17371 16068
rect 17313 16059 17371 16065
rect 17402 16056 17408 16068
rect 17460 16056 17466 16108
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16096 18383 16099
rect 18598 16096 18604 16108
rect 18371 16068 18604 16096
rect 18371 16065 18383 16068
rect 18325 16059 18383 16065
rect 18598 16056 18604 16068
rect 18656 16096 18662 16108
rect 19153 16099 19211 16105
rect 19153 16096 19165 16099
rect 18656 16068 19165 16096
rect 18656 16056 18662 16068
rect 19153 16065 19165 16068
rect 19199 16096 19211 16099
rect 19242 16096 19248 16108
rect 19199 16068 19248 16096
rect 19199 16065 19211 16068
rect 19153 16059 19211 16065
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 23750 16096 23756 16108
rect 23711 16068 23756 16096
rect 23750 16056 23756 16068
rect 23808 16056 23814 16108
rect 24394 16096 24400 16108
rect 24355 16068 24400 16096
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 30098 16096 30104 16108
rect 30011 16068 30104 16096
rect 30098 16056 30104 16068
rect 30156 16096 30162 16108
rect 35866 16096 35894 16204
rect 46474 16192 46480 16204
rect 46532 16192 46538 16244
rect 47670 16232 47676 16244
rect 47631 16204 47676 16232
rect 47670 16192 47676 16204
rect 47728 16192 47734 16244
rect 46658 16124 46664 16176
rect 46716 16164 46722 16176
rect 46934 16164 46940 16176
rect 46716 16136 46940 16164
rect 46716 16124 46722 16136
rect 46934 16124 46940 16136
rect 46992 16164 46998 16176
rect 46992 16136 47624 16164
rect 46992 16124 46998 16136
rect 47026 16096 47032 16108
rect 30156 16068 35894 16096
rect 46987 16068 47032 16096
rect 30156 16056 30162 16068
rect 47026 16056 47032 16068
rect 47084 16056 47090 16108
rect 47596 16105 47624 16136
rect 47581 16099 47639 16105
rect 47581 16065 47593 16099
rect 47627 16065 47639 16099
rect 47581 16059 47639 16065
rect 15948 16000 17080 16028
rect 17052 15969 17080 16000
rect 17037 15963 17095 15969
rect 17037 15929 17049 15963
rect 17083 15929 17095 15963
rect 17037 15923 17095 15929
rect 15933 15895 15991 15901
rect 15933 15861 15945 15895
rect 15979 15892 15991 15895
rect 17218 15892 17224 15904
rect 15979 15864 17224 15892
rect 15979 15861 15991 15864
rect 15933 15855 15991 15861
rect 17218 15852 17224 15864
rect 17276 15852 17282 15904
rect 18322 15852 18328 15904
rect 18380 15892 18386 15904
rect 18417 15895 18475 15901
rect 18417 15892 18429 15895
rect 18380 15864 18429 15892
rect 18380 15852 18386 15864
rect 18417 15861 18429 15864
rect 18463 15861 18475 15895
rect 18417 15855 18475 15861
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 18966 15648 18972 15700
rect 19024 15688 19030 15700
rect 19024 15660 21036 15688
rect 19024 15648 19030 15660
rect 2038 15580 2044 15632
rect 2096 15620 2102 15632
rect 21008 15620 21036 15660
rect 22002 15648 22008 15700
rect 22060 15688 22066 15700
rect 23109 15691 23167 15697
rect 23109 15688 23121 15691
rect 22060 15660 23121 15688
rect 22060 15648 22066 15660
rect 23109 15657 23121 15660
rect 23155 15688 23167 15691
rect 23934 15688 23940 15700
rect 23155 15660 23940 15688
rect 23155 15657 23167 15660
rect 23109 15651 23167 15657
rect 23934 15648 23940 15660
rect 23992 15648 23998 15700
rect 24394 15648 24400 15700
rect 24452 15688 24458 15700
rect 24489 15691 24547 15697
rect 24489 15688 24501 15691
rect 24452 15660 24501 15688
rect 24452 15648 24458 15660
rect 24489 15657 24501 15660
rect 24535 15657 24547 15691
rect 24489 15651 24547 15657
rect 27062 15620 27068 15632
rect 2096 15592 20852 15620
rect 21008 15592 27068 15620
rect 2096 15580 2102 15592
rect 9214 15512 9220 15564
rect 9272 15552 9278 15564
rect 10137 15555 10195 15561
rect 10137 15552 10149 15555
rect 9272 15524 10149 15552
rect 9272 15512 9278 15524
rect 10137 15521 10149 15524
rect 10183 15521 10195 15555
rect 10137 15515 10195 15521
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15521 13139 15555
rect 13354 15552 13360 15564
rect 13315 15524 13360 15552
rect 13081 15515 13139 15521
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 9674 15484 9680 15496
rect 9635 15456 9680 15484
rect 2041 15447 2099 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15453 13047 15487
rect 13096 15484 13124 15515
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 14274 15552 14280 15564
rect 13464 15524 14280 15552
rect 13464 15484 13492 15524
rect 14274 15512 14280 15524
rect 14332 15552 14338 15564
rect 15010 15552 15016 15564
rect 14332 15524 15016 15552
rect 14332 15512 14338 15524
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15552 15991 15555
rect 16206 15552 16212 15564
rect 15979 15524 16212 15552
rect 15979 15521 15991 15524
rect 15933 15515 15991 15521
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 20824 15561 20852 15592
rect 21100 15561 21128 15592
rect 27062 15580 27068 15592
rect 27120 15580 27126 15632
rect 20809 15555 20867 15561
rect 20809 15521 20821 15555
rect 20855 15521 20867 15555
rect 20809 15515 20867 15521
rect 21085 15555 21143 15561
rect 21085 15521 21097 15555
rect 21131 15552 21143 15555
rect 23385 15555 23443 15561
rect 21131 15524 21165 15552
rect 21131 15521 21143 15524
rect 21085 15515 21143 15521
rect 23385 15521 23397 15555
rect 23431 15552 23443 15555
rect 23474 15552 23480 15564
rect 23431 15524 23480 15552
rect 23431 15521 23443 15524
rect 23385 15515 23443 15521
rect 23474 15512 23480 15524
rect 23532 15512 23538 15564
rect 23750 15512 23756 15564
rect 23808 15552 23814 15564
rect 47949 15555 48007 15561
rect 47949 15552 47961 15555
rect 23808 15524 24624 15552
rect 23808 15512 23814 15524
rect 13096 15456 13492 15484
rect 12989 15447 13047 15453
rect 9858 15416 9864 15428
rect 9819 15388 9864 15416
rect 9858 15376 9864 15388
rect 9916 15376 9922 15428
rect 13004 15416 13032 15447
rect 13630 15444 13636 15496
rect 13688 15484 13694 15496
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13688 15456 14105 15484
rect 13688 15444 13694 15456
rect 14093 15453 14105 15456
rect 14139 15486 14151 15487
rect 14139 15484 14228 15486
rect 14826 15484 14832 15496
rect 14139 15458 14688 15484
rect 14139 15453 14151 15458
rect 14200 15456 14688 15458
rect 14787 15456 14832 15484
rect 14093 15447 14151 15453
rect 13998 15416 14004 15428
rect 13004 15388 14004 15416
rect 13998 15376 14004 15388
rect 14056 15376 14062 15428
rect 14660 15416 14688 15456
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 18233 15487 18291 15493
rect 18233 15484 18245 15487
rect 17328 15456 18245 15484
rect 16114 15416 16120 15428
rect 14660 15388 15976 15416
rect 16075 15388 16120 15416
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14277 15351 14335 15357
rect 14277 15348 14289 15351
rect 13872 15320 14289 15348
rect 13872 15308 13878 15320
rect 14277 15317 14289 15320
rect 14323 15317 14335 15351
rect 14918 15348 14924 15360
rect 14879 15320 14924 15348
rect 14277 15311 14335 15317
rect 14918 15308 14924 15320
rect 14976 15308 14982 15360
rect 15948 15348 15976 15388
rect 16114 15376 16120 15388
rect 16172 15376 16178 15428
rect 17328 15348 17356 15456
rect 18233 15453 18245 15456
rect 18279 15484 18291 15487
rect 19334 15484 19340 15496
rect 18279 15456 19340 15484
rect 18279 15453 18291 15456
rect 18233 15447 18291 15453
rect 19334 15444 19340 15456
rect 19392 15484 19398 15496
rect 19978 15484 19984 15496
rect 19392 15456 19984 15484
rect 19392 15444 19398 15456
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 20625 15487 20683 15493
rect 20625 15453 20637 15487
rect 20671 15453 20683 15487
rect 20625 15447 20683 15453
rect 17770 15416 17776 15428
rect 17731 15388 17776 15416
rect 17770 15376 17776 15388
rect 17828 15376 17834 15428
rect 15948 15320 17356 15348
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18417 15351 18475 15357
rect 18417 15348 18429 15351
rect 18012 15320 18429 15348
rect 18012 15308 18018 15320
rect 18417 15317 18429 15320
rect 18463 15317 18475 15351
rect 20640 15348 20668 15447
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 23017 15487 23075 15493
rect 23017 15484 23029 15487
rect 22152 15456 23029 15484
rect 22152 15444 22158 15456
rect 23017 15453 23029 15456
rect 23063 15453 23075 15487
rect 23017 15447 23075 15453
rect 23293 15487 23351 15493
rect 23293 15453 23305 15487
rect 23339 15484 23351 15487
rect 23658 15484 23664 15496
rect 23339 15456 23664 15484
rect 23339 15453 23351 15456
rect 23293 15447 23351 15453
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 24596 15493 24624 15524
rect 47044 15524 47961 15552
rect 24489 15487 24547 15493
rect 24489 15453 24501 15487
rect 24535 15453 24547 15487
rect 24489 15447 24547 15453
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15453 24639 15487
rect 46382 15484 46388 15496
rect 46343 15456 46388 15484
rect 24581 15447 24639 15453
rect 23842 15416 23848 15428
rect 23216 15388 23848 15416
rect 23216 15348 23244 15388
rect 23842 15376 23848 15388
rect 23900 15376 23906 15428
rect 24504 15416 24532 15447
rect 46382 15444 46388 15456
rect 46440 15444 46446 15496
rect 47044 15470 47072 15524
rect 47949 15521 47961 15524
rect 47995 15521 48007 15555
rect 47949 15515 48007 15521
rect 47854 15484 47860 15496
rect 47815 15456 47860 15484
rect 47854 15444 47860 15456
rect 47912 15444 47918 15496
rect 48041 15487 48099 15493
rect 48041 15453 48053 15487
rect 48087 15453 48099 15487
rect 48041 15447 48099 15453
rect 24854 15416 24860 15428
rect 24504 15388 24860 15416
rect 24854 15376 24860 15388
rect 24912 15376 24918 15428
rect 45186 15376 45192 15428
rect 45244 15416 45250 15428
rect 47121 15419 47179 15425
rect 47121 15416 47133 15419
rect 45244 15388 47133 15416
rect 45244 15376 45250 15388
rect 47121 15385 47133 15388
rect 47167 15385 47179 15419
rect 48056 15416 48084 15447
rect 47121 15379 47179 15385
rect 47872 15388 48084 15416
rect 47872 15360 47900 15388
rect 23382 15348 23388 15360
rect 20640 15320 23244 15348
rect 23343 15320 23388 15348
rect 18417 15311 18475 15317
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 47854 15308 47860 15360
rect 47912 15308 47918 15360
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 9858 15104 9864 15156
rect 9916 15144 9922 15156
rect 10413 15147 10471 15153
rect 10413 15144 10425 15147
rect 9916 15116 10425 15144
rect 9916 15104 9922 15116
rect 10413 15113 10425 15116
rect 10459 15113 10471 15147
rect 10413 15107 10471 15113
rect 16025 15147 16083 15153
rect 16025 15113 16037 15147
rect 16071 15144 16083 15147
rect 16114 15144 16120 15156
rect 16071 15116 16120 15144
rect 16071 15113 16083 15116
rect 16025 15107 16083 15113
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 17954 15144 17960 15156
rect 16960 15116 17960 15144
rect 13354 15036 13360 15088
rect 13412 15076 13418 15088
rect 13449 15079 13507 15085
rect 13449 15076 13461 15079
rect 13412 15048 13461 15076
rect 13412 15036 13418 15048
rect 13449 15045 13461 15048
rect 13495 15045 13507 15079
rect 14918 15076 14924 15088
rect 14674 15048 14924 15076
rect 13449 15039 13507 15045
rect 14918 15036 14924 15048
rect 14976 15036 14982 15088
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 11054 15008 11060 15020
rect 10367 14980 11060 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 15930 15008 15936 15020
rect 15891 14980 15936 15008
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 16960 15017 16988 15116
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 18693 15147 18751 15153
rect 18693 15144 18705 15147
rect 18104 15116 18705 15144
rect 18104 15104 18110 15116
rect 18693 15113 18705 15116
rect 18739 15113 18751 15147
rect 18693 15107 18751 15113
rect 22189 15147 22247 15153
rect 22189 15113 22201 15147
rect 22235 15144 22247 15147
rect 23750 15144 23756 15156
rect 22235 15116 23756 15144
rect 22235 15113 22247 15116
rect 22189 15107 22247 15113
rect 17218 15076 17224 15088
rect 17179 15048 17224 15076
rect 17218 15036 17224 15048
rect 17276 15036 17282 15088
rect 22848 15076 22876 15116
rect 23750 15104 23756 15116
rect 23808 15104 23814 15156
rect 23845 15147 23903 15153
rect 23845 15113 23857 15147
rect 23891 15144 23903 15147
rect 24486 15144 24492 15156
rect 23891 15116 24492 15144
rect 23891 15113 23903 15116
rect 23845 15107 23903 15113
rect 24486 15104 24492 15116
rect 24544 15104 24550 15156
rect 24854 15144 24860 15156
rect 24815 15116 24860 15144
rect 24854 15104 24860 15116
rect 24912 15104 24918 15156
rect 26206 15116 40724 15144
rect 26206 15088 26234 15116
rect 22756 15048 22876 15076
rect 16945 15011 17003 15017
rect 16945 14977 16957 15011
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 18322 14968 18328 15020
rect 18380 14968 18386 15020
rect 20346 14968 20352 15020
rect 20404 15008 20410 15020
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 20404 14980 20453 15008
rect 20404 14968 20410 14980
rect 20441 14977 20453 14980
rect 20487 15008 20499 15011
rect 21085 15011 21143 15017
rect 21085 15008 21097 15011
rect 20487 14980 21097 15008
rect 20487 14977 20499 14980
rect 20441 14971 20499 14977
rect 21085 14977 21097 14980
rect 21131 14977 21143 15011
rect 22002 15008 22008 15020
rect 21963 14980 22008 15008
rect 21085 14971 21143 14977
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 22756 15017 22784 15048
rect 23382 15036 23388 15088
rect 23440 15076 23446 15088
rect 23661 15079 23719 15085
rect 23661 15076 23673 15079
rect 23440 15048 23673 15076
rect 23440 15036 23446 15048
rect 23661 15045 23673 15048
rect 23707 15045 23719 15079
rect 23661 15039 23719 15045
rect 23934 15036 23940 15088
rect 23992 15076 23998 15088
rect 25958 15076 25964 15088
rect 23992 15048 25964 15076
rect 23992 15036 23998 15048
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 22152 14980 22201 15008
rect 22152 14968 22158 14980
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 22741 15011 22799 15017
rect 22741 14977 22753 15011
rect 22787 14977 22799 15011
rect 22741 14971 22799 14977
rect 22833 15011 22891 15017
rect 22833 14977 22845 15011
rect 22879 15008 22891 15011
rect 23400 15008 23428 15036
rect 22879 14980 23428 15008
rect 22879 14977 22891 14980
rect 22833 14971 22891 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 13173 14943 13231 14949
rect 2832 14912 2877 14940
rect 2832 14900 2838 14912
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13814 14940 13820 14952
rect 13219 14912 13820 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 15102 14900 15108 14952
rect 15160 14940 15166 14952
rect 15197 14943 15255 14949
rect 15197 14940 15209 14943
rect 15160 14912 15209 14940
rect 15160 14900 15166 14912
rect 15197 14909 15209 14912
rect 15243 14940 15255 14943
rect 20254 14940 20260 14952
rect 15243 14912 20260 14940
rect 15243 14909 15255 14912
rect 15197 14903 15255 14909
rect 20254 14900 20260 14912
rect 20312 14900 20318 14952
rect 22204 14940 22232 14971
rect 23750 14968 23756 15020
rect 23808 15008 23814 15020
rect 24504 15017 24532 15048
rect 25958 15036 25964 15048
rect 26016 15036 26022 15088
rect 26142 15036 26148 15088
rect 26200 15048 26234 15088
rect 26200 15036 26206 15048
rect 24029 15011 24087 15017
rect 24029 15008 24041 15011
rect 23808 14980 24041 15008
rect 23808 14968 23814 14980
rect 24029 14977 24041 14980
rect 24075 14977 24087 15011
rect 24029 14971 24087 14977
rect 24489 15011 24547 15017
rect 24489 14977 24501 15011
rect 24535 14977 24547 15011
rect 24673 15011 24731 15017
rect 24673 15008 24685 15011
rect 24489 14971 24547 14977
rect 24596 14980 24685 15008
rect 24596 14940 24624 14980
rect 24673 14977 24685 14980
rect 24719 14977 24731 15011
rect 24673 14971 24731 14977
rect 22204 14912 24624 14940
rect 24688 14912 26234 14940
rect 23477 14875 23535 14881
rect 23477 14841 23489 14875
rect 23523 14872 23535 14875
rect 24688 14872 24716 14912
rect 23523 14844 24716 14872
rect 23523 14841 23535 14844
rect 23477 14835 23535 14841
rect 20533 14807 20591 14813
rect 20533 14773 20545 14807
rect 20579 14804 20591 14807
rect 20714 14804 20720 14816
rect 20579 14776 20720 14804
rect 20579 14773 20591 14776
rect 20533 14767 20591 14773
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 21174 14804 21180 14816
rect 21135 14776 21180 14804
rect 21174 14764 21180 14776
rect 21232 14764 21238 14816
rect 23014 14804 23020 14816
rect 22975 14776 23020 14804
rect 23014 14764 23020 14776
rect 23072 14764 23078 14816
rect 26206 14804 26234 14912
rect 40696 14872 40724 15116
rect 46198 15036 46204 15088
rect 46256 15076 46262 15088
rect 47762 15076 47768 15088
rect 46256 15048 47768 15076
rect 46256 15036 46262 15048
rect 47762 15036 47768 15048
rect 47820 15036 47826 15088
rect 45186 15008 45192 15020
rect 45147 14980 45192 15008
rect 45186 14968 45192 14980
rect 45244 14968 45250 15020
rect 47581 15011 47639 15017
rect 47581 14977 47593 15011
rect 47627 15008 47639 15011
rect 47670 15008 47676 15020
rect 47627 14980 47676 15008
rect 47627 14977 47639 14980
rect 47581 14971 47639 14977
rect 47670 14968 47676 14980
rect 47728 14968 47734 15020
rect 45373 14943 45431 14949
rect 45373 14909 45385 14943
rect 45419 14940 45431 14943
rect 45646 14940 45652 14952
rect 45419 14912 45652 14940
rect 45419 14909 45431 14912
rect 45373 14903 45431 14909
rect 45646 14900 45652 14912
rect 45704 14900 45710 14952
rect 45741 14943 45799 14949
rect 45741 14909 45753 14943
rect 45787 14909 45799 14943
rect 45741 14903 45799 14909
rect 45756 14872 45784 14903
rect 40696 14844 45784 14872
rect 46382 14804 46388 14816
rect 26206 14776 46388 14804
rect 46382 14764 46388 14776
rect 46440 14804 46446 14816
rect 46842 14804 46848 14816
rect 46440 14776 46848 14804
rect 46440 14764 46446 14776
rect 46842 14764 46848 14776
rect 46900 14764 46906 14816
rect 47946 14804 47952 14816
rect 47907 14776 47952 14804
rect 47946 14764 47952 14776
rect 48004 14764 48010 14816
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 16209 14603 16267 14609
rect 16209 14569 16221 14603
rect 16255 14569 16267 14603
rect 16390 14600 16396 14612
rect 16351 14572 16396 14600
rect 16209 14563 16267 14569
rect 16224 14532 16252 14563
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 17037 14603 17095 14609
rect 17037 14569 17049 14603
rect 17083 14600 17095 14603
rect 17126 14600 17132 14612
rect 17083 14572 17132 14600
rect 17083 14569 17095 14572
rect 17037 14563 17095 14569
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 22922 14600 22928 14612
rect 17236 14572 22928 14600
rect 16850 14532 16856 14544
rect 16224 14504 16856 14532
rect 16850 14492 16856 14504
rect 16908 14492 16914 14544
rect 17236 14532 17264 14572
rect 22922 14560 22928 14572
rect 22980 14560 22986 14612
rect 24486 14600 24492 14612
rect 24447 14572 24492 14600
rect 24486 14560 24492 14572
rect 24544 14560 24550 14612
rect 45646 14600 45652 14612
rect 45607 14572 45652 14600
rect 45646 14560 45652 14572
rect 45704 14560 45710 14612
rect 16960 14504 17264 14532
rect 3878 14424 3884 14476
rect 3936 14464 3942 14476
rect 16960 14464 16988 14504
rect 17402 14492 17408 14544
rect 17460 14532 17466 14544
rect 26142 14532 26148 14544
rect 17460 14504 26148 14532
rect 17460 14492 17466 14504
rect 26142 14492 26148 14504
rect 26200 14492 26206 14544
rect 46566 14492 46572 14544
rect 46624 14532 46630 14544
rect 46624 14504 47256 14532
rect 46624 14492 46630 14504
rect 3936 14436 16988 14464
rect 3936 14424 3942 14436
rect 17218 14424 17224 14476
rect 17276 14464 17282 14476
rect 21818 14464 21824 14476
rect 17276 14436 21680 14464
rect 21779 14436 21824 14464
rect 17276 14424 17282 14436
rect 2130 14396 2136 14408
rect 2091 14368 2136 14396
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14396 14151 14399
rect 14826 14396 14832 14408
rect 14139 14368 14832 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 14921 14399 14979 14405
rect 14921 14365 14933 14399
rect 14967 14396 14979 14399
rect 15010 14396 15016 14408
rect 14967 14368 15016 14396
rect 14967 14365 14979 14368
rect 14921 14359 14979 14365
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15197 14399 15255 14405
rect 15197 14365 15209 14399
rect 15243 14365 15255 14399
rect 15378 14396 15384 14408
rect 15339 14368 15384 14396
rect 15197 14359 15255 14365
rect 14185 14331 14243 14337
rect 14185 14297 14197 14331
rect 14231 14328 14243 14331
rect 14458 14328 14464 14340
rect 14231 14300 14464 14328
rect 14231 14297 14243 14300
rect 14185 14291 14243 14297
rect 14458 14288 14464 14300
rect 14516 14288 14522 14340
rect 15212 14328 15240 14359
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 15488 14390 16988 14396
rect 15488 14368 17172 14390
rect 15488 14328 15516 14368
rect 16960 14362 17172 14368
rect 15212 14300 15516 14328
rect 16025 14331 16083 14337
rect 16025 14297 16037 14331
rect 16071 14297 16083 14331
rect 16850 14328 16856 14340
rect 16811 14300 16856 14328
rect 16025 14291 16083 14297
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 14737 14263 14795 14269
rect 14737 14260 14749 14263
rect 14332 14232 14749 14260
rect 14332 14220 14338 14232
rect 14737 14229 14749 14232
rect 14783 14229 14795 14263
rect 14737 14223 14795 14229
rect 15378 14220 15384 14272
rect 15436 14260 15442 14272
rect 16040 14260 16068 14291
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 17144 14328 17172 14362
rect 19242 14356 19248 14408
rect 19300 14396 19306 14408
rect 19337 14399 19395 14405
rect 19337 14396 19349 14399
rect 19300 14368 19349 14396
rect 19300 14356 19306 14368
rect 19337 14365 19349 14368
rect 19383 14365 19395 14399
rect 20254 14396 20260 14408
rect 20215 14368 20260 14396
rect 19337 14359 19395 14365
rect 20254 14356 20260 14368
rect 20312 14356 20318 14408
rect 20441 14331 20499 14337
rect 17144 14300 17264 14328
rect 15436 14232 16068 14260
rect 16235 14263 16293 14269
rect 15436 14220 15442 14232
rect 16235 14229 16247 14263
rect 16281 14260 16293 14263
rect 16942 14260 16948 14272
rect 16281 14232 16948 14260
rect 16281 14229 16293 14232
rect 16235 14223 16293 14229
rect 16942 14220 16948 14232
rect 17000 14220 17006 14272
rect 17034 14220 17040 14272
rect 17092 14269 17098 14272
rect 17236 14269 17264 14300
rect 20441 14297 20453 14331
rect 20487 14297 20499 14331
rect 21652 14328 21680 14436
rect 21818 14424 21824 14436
rect 21876 14424 21882 14476
rect 22922 14424 22928 14476
rect 22980 14464 22986 14476
rect 23293 14467 23351 14473
rect 22980 14436 23152 14464
rect 22980 14424 22986 14436
rect 23014 14396 23020 14408
rect 22975 14368 23020 14396
rect 23014 14356 23020 14368
rect 23072 14356 23078 14408
rect 23124 14396 23152 14436
rect 23293 14433 23305 14467
rect 23339 14464 23351 14467
rect 25133 14467 25191 14473
rect 25133 14464 25145 14467
rect 23339 14436 25145 14464
rect 23339 14433 23351 14436
rect 23293 14427 23351 14433
rect 25133 14433 25145 14436
rect 25179 14433 25191 14467
rect 46658 14464 46664 14476
rect 46619 14436 46664 14464
rect 25133 14427 25191 14433
rect 46658 14424 46664 14436
rect 46716 14424 46722 14476
rect 47228 14473 47256 14504
rect 47762 14492 47768 14544
rect 47820 14492 47826 14544
rect 47213 14467 47271 14473
rect 47213 14433 47225 14467
rect 47259 14433 47271 14467
rect 47780 14464 47808 14492
rect 47780 14436 47992 14464
rect 47213 14427 47271 14433
rect 24397 14399 24455 14405
rect 24397 14396 24409 14399
rect 23124 14368 24409 14396
rect 24397 14365 24409 14368
rect 24443 14365 24455 14399
rect 24397 14359 24455 14365
rect 24581 14399 24639 14405
rect 24581 14365 24593 14399
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 25041 14399 25099 14405
rect 25041 14365 25053 14399
rect 25087 14365 25099 14399
rect 25222 14396 25228 14408
rect 25183 14368 25228 14396
rect 25041 14359 25099 14365
rect 22278 14328 22284 14340
rect 21652 14300 22284 14328
rect 20441 14291 20499 14297
rect 17092 14263 17111 14269
rect 17099 14229 17111 14263
rect 17092 14223 17111 14229
rect 17221 14263 17279 14269
rect 17221 14229 17233 14263
rect 17267 14229 17279 14263
rect 19426 14260 19432 14272
rect 19387 14232 19432 14260
rect 17221 14223 17279 14229
rect 17092 14220 17098 14223
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 20456 14260 20484 14291
rect 22278 14288 22284 14300
rect 22336 14288 22342 14340
rect 23750 14288 23756 14340
rect 23808 14328 23814 14340
rect 23808 14300 23980 14328
rect 23808 14288 23814 14300
rect 21174 14260 21180 14272
rect 20456 14232 21180 14260
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 23842 14260 23848 14272
rect 23803 14232 23848 14260
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 23952 14260 23980 14300
rect 24026 14288 24032 14340
rect 24084 14328 24090 14340
rect 24596 14328 24624 14359
rect 24084 14300 24624 14328
rect 24084 14288 24090 14300
rect 25056 14260 25084 14359
rect 25222 14356 25228 14368
rect 25280 14356 25286 14408
rect 45557 14399 45615 14405
rect 45557 14365 45569 14399
rect 45603 14365 45615 14399
rect 45557 14359 45615 14365
rect 45572 14328 45600 14359
rect 46290 14356 46296 14408
rect 46348 14396 46354 14408
rect 46477 14399 46535 14405
rect 46477 14396 46489 14399
rect 46348 14368 46489 14396
rect 46348 14356 46354 14368
rect 46477 14365 46489 14368
rect 46523 14365 46535 14399
rect 46477 14359 46535 14365
rect 47670 14356 47676 14408
rect 47728 14396 47734 14408
rect 47964 14405 47992 14436
rect 47765 14399 47823 14405
rect 47765 14396 47777 14399
rect 47728 14368 47777 14396
rect 47728 14356 47734 14368
rect 47765 14365 47777 14368
rect 47811 14365 47823 14399
rect 47765 14359 47823 14365
rect 47949 14399 48007 14405
rect 47949 14365 47961 14399
rect 47995 14365 48007 14399
rect 47949 14359 48007 14365
rect 47210 14328 47216 14340
rect 45572 14300 47216 14328
rect 47210 14288 47216 14300
rect 47268 14288 47274 14340
rect 47780 14328 47808 14359
rect 48222 14328 48228 14340
rect 47780 14300 48228 14328
rect 48222 14288 48228 14300
rect 48280 14288 48286 14340
rect 47854 14260 47860 14272
rect 23952 14232 25084 14260
rect 47815 14232 47860 14260
rect 47854 14220 47860 14232
rect 47912 14220 47918 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 2130 14016 2136 14068
rect 2188 14056 2194 14068
rect 17218 14056 17224 14068
rect 2188 14028 17224 14056
rect 2188 14016 2194 14028
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 19334 14056 19340 14068
rect 18432 14028 19340 14056
rect 14001 13991 14059 13997
rect 14001 13957 14013 13991
rect 14047 13988 14059 13991
rect 14274 13988 14280 14000
rect 14047 13960 14280 13988
rect 14047 13957 14059 13960
rect 14001 13951 14059 13957
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 14458 13948 14464 14000
rect 14516 13948 14522 14000
rect 16850 13948 16856 14000
rect 16908 13988 16914 14000
rect 17954 13988 17960 14000
rect 16908 13960 17960 13988
rect 16908 13948 16914 13960
rect 17954 13948 17960 13960
rect 18012 13948 18018 14000
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13630 13920 13636 13932
rect 13219 13892 13636 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 15930 13920 15936 13932
rect 15891 13892 15936 13920
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 16666 13880 16672 13932
rect 16724 13920 16730 13932
rect 16761 13923 16819 13929
rect 16761 13920 16773 13923
rect 16724 13892 16773 13920
rect 16724 13880 16730 13892
rect 16761 13889 16773 13892
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 16942 13880 16948 13932
rect 17000 13920 17006 13932
rect 18432 13929 18460 14028
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 23750 14056 23756 14068
rect 23711 14028 23756 14056
rect 23750 14016 23756 14028
rect 23808 14016 23814 14068
rect 24397 14059 24455 14065
rect 24397 14025 24409 14059
rect 24443 14056 24455 14059
rect 25222 14056 25228 14068
rect 24443 14028 25228 14056
rect 24443 14025 24455 14028
rect 24397 14019 24455 14025
rect 25222 14016 25228 14028
rect 25280 14016 25286 14068
rect 46385 14059 46443 14065
rect 46385 14025 46397 14059
rect 46431 14056 46443 14059
rect 47946 14056 47952 14068
rect 46431 14028 47952 14056
rect 46431 14025 46443 14028
rect 46385 14019 46443 14025
rect 47946 14016 47952 14028
rect 48004 14016 48010 14068
rect 19426 13948 19432 14000
rect 19484 13948 19490 14000
rect 46474 13948 46480 14000
rect 46532 13988 46538 14000
rect 47673 13991 47731 13997
rect 47673 13988 47685 13991
rect 46532 13960 47685 13988
rect 46532 13948 46538 13960
rect 47673 13957 47685 13960
rect 47719 13957 47731 13991
rect 47673 13951 47731 13957
rect 17589 13923 17647 13929
rect 17589 13920 17601 13923
rect 17000 13892 17601 13920
rect 17000 13880 17006 13892
rect 17589 13889 17601 13892
rect 17635 13920 17647 13923
rect 18417 13923 18475 13929
rect 17635 13892 17908 13920
rect 17635 13889 17647 13892
rect 17589 13883 17647 13889
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13852 13323 13855
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 13311 13824 13737 13852
rect 13311 13821 13323 13824
rect 13265 13815 13323 13821
rect 13725 13821 13737 13824
rect 13771 13821 13783 13855
rect 15470 13852 15476 13864
rect 15431 13824 15476 13852
rect 13725 13815 13783 13821
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 16684 13784 16712 13880
rect 16850 13852 16856 13864
rect 16811 13824 16856 13852
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 17034 13852 17040 13864
rect 16960 13824 17040 13852
rect 16960 13784 16988 13824
rect 17034 13812 17040 13824
rect 17092 13852 17098 13864
rect 17497 13855 17555 13861
rect 17497 13852 17509 13855
rect 17092 13824 17509 13852
rect 17092 13812 17098 13824
rect 17497 13821 17509 13824
rect 17543 13821 17555 13855
rect 17497 13815 17555 13821
rect 16684 13756 16988 13784
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 13814 13716 13820 13728
rect 4028 13688 13820 13716
rect 4028 13676 4034 13688
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 16022 13716 16028 13728
rect 15983 13688 16028 13716
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 17880 13716 17908 13892
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 22922 13880 22928 13932
rect 22980 13920 22986 13932
rect 23661 13923 23719 13929
rect 23661 13920 23673 13923
rect 22980 13892 23673 13920
rect 22980 13880 22986 13892
rect 23661 13889 23673 13892
rect 23707 13889 23719 13923
rect 23661 13883 23719 13889
rect 23845 13923 23903 13929
rect 23845 13889 23857 13923
rect 23891 13920 23903 13923
rect 24026 13920 24032 13932
rect 23891 13892 24032 13920
rect 23891 13889 23903 13892
rect 23845 13883 23903 13889
rect 24026 13880 24032 13892
rect 24084 13880 24090 13932
rect 24305 13923 24363 13929
rect 24305 13889 24317 13923
rect 24351 13920 24363 13923
rect 24486 13920 24492 13932
rect 24351 13892 24492 13920
rect 24351 13889 24363 13892
rect 24305 13883 24363 13889
rect 24486 13880 24492 13892
rect 24544 13880 24550 13932
rect 46290 13880 46296 13932
rect 46348 13920 46354 13932
rect 47029 13923 47087 13929
rect 47029 13920 47041 13923
rect 46348 13892 47041 13920
rect 46348 13880 46354 13892
rect 47029 13889 47041 13892
rect 47075 13889 47087 13923
rect 47029 13883 47087 13889
rect 47210 13880 47216 13932
rect 47268 13920 47274 13932
rect 47581 13923 47639 13929
rect 47581 13920 47593 13923
rect 47268 13892 47593 13920
rect 47268 13880 47274 13892
rect 47581 13889 47593 13892
rect 47627 13889 47639 13923
rect 47581 13883 47639 13889
rect 18693 13855 18751 13861
rect 18693 13852 18705 13855
rect 18524 13824 18705 13852
rect 17957 13787 18015 13793
rect 17957 13753 17969 13787
rect 18003 13784 18015 13787
rect 18524 13784 18552 13824
rect 18693 13821 18705 13824
rect 18739 13821 18751 13855
rect 18693 13815 18751 13821
rect 22278 13812 22284 13864
rect 22336 13852 22342 13864
rect 22830 13852 22836 13864
rect 22336 13824 22836 13852
rect 22336 13812 22342 13824
rect 22830 13812 22836 13824
rect 22888 13812 22894 13864
rect 46753 13855 46811 13861
rect 46753 13821 46765 13855
rect 46799 13821 46811 13855
rect 46753 13815 46811 13821
rect 18003 13756 18552 13784
rect 46768 13784 46796 13815
rect 46842 13812 46848 13864
rect 46900 13852 46906 13864
rect 47854 13852 47860 13864
rect 46900 13824 46945 13852
rect 47044 13824 47860 13852
rect 46900 13812 46906 13824
rect 47044 13784 47072 13824
rect 47854 13812 47860 13824
rect 47912 13812 47918 13864
rect 46768 13756 47072 13784
rect 18003 13753 18015 13756
rect 17957 13747 18015 13753
rect 20162 13716 20168 13728
rect 17880 13688 20168 13716
rect 20162 13676 20168 13688
rect 20220 13676 20226 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19392 13484 19441 13512
rect 19392 13472 19398 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 46658 13512 46664 13524
rect 46619 13484 46664 13512
rect 19429 13475 19487 13481
rect 46658 13472 46664 13484
rect 46716 13472 46722 13524
rect 12434 13404 12440 13456
rect 12492 13444 12498 13456
rect 12492 13416 16160 13444
rect 12492 13404 12498 13416
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 16022 13376 16028 13388
rect 15335 13348 16028 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16132 13385 16160 13416
rect 19242 13404 19248 13456
rect 19300 13404 19306 13456
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13345 16175 13379
rect 19260 13376 19288 13404
rect 16117 13339 16175 13345
rect 18432 13348 19288 13376
rect 18432 13317 18460 13348
rect 20162 13336 20168 13388
rect 20220 13376 20226 13388
rect 20533 13379 20591 13385
rect 20533 13376 20545 13379
rect 20220 13348 20545 13376
rect 20220 13336 20226 13348
rect 20533 13345 20545 13348
rect 20579 13345 20591 13379
rect 20714 13376 20720 13388
rect 20675 13348 20720 13376
rect 20533 13339 20591 13345
rect 20714 13336 20720 13348
rect 20772 13336 20778 13388
rect 45370 13336 45376 13388
rect 45428 13376 45434 13388
rect 45833 13379 45891 13385
rect 45833 13376 45845 13379
rect 45428 13348 45845 13376
rect 45428 13336 45434 13348
rect 45833 13345 45845 13348
rect 45879 13376 45891 13379
rect 47210 13376 47216 13388
rect 45879 13348 47216 13376
rect 45879 13345 45891 13348
rect 45833 13339 45891 13345
rect 47210 13336 47216 13348
rect 47268 13336 47274 13388
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13277 15163 13311
rect 15105 13271 15163 13277
rect 17589 13311 17647 13317
rect 17589 13277 17601 13311
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 18417 13311 18475 13317
rect 18417 13277 18429 13311
rect 18463 13277 18475 13311
rect 18417 13271 18475 13277
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13308 19487 13311
rect 19978 13308 19984 13320
rect 19475 13280 19984 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 15120 13240 15148 13271
rect 15470 13240 15476 13252
rect 15120 13212 15476 13240
rect 15470 13200 15476 13212
rect 15528 13200 15534 13252
rect 17604 13240 17632 13271
rect 19444 13240 19472 13271
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 46017 13311 46075 13317
rect 46017 13277 46029 13311
rect 46063 13277 46075 13311
rect 46017 13271 46075 13277
rect 17604 13212 19472 13240
rect 22373 13243 22431 13249
rect 22373 13209 22385 13243
rect 22419 13240 22431 13243
rect 30466 13240 30472 13252
rect 22419 13212 30472 13240
rect 22419 13209 22431 13212
rect 22373 13203 22431 13209
rect 30466 13200 30472 13212
rect 30524 13200 30530 13252
rect 45186 13200 45192 13252
rect 45244 13240 45250 13252
rect 46032 13240 46060 13271
rect 46106 13268 46112 13320
rect 46164 13308 46170 13320
rect 46661 13311 46719 13317
rect 46661 13308 46673 13311
rect 46164 13280 46673 13308
rect 46164 13268 46170 13280
rect 46661 13277 46673 13280
rect 46707 13277 46719 13311
rect 46661 13271 46719 13277
rect 46845 13311 46903 13317
rect 46845 13277 46857 13311
rect 46891 13277 46903 13311
rect 47670 13308 47676 13320
rect 47631 13280 47676 13308
rect 46845 13271 46903 13277
rect 45244 13212 46060 13240
rect 46201 13243 46259 13249
rect 45244 13200 45250 13212
rect 46201 13209 46213 13243
rect 46247 13240 46259 13243
rect 46860 13240 46888 13271
rect 47670 13268 47676 13280
rect 47728 13268 47734 13320
rect 46247 13212 46888 13240
rect 46247 13209 46259 13212
rect 46201 13203 46259 13209
rect 17126 13132 17132 13184
rect 17184 13172 17190 13184
rect 17589 13175 17647 13181
rect 17589 13172 17601 13175
rect 17184 13144 17601 13172
rect 17184 13132 17190 13144
rect 17589 13141 17601 13144
rect 17635 13141 17647 13175
rect 18506 13172 18512 13184
rect 18467 13144 18512 13172
rect 17589 13135 17647 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 23477 12903 23535 12909
rect 23477 12869 23489 12903
rect 23523 12900 23535 12903
rect 24213 12903 24271 12909
rect 24213 12900 24225 12903
rect 23523 12872 24225 12900
rect 23523 12869 23535 12872
rect 23477 12863 23535 12869
rect 24213 12869 24225 12872
rect 24259 12869 24271 12903
rect 24213 12863 24271 12869
rect 45281 12903 45339 12909
rect 45281 12869 45293 12903
rect 45327 12900 45339 12903
rect 46201 12903 46259 12909
rect 45327 12872 46060 12900
rect 45327 12869 45339 12872
rect 45281 12863 45339 12869
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 17126 12832 17132 12844
rect 17087 12804 17132 12832
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 18506 12792 18512 12844
rect 18564 12792 18570 12844
rect 21542 12792 21548 12844
rect 21600 12832 21606 12844
rect 21726 12832 21732 12844
rect 21600 12804 21732 12832
rect 21600 12792 21606 12804
rect 21726 12792 21732 12804
rect 21784 12832 21790 12844
rect 23385 12835 23443 12841
rect 23385 12832 23397 12835
rect 21784 12804 23397 12832
rect 21784 12792 21790 12804
rect 23385 12801 23397 12804
rect 23431 12801 23443 12835
rect 23385 12795 23443 12801
rect 23842 12792 23848 12844
rect 23900 12832 23906 12844
rect 24029 12835 24087 12841
rect 24029 12832 24041 12835
rect 23900 12804 24041 12832
rect 23900 12792 23906 12804
rect 24029 12801 24041 12804
rect 24075 12801 24087 12835
rect 45186 12832 45192 12844
rect 45147 12804 45192 12832
rect 24029 12795 24087 12801
rect 45186 12792 45192 12804
rect 45244 12792 45250 12844
rect 45370 12832 45376 12844
rect 45331 12804 45376 12832
rect 45370 12792 45376 12804
rect 45428 12792 45434 12844
rect 46032 12841 46060 12872
rect 46201 12869 46213 12903
rect 46247 12900 46259 12903
rect 46845 12903 46903 12909
rect 46845 12900 46857 12903
rect 46247 12872 46857 12900
rect 46247 12869 46259 12872
rect 46201 12863 46259 12869
rect 46845 12869 46857 12872
rect 46891 12869 46903 12903
rect 46845 12863 46903 12869
rect 46017 12835 46075 12841
rect 46017 12801 46029 12835
rect 46063 12832 46075 12835
rect 46106 12832 46112 12844
rect 46063 12804 46112 12832
rect 46063 12801 46075 12804
rect 46017 12795 46075 12801
rect 46106 12792 46112 12804
rect 46164 12792 46170 12844
rect 46290 12832 46296 12844
rect 46251 12804 46296 12832
rect 46290 12792 46296 12804
rect 46348 12792 46354 12844
rect 46753 12835 46811 12841
rect 46753 12801 46765 12835
rect 46799 12801 46811 12835
rect 46753 12795 46811 12801
rect 46937 12835 46995 12841
rect 46937 12801 46949 12835
rect 46983 12832 46995 12835
rect 47210 12832 47216 12844
rect 46983 12804 47216 12832
rect 46983 12801 46995 12804
rect 46937 12795 46995 12801
rect 17034 12724 17040 12776
rect 17092 12764 17098 12776
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 17092 12736 17417 12764
rect 17092 12724 17098 12736
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 25866 12764 25872 12776
rect 25827 12736 25872 12764
rect 17405 12727 17463 12733
rect 25866 12724 25872 12736
rect 25924 12724 25930 12776
rect 45204 12764 45232 12792
rect 46768 12764 46796 12795
rect 47210 12792 47216 12804
rect 47268 12792 47274 12844
rect 45204 12736 46796 12764
rect 25038 12696 25044 12708
rect 18432 12668 25044 12696
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 18432 12628 18460 12668
rect 25038 12656 25044 12668
rect 25096 12656 25102 12708
rect 18874 12628 18880 12640
rect 1627 12600 18460 12628
rect 18835 12600 18880 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 45830 12628 45836 12640
rect 45791 12600 45836 12628
rect 45830 12588 45836 12600
rect 45888 12588 45894 12640
rect 46014 12588 46020 12640
rect 46072 12628 46078 12640
rect 46198 12628 46204 12640
rect 46072 12600 46204 12628
rect 46072 12588 46078 12600
rect 46198 12588 46204 12600
rect 46256 12588 46262 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 45373 12427 45431 12433
rect 45373 12393 45385 12427
rect 45419 12424 45431 12427
rect 45738 12424 45744 12436
rect 45419 12396 45744 12424
rect 45419 12393 45431 12396
rect 45373 12387 45431 12393
rect 45738 12384 45744 12396
rect 45796 12384 45802 12436
rect 17034 12356 17040 12368
rect 16995 12328 17040 12356
rect 17034 12316 17040 12328
rect 17092 12316 17098 12368
rect 47670 12356 47676 12368
rect 46308 12328 47676 12356
rect 16761 12291 16819 12297
rect 16761 12257 16773 12291
rect 16807 12288 16819 12291
rect 16850 12288 16856 12300
rect 16807 12260 16856 12288
rect 16807 12257 16819 12260
rect 16761 12251 16819 12257
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 45738 12288 45744 12300
rect 45699 12260 45744 12288
rect 45738 12248 45744 12260
rect 45796 12248 45802 12300
rect 46308 12297 46336 12328
rect 47670 12316 47676 12328
rect 47728 12316 47734 12368
rect 46293 12291 46351 12297
rect 46293 12257 46305 12291
rect 46339 12257 46351 12291
rect 46474 12288 46480 12300
rect 46435 12260 46480 12288
rect 46293 12251 46351 12257
rect 46474 12248 46480 12260
rect 46532 12248 46538 12300
rect 48130 12288 48136 12300
rect 48091 12260 48136 12288
rect 48130 12248 48136 12260
rect 48188 12248 48194 12300
rect 15010 12180 15016 12232
rect 15068 12220 15074 12232
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 15068 12192 16681 12220
rect 15068 12180 15074 12192
rect 16669 12189 16681 12192
rect 16715 12220 16727 12223
rect 17954 12220 17960 12232
rect 16715 12192 17960 12220
rect 16715 12189 16727 12192
rect 16669 12183 16727 12189
rect 17954 12180 17960 12192
rect 18012 12220 18018 12232
rect 18874 12220 18880 12232
rect 18012 12192 18880 12220
rect 18012 12180 18018 12192
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 45557 12223 45615 12229
rect 45557 12189 45569 12223
rect 45603 12220 45615 12223
rect 45646 12220 45652 12232
rect 45603 12192 45652 12220
rect 45603 12189 45615 12192
rect 45557 12183 45615 12189
rect 45646 12180 45652 12192
rect 45704 12180 45710 12232
rect 45833 12223 45891 12229
rect 45833 12189 45845 12223
rect 45879 12220 45891 12223
rect 45879 12192 45968 12220
rect 45879 12189 45891 12192
rect 45833 12183 45891 12189
rect 45370 12112 45376 12164
rect 45428 12152 45434 12164
rect 45940 12152 45968 12192
rect 45428 12124 45968 12152
rect 45428 12112 45434 12124
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 15105 11747 15163 11753
rect 15105 11713 15117 11747
rect 15151 11744 15163 11747
rect 15654 11744 15660 11756
rect 15151 11716 15660 11744
rect 15151 11713 15163 11716
rect 15105 11707 15163 11713
rect 15654 11704 15660 11716
rect 15712 11744 15718 11756
rect 21358 11744 21364 11756
rect 15712 11716 21364 11744
rect 15712 11704 15718 11716
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 45738 11744 45744 11756
rect 45699 11716 45744 11744
rect 45738 11704 45744 11716
rect 45796 11704 45802 11756
rect 45830 11704 45836 11756
rect 45888 11744 45894 11756
rect 46201 11747 46259 11753
rect 46201 11744 46213 11747
rect 45888 11716 46213 11744
rect 45888 11704 45894 11716
rect 46201 11713 46213 11716
rect 46247 11713 46259 11747
rect 46201 11707 46259 11713
rect 45554 11568 45560 11620
rect 45612 11608 45618 11620
rect 46385 11611 46443 11617
rect 46385 11608 46397 11611
rect 45612 11580 46397 11608
rect 45612 11568 45618 11580
rect 46385 11577 46397 11580
rect 46431 11608 46443 11611
rect 46750 11608 46756 11620
rect 46431 11580 46756 11608
rect 46431 11577 46443 11580
rect 46385 11571 46443 11577
rect 46750 11568 46756 11580
rect 46808 11568 46814 11620
rect 15194 11540 15200 11552
rect 15155 11512 15200 11540
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 47762 11540 47768 11552
rect 47723 11512 47768 11540
rect 47762 11500 47768 11512
rect 47820 11500 47826 11552
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 3326 11296 3332 11348
rect 3384 11336 3390 11348
rect 3384 11308 12434 11336
rect 3384 11296 3390 11308
rect 12406 11064 12434 11308
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 14884 11308 15424 11336
rect 14884 11296 14890 11308
rect 15010 11200 15016 11212
rect 14971 11172 15016 11200
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 15194 11200 15200 11212
rect 15155 11172 15200 11200
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 15396 11200 15424 11308
rect 21726 11296 21732 11348
rect 21784 11336 21790 11348
rect 45554 11336 45560 11348
rect 21784 11308 45560 11336
rect 21784 11296 21790 11308
rect 45554 11296 45560 11308
rect 45612 11296 45618 11348
rect 45830 11336 45836 11348
rect 45791 11308 45836 11336
rect 45830 11296 45836 11308
rect 45888 11296 45894 11348
rect 45646 11268 45652 11280
rect 21652 11240 22232 11268
rect 45607 11240 45652 11268
rect 15473 11203 15531 11209
rect 15473 11200 15485 11203
rect 15396 11172 15485 11200
rect 15473 11169 15485 11172
rect 15519 11169 15531 11203
rect 21652 11200 21680 11240
rect 22204 11209 22232 11240
rect 45646 11228 45652 11240
rect 45704 11228 45710 11280
rect 15473 11163 15531 11169
rect 16408 11172 21680 11200
rect 22189 11203 22247 11209
rect 16408 11064 16436 11172
rect 22189 11169 22201 11203
rect 22235 11169 22247 11203
rect 45370 11200 45376 11212
rect 45331 11172 45376 11200
rect 22189 11163 22247 11169
rect 45370 11160 45376 11172
rect 45428 11160 45434 11212
rect 46293 11203 46351 11209
rect 46293 11169 46305 11203
rect 46339 11200 46351 11203
rect 47762 11200 47768 11212
rect 46339 11172 47768 11200
rect 46339 11169 46351 11172
rect 46293 11163 46351 11169
rect 47762 11160 47768 11172
rect 47820 11160 47826 11212
rect 21726 11132 21732 11144
rect 21687 11104 21732 11132
rect 21726 11092 21732 11104
rect 21784 11092 21790 11144
rect 21910 11064 21916 11076
rect 12406 11036 16436 11064
rect 21871 11036 21916 11064
rect 21910 11024 21916 11036
rect 21968 11024 21974 11076
rect 46014 11024 46020 11076
rect 46072 11064 46078 11076
rect 46477 11067 46535 11073
rect 46477 11064 46489 11067
rect 46072 11036 46489 11064
rect 46072 11024 46078 11036
rect 46477 11033 46489 11036
rect 46523 11033 46535 11067
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 46477 11027 46535 11033
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 21910 10792 21916 10804
rect 21871 10764 21916 10792
rect 21910 10752 21916 10764
rect 21968 10752 21974 10804
rect 45370 10792 45376 10804
rect 45331 10764 45376 10792
rect 45370 10752 45376 10764
rect 45428 10752 45434 10804
rect 46106 10724 46112 10736
rect 46067 10696 46112 10724
rect 46106 10684 46112 10696
rect 46164 10684 46170 10736
rect 21634 10616 21640 10668
rect 21692 10656 21698 10668
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 21692 10628 21833 10656
rect 21692 10616 21698 10628
rect 21821 10625 21833 10628
rect 21867 10625 21879 10659
rect 21821 10619 21879 10625
rect 45281 10659 45339 10665
rect 45281 10625 45293 10659
rect 45327 10625 45339 10659
rect 45462 10656 45468 10668
rect 45423 10628 45468 10656
rect 45281 10619 45339 10625
rect 45296 10520 45324 10619
rect 45462 10616 45468 10628
rect 45520 10616 45526 10668
rect 45370 10548 45376 10600
rect 45428 10588 45434 10600
rect 46017 10591 46075 10597
rect 46017 10588 46029 10591
rect 45428 10560 46029 10588
rect 45428 10548 45434 10560
rect 46017 10557 46029 10560
rect 46063 10557 46075 10591
rect 46017 10551 46075 10557
rect 46198 10548 46204 10600
rect 46256 10588 46262 10600
rect 46293 10591 46351 10597
rect 46293 10588 46305 10591
rect 46256 10560 46305 10588
rect 46256 10548 46262 10560
rect 46293 10557 46305 10560
rect 46339 10557 46351 10591
rect 46293 10551 46351 10557
rect 45554 10520 45560 10532
rect 45296 10492 45560 10520
rect 45554 10480 45560 10492
rect 45612 10520 45618 10532
rect 46216 10520 46244 10548
rect 45612 10492 46244 10520
rect 45612 10480 45618 10492
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 9214 10452 9220 10464
rect 3568 10424 9220 10452
rect 3568 10412 3574 10424
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 46290 10412 46296 10464
rect 46348 10452 46354 10464
rect 47765 10455 47823 10461
rect 47765 10452 47777 10455
rect 46348 10424 47777 10452
rect 46348 10412 46354 10424
rect 47765 10421 47777 10424
rect 47811 10421 47823 10455
rect 47765 10415 47823 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 45646 10248 45652 10260
rect 45607 10220 45652 10248
rect 45646 10208 45652 10220
rect 45704 10208 45710 10260
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 45554 10044 45560 10056
rect 45515 10016 45560 10044
rect 45554 10004 45560 10016
rect 45612 10004 45618 10056
rect 45741 10047 45799 10053
rect 45741 10013 45753 10047
rect 45787 10013 45799 10047
rect 45741 10007 45799 10013
rect 45094 9936 45100 9988
rect 45152 9976 45158 9988
rect 45462 9976 45468 9988
rect 45152 9948 45468 9976
rect 45152 9936 45158 9948
rect 45462 9936 45468 9948
rect 45520 9976 45526 9988
rect 45756 9976 45784 10007
rect 45520 9948 45784 9976
rect 46477 9979 46535 9985
rect 45520 9936 45526 9948
rect 46477 9945 46489 9979
rect 46523 9976 46535 9979
rect 47670 9976 47676 9988
rect 46523 9948 47676 9976
rect 46523 9945 46535 9948
rect 46477 9939 46535 9945
rect 47670 9936 47676 9948
rect 47728 9936 47734 9988
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 46106 9664 46112 9716
rect 46164 9704 46170 9716
rect 46845 9707 46903 9713
rect 46845 9704 46857 9707
rect 46164 9676 46857 9704
rect 46164 9664 46170 9676
rect 46845 9673 46857 9676
rect 46891 9673 46903 9707
rect 46845 9667 46903 9673
rect 47670 9636 47676 9648
rect 47631 9608 47676 9636
rect 47670 9596 47676 9608
rect 47728 9596 47734 9648
rect 46842 9528 46848 9580
rect 46900 9568 46906 9580
rect 47029 9571 47087 9577
rect 47029 9568 47041 9571
rect 46900 9540 47041 9568
rect 46900 9528 46906 9540
rect 47029 9537 47041 9540
rect 47075 9537 47087 9571
rect 47029 9531 47087 9537
rect 47486 9528 47492 9580
rect 47544 9568 47550 9580
rect 47581 9571 47639 9577
rect 47581 9568 47593 9571
rect 47544 9540 47593 9568
rect 47544 9528 47550 9540
rect 47581 9537 47593 9540
rect 47627 9537 47639 9571
rect 47581 9531 47639 9537
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 9024 16359 9027
rect 16574 9024 16580 9036
rect 16347 8996 16580 9024
rect 16347 8993 16359 8996
rect 16301 8987 16359 8993
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 16666 8984 16672 9036
rect 16724 9024 16730 9036
rect 16761 9027 16819 9033
rect 16761 9024 16773 9027
rect 16724 8996 16773 9024
rect 16724 8984 16730 8996
rect 16761 8993 16773 8996
rect 16807 8993 16819 9027
rect 16761 8987 16819 8993
rect 15654 8956 15660 8968
rect 15615 8928 15660 8956
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 47302 8956 47308 8968
rect 47263 8928 47308 8956
rect 47302 8916 47308 8928
rect 47360 8916 47366 8968
rect 47394 8916 47400 8968
rect 47452 8956 47458 8968
rect 47581 8959 47639 8965
rect 47581 8956 47593 8959
rect 47452 8928 47593 8956
rect 47452 8916 47458 8928
rect 47581 8925 47593 8928
rect 47627 8925 47639 8959
rect 47581 8919 47639 8925
rect 15749 8891 15807 8897
rect 15749 8857 15761 8891
rect 15795 8888 15807 8891
rect 16485 8891 16543 8897
rect 16485 8888 16497 8891
rect 15795 8860 16497 8888
rect 15795 8857 15807 8860
rect 15749 8851 15807 8857
rect 16485 8857 16497 8860
rect 16531 8857 16543 8891
rect 16485 8851 16543 8857
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 47762 8548 47768 8560
rect 47723 8520 47768 8548
rect 47762 8508 47768 8520
rect 47820 8508 47826 8560
rect 24946 8304 24952 8356
rect 25004 8344 25010 8356
rect 47949 8347 48007 8353
rect 47949 8344 47961 8347
rect 25004 8316 47961 8344
rect 25004 8304 25010 8316
rect 47949 8313 47961 8316
rect 47995 8313 48007 8347
rect 47949 8307 48007 8313
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 12434 8276 12440 8288
rect 3016 8248 12440 8276
rect 3016 8236 3022 8248
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 21818 8236 21824 8288
rect 21876 8276 21882 8288
rect 45554 8276 45560 8288
rect 21876 8248 45560 8276
rect 21876 8236 21882 8248
rect 45554 8236 45560 8248
rect 45612 8236 45618 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 30926 7964 30932 8016
rect 30984 8004 30990 8016
rect 33870 8004 33876 8016
rect 30984 7976 33876 8004
rect 30984 7964 30990 7976
rect 33870 7964 33876 7976
rect 33928 7964 33934 8016
rect 47118 8004 47124 8016
rect 46308 7976 47124 8004
rect 46308 7945 46336 7976
rect 47118 7964 47124 7976
rect 47176 7964 47182 8016
rect 46293 7939 46351 7945
rect 46293 7905 46305 7939
rect 46339 7905 46351 7939
rect 46293 7899 46351 7905
rect 46477 7939 46535 7945
rect 46477 7905 46489 7939
rect 46523 7936 46535 7939
rect 47394 7936 47400 7948
rect 46523 7908 47400 7936
rect 46523 7905 46535 7908
rect 46477 7899 46535 7905
rect 47394 7896 47400 7908
rect 47452 7896 47458 7948
rect 47670 7936 47676 7948
rect 47631 7908 47676 7936
rect 47670 7896 47676 7908
rect 47728 7896 47734 7948
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 48130 7392 48136 7404
rect 48091 7364 48136 7392
rect 48130 7352 48136 7364
rect 48188 7352 48194 7404
rect 47118 7148 47124 7200
rect 47176 7188 47182 7200
rect 47949 7191 48007 7197
rect 47949 7188 47961 7191
rect 47176 7160 47961 7188
rect 47176 7148 47182 7160
rect 47949 7157 47961 7160
rect 47995 7157 48007 7191
rect 47949 7151 48007 7157
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 17770 6848 17776 6860
rect 3568 6820 17776 6848
rect 3568 6808 3574 6820
rect 17770 6808 17776 6820
rect 17828 6808 17834 6860
rect 47118 6848 47124 6860
rect 47079 6820 47124 6848
rect 47118 6808 47124 6820
rect 47176 6808 47182 6860
rect 48133 6851 48191 6857
rect 48133 6817 48145 6851
rect 48179 6848 48191 6851
rect 48222 6848 48228 6860
rect 48179 6820 48228 6848
rect 48179 6817 48191 6820
rect 48133 6811 48191 6817
rect 48222 6808 48228 6820
rect 48280 6808 48286 6860
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6780 7619 6783
rect 22370 6780 22376 6792
rect 7607 6752 22376 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 22370 6740 22376 6752
rect 22428 6740 22434 6792
rect 1670 6672 1676 6724
rect 1728 6712 1734 6724
rect 47213 6715 47271 6721
rect 47213 6712 47225 6715
rect 1728 6684 26234 6712
rect 1728 6672 1734 6684
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7653 6647 7711 6653
rect 7653 6644 7665 6647
rect 6972 6616 7665 6644
rect 6972 6604 6978 6616
rect 7653 6613 7665 6616
rect 7699 6613 7711 6647
rect 26206 6644 26234 6684
rect 41386 6684 47225 6712
rect 41386 6644 41414 6684
rect 47213 6681 47225 6684
rect 47259 6681 47271 6715
rect 47213 6675 47271 6681
rect 26206 6616 41414 6644
rect 7653 6607 7711 6613
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 6914 6332 6920 6384
rect 6972 6372 6978 6384
rect 6972 6344 7017 6372
rect 6972 6332 6978 6344
rect 6733 6239 6791 6245
rect 6733 6205 6745 6239
rect 6779 6236 6791 6239
rect 6914 6236 6920 6248
rect 6779 6208 6920 6236
rect 6779 6205 6791 6208
rect 6733 6199 6791 6205
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7193 6239 7251 6245
rect 7193 6205 7205 6239
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 6454 6128 6460 6180
rect 6512 6168 6518 6180
rect 7208 6168 7236 6199
rect 6512 6140 7236 6168
rect 6512 6128 6518 6140
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 6972 5868 7017 5896
rect 6972 5856 6978 5868
rect 46842 5720 46848 5772
rect 46900 5760 46906 5772
rect 47305 5763 47363 5769
rect 47305 5760 47317 5763
rect 46900 5732 47317 5760
rect 46900 5720 46906 5732
rect 47305 5729 47317 5732
rect 47351 5729 47363 5763
rect 47305 5723 47363 5729
rect 21082 5652 21088 5704
rect 21140 5692 21146 5704
rect 22189 5695 22247 5701
rect 22189 5692 22201 5695
rect 21140 5664 22201 5692
rect 21140 5652 21146 5664
rect 22189 5661 22201 5664
rect 22235 5661 22247 5695
rect 22189 5655 22247 5661
rect 47210 5652 47216 5704
rect 47268 5692 47274 5704
rect 47581 5695 47639 5701
rect 47581 5692 47593 5695
rect 47268 5664 47593 5692
rect 47268 5652 47274 5664
rect 47581 5661 47593 5664
rect 47627 5661 47639 5695
rect 47581 5655 47639 5661
rect 20622 5516 20628 5568
rect 20680 5556 20686 5568
rect 22281 5559 22339 5565
rect 22281 5556 22293 5559
rect 20680 5528 22293 5556
rect 20680 5516 20686 5528
rect 22281 5525 22293 5528
rect 22327 5525 22339 5559
rect 22281 5519 22339 5525
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 18874 5216 18880 5228
rect 18835 5188 18880 5216
rect 18874 5176 18880 5188
rect 18932 5176 18938 5228
rect 19889 5219 19947 5225
rect 19889 5185 19901 5219
rect 19935 5216 19947 5219
rect 20806 5216 20812 5228
rect 19935 5188 20812 5216
rect 19935 5185 19947 5188
rect 19889 5179 19947 5185
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 21821 5219 21879 5225
rect 21821 5185 21833 5219
rect 21867 5216 21879 5219
rect 22370 5216 22376 5228
rect 21867 5188 22376 5216
rect 21867 5185 21879 5188
rect 21821 5179 21879 5185
rect 22370 5176 22376 5188
rect 22428 5176 22434 5228
rect 22465 5219 22523 5225
rect 22465 5185 22477 5219
rect 22511 5216 22523 5219
rect 22738 5216 22744 5228
rect 22511 5188 22744 5216
rect 22511 5185 22523 5188
rect 22465 5179 22523 5185
rect 22738 5176 22744 5188
rect 22796 5176 22802 5228
rect 23474 5216 23480 5228
rect 23435 5188 23480 5216
rect 23474 5176 23480 5188
rect 23532 5176 23538 5228
rect 46842 5176 46848 5228
rect 46900 5216 46906 5228
rect 47029 5219 47087 5225
rect 47029 5216 47041 5219
rect 46900 5188 47041 5216
rect 46900 5176 46906 5188
rect 47029 5185 47041 5188
rect 47075 5185 47087 5219
rect 47029 5179 47087 5185
rect 47857 5219 47915 5225
rect 47857 5185 47869 5219
rect 47903 5216 47915 5219
rect 48314 5216 48320 5228
rect 47903 5188 48320 5216
rect 47903 5185 47915 5188
rect 47857 5179 47915 5185
rect 48314 5176 48320 5188
rect 48372 5176 48378 5228
rect 44726 5040 44732 5092
rect 44784 5080 44790 5092
rect 44784 5052 48084 5080
rect 44784 5040 44790 5052
rect 18598 4972 18604 5024
rect 18656 5012 18662 5024
rect 18969 5015 19027 5021
rect 18969 5012 18981 5015
rect 18656 4984 18981 5012
rect 18656 4972 18662 4984
rect 18969 4981 18981 4984
rect 19015 4981 19027 5015
rect 18969 4975 19027 4981
rect 19981 5015 20039 5021
rect 19981 4981 19993 5015
rect 20027 5012 20039 5015
rect 21358 5012 21364 5024
rect 20027 4984 21364 5012
rect 20027 4981 20039 4984
rect 19981 4975 20039 4981
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 21913 5015 21971 5021
rect 21913 4981 21925 5015
rect 21959 5012 21971 5015
rect 22462 5012 22468 5024
rect 21959 4984 22468 5012
rect 21959 4981 21971 4984
rect 21913 4975 21971 4981
rect 22462 4972 22468 4984
rect 22520 4972 22526 5024
rect 22557 5015 22615 5021
rect 22557 4981 22569 5015
rect 22603 5012 22615 5015
rect 23198 5012 23204 5024
rect 22603 4984 23204 5012
rect 22603 4981 22615 4984
rect 22557 4975 22615 4981
rect 23198 4972 23204 4984
rect 23256 4972 23262 5024
rect 23293 5015 23351 5021
rect 23293 4981 23305 5015
rect 23339 5012 23351 5015
rect 24670 5012 24676 5024
rect 23339 4984 24676 5012
rect 23339 4981 23351 4984
rect 23293 4975 23351 4981
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 46845 5015 46903 5021
rect 46845 4981 46857 5015
rect 46891 5012 46903 5015
rect 47210 5012 47216 5024
rect 46891 4984 47216 5012
rect 46891 4981 46903 4984
rect 46845 4975 46903 4981
rect 47210 4972 47216 4984
rect 47268 4972 47274 5024
rect 48056 5021 48084 5052
rect 48041 5015 48099 5021
rect 48041 4981 48053 5015
rect 48087 4981 48099 5015
rect 48041 4975 48099 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 20806 4808 20812 4820
rect 20767 4780 20812 4808
rect 20806 4768 20812 4780
rect 20864 4768 20870 4820
rect 22738 4808 22744 4820
rect 22699 4780 22744 4808
rect 22738 4768 22744 4780
rect 22796 4768 22802 4820
rect 46382 4768 46388 4820
rect 46440 4808 46446 4820
rect 47578 4808 47584 4820
rect 46440 4780 47584 4808
rect 46440 4768 46446 4780
rect 47578 4768 47584 4780
rect 47636 4768 47642 4820
rect 24486 4632 24492 4684
rect 24544 4672 24550 4684
rect 25225 4675 25283 4681
rect 25225 4672 25237 4675
rect 24544 4644 25237 4672
rect 24544 4632 24550 4644
rect 25225 4641 25237 4644
rect 25271 4641 25283 4675
rect 25225 4635 25283 4641
rect 25409 4675 25467 4681
rect 25409 4641 25421 4675
rect 25455 4672 25467 4675
rect 44726 4672 44732 4684
rect 25455 4644 44732 4672
rect 25455 4641 25467 4644
rect 25409 4635 25467 4641
rect 44726 4632 44732 4644
rect 44784 4632 44790 4684
rect 45370 4632 45376 4684
rect 45428 4672 45434 4684
rect 47121 4675 47179 4681
rect 47121 4672 47133 4675
rect 45428 4644 47133 4672
rect 45428 4632 45434 4644
rect 47121 4641 47133 4644
rect 47167 4641 47179 4675
rect 47121 4635 47179 4641
rect 48133 4675 48191 4681
rect 48133 4641 48145 4675
rect 48179 4672 48191 4675
rect 48222 4672 48228 4684
rect 48179 4644 48228 4672
rect 48179 4641 48191 4644
rect 48133 4635 48191 4641
rect 48222 4632 48228 4644
rect 48280 4632 48286 4684
rect 10318 4564 10324 4616
rect 10376 4604 10382 4616
rect 10597 4607 10655 4613
rect 10597 4604 10609 4607
rect 10376 4576 10609 4604
rect 10376 4564 10382 4576
rect 10597 4573 10609 4576
rect 10643 4573 10655 4607
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 10597 4567 10655 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18966 4564 18972 4616
rect 19024 4604 19030 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19024 4576 19441 4604
rect 19024 4564 19030 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 20070 4604 20076 4616
rect 20031 4576 20076 4604
rect 19429 4567 19487 4573
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20714 4604 20720 4616
rect 20675 4576 20720 4604
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 21358 4604 21364 4616
rect 21319 4576 21364 4604
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 22002 4604 22008 4616
rect 21963 4576 22008 4604
rect 22002 4564 22008 4576
rect 22060 4564 22066 4616
rect 22462 4564 22468 4616
rect 22520 4604 22526 4616
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 22520 4576 22661 4604
rect 22520 4564 22526 4576
rect 22649 4573 22661 4576
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 23198 4564 23204 4616
rect 23256 4604 23262 4616
rect 23293 4607 23351 4613
rect 23293 4604 23305 4607
rect 23256 4576 23305 4604
rect 23256 4564 23262 4576
rect 23293 4573 23305 4576
rect 23339 4573 23351 4607
rect 23293 4567 23351 4573
rect 43806 4564 43812 4616
rect 43864 4604 43870 4616
rect 44085 4607 44143 4613
rect 44085 4604 44097 4607
rect 43864 4576 44097 4604
rect 43864 4564 43870 4576
rect 44085 4573 44097 4576
rect 44131 4573 44143 4607
rect 44085 4567 44143 4573
rect 45925 4607 45983 4613
rect 45925 4573 45937 4607
rect 45971 4573 45983 4607
rect 46382 4604 46388 4616
rect 46343 4576 46388 4604
rect 45925 4567 45983 4573
rect 19334 4496 19340 4548
rect 19392 4536 19398 4548
rect 20165 4539 20223 4545
rect 20165 4536 20177 4539
rect 19392 4508 20177 4536
rect 19392 4496 19398 4508
rect 20165 4505 20177 4508
rect 20211 4505 20223 4539
rect 27062 4536 27068 4548
rect 26975 4508 27068 4536
rect 20165 4499 20223 4505
rect 27062 4496 27068 4508
rect 27120 4536 27126 4548
rect 27246 4536 27252 4548
rect 27120 4508 27252 4536
rect 27120 4496 27126 4508
rect 27246 4496 27252 4508
rect 27304 4496 27310 4548
rect 39666 4496 39672 4548
rect 39724 4536 39730 4548
rect 45186 4536 45192 4548
rect 39724 4508 45192 4536
rect 39724 4496 39730 4508
rect 45186 4496 45192 4508
rect 45244 4496 45250 4548
rect 45940 4536 45968 4567
rect 46382 4564 46388 4576
rect 46440 4564 46446 4616
rect 45940 4508 46980 4536
rect 18601 4471 18659 4477
rect 18601 4437 18613 4471
rect 18647 4468 18659 4471
rect 18782 4468 18788 4480
rect 18647 4440 18788 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 19521 4471 19579 4477
rect 19521 4468 19533 4471
rect 19484 4440 19533 4468
rect 19484 4428 19490 4440
rect 19521 4437 19533 4440
rect 19567 4437 19579 4471
rect 19521 4431 19579 4437
rect 21453 4471 21511 4477
rect 21453 4437 21465 4471
rect 21499 4468 21511 4471
rect 21818 4468 21824 4480
rect 21499 4440 21824 4468
rect 21499 4437 21511 4440
rect 21453 4431 21511 4437
rect 21818 4428 21824 4440
rect 21876 4428 21882 4480
rect 22097 4471 22155 4477
rect 22097 4437 22109 4471
rect 22143 4468 22155 4471
rect 23198 4468 23204 4480
rect 22143 4440 23204 4468
rect 22143 4437 22155 4440
rect 22097 4431 22155 4437
rect 23198 4428 23204 4440
rect 23256 4428 23262 4480
rect 23385 4471 23443 4477
rect 23385 4437 23397 4471
rect 23431 4468 23443 4471
rect 23842 4468 23848 4480
rect 23431 4440 23848 4468
rect 23431 4437 23443 4440
rect 23385 4431 23443 4437
rect 23842 4428 23848 4440
rect 23900 4428 23906 4480
rect 43714 4428 43720 4480
rect 43772 4468 43778 4480
rect 43901 4471 43959 4477
rect 43901 4468 43913 4471
rect 43772 4440 43913 4468
rect 43772 4428 43778 4440
rect 43901 4437 43913 4440
rect 43947 4437 43959 4471
rect 45738 4468 45744 4480
rect 45699 4440 45744 4468
rect 43901 4431 43959 4437
rect 45738 4428 45744 4440
rect 45796 4428 45802 4480
rect 46474 4468 46480 4480
rect 46435 4440 46480 4468
rect 46474 4428 46480 4440
rect 46532 4428 46538 4480
rect 46952 4468 46980 4508
rect 47210 4496 47216 4548
rect 47268 4536 47274 4548
rect 47268 4508 47313 4536
rect 47268 4496 47274 4508
rect 47026 4468 47032 4480
rect 46952 4440 47032 4468
rect 47026 4428 47032 4440
rect 47084 4428 47090 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 18141 4267 18199 4273
rect 18141 4233 18153 4267
rect 18187 4264 18199 4267
rect 18506 4264 18512 4276
rect 18187 4236 18512 4264
rect 18187 4233 18199 4236
rect 18141 4227 18199 4233
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 19521 4267 19579 4273
rect 19521 4233 19533 4267
rect 19567 4264 19579 4267
rect 20070 4264 20076 4276
rect 19567 4236 20076 4264
rect 19567 4233 19579 4236
rect 19521 4227 19579 4233
rect 20070 4224 20076 4236
rect 20128 4224 20134 4276
rect 40586 4264 40592 4276
rect 24596 4236 24992 4264
rect 40547 4236 40592 4264
rect 17604 4168 18184 4196
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4128 10195 4131
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 10183 4100 10425 4128
rect 10183 4097 10195 4100
rect 10137 4091 10195 4097
rect 10413 4097 10425 4100
rect 10459 4128 10471 4131
rect 17405 4131 17463 4137
rect 10459 4100 17264 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 8772 4060 8800 4091
rect 15654 4060 15660 4072
rect 3476 4032 6914 4060
rect 8772 4032 15660 4060
rect 3476 4020 3482 4032
rect 6886 3992 6914 4032
rect 15654 4020 15660 4032
rect 15712 4020 15718 4072
rect 16666 3992 16672 4004
rect 6886 3964 16672 3992
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1728 3896 2145 3924
rect 1728 3884 1734 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2133 3887 2191 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2832 3896 2881 3924
rect 2832 3884 2838 3896
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 2869 3887 2927 3893
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8849 3927 8907 3933
rect 8849 3924 8861 3927
rect 8168 3896 8861 3924
rect 8168 3884 8174 3896
rect 8849 3893 8861 3896
rect 8895 3893 8907 3927
rect 8849 3887 8907 3893
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 9180 3896 9597 3924
rect 9180 3884 9186 3896
rect 9585 3893 9597 3896
rect 9631 3893 9643 3927
rect 10502 3924 10508 3936
rect 10463 3896 10508 3924
rect 9585 3887 9643 3893
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 17236 3924 17264 4100
rect 17405 4097 17417 4131
rect 17451 4128 17463 4131
rect 17604 4128 17632 4168
rect 17451 4100 17632 4128
rect 17451 4097 17463 4100
rect 17405 4091 17463 4097
rect 17678 4088 17684 4140
rect 17736 4128 17742 4140
rect 18049 4131 18107 4137
rect 18049 4128 18061 4131
rect 17736 4100 18061 4128
rect 17736 4088 17742 4100
rect 18049 4097 18061 4100
rect 18095 4097 18107 4131
rect 18156 4128 18184 4168
rect 18506 4128 18512 4140
rect 18156 4100 18512 4128
rect 18049 4091 18107 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18785 4131 18843 4137
rect 18785 4097 18797 4131
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4128 18935 4131
rect 18966 4128 18972 4140
rect 18923 4100 18972 4128
rect 18923 4097 18935 4100
rect 18877 4091 18935 4097
rect 17497 4063 17555 4069
rect 17497 4029 17509 4063
rect 17543 4060 17555 4063
rect 18800 4060 18828 4091
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19426 4128 19432 4140
rect 19387 4100 19432 4128
rect 19426 4088 19432 4100
rect 19484 4088 19490 4140
rect 20625 4131 20683 4137
rect 20625 4097 20637 4131
rect 20671 4128 20683 4131
rect 21634 4128 21640 4140
rect 20671 4100 21640 4128
rect 20671 4097 20683 4100
rect 20625 4091 20683 4097
rect 21634 4088 21640 4100
rect 21692 4088 21698 4140
rect 21818 4128 21824 4140
rect 21779 4100 21824 4128
rect 21818 4088 21824 4100
rect 21876 4088 21882 4140
rect 21913 4131 21971 4137
rect 21913 4097 21925 4131
rect 21959 4128 21971 4131
rect 22465 4131 22523 4137
rect 22465 4128 22477 4131
rect 21959 4100 22477 4128
rect 21959 4097 21971 4100
rect 21913 4091 21971 4097
rect 22465 4097 22477 4100
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 23201 4131 23259 4137
rect 23201 4097 23213 4131
rect 23247 4097 23259 4131
rect 23842 4128 23848 4140
rect 23803 4100 23848 4128
rect 23201 4091 23259 4097
rect 17543 4032 18828 4060
rect 23216 4060 23244 4091
rect 23842 4088 23848 4100
rect 23900 4088 23906 4140
rect 24596 4060 24624 4236
rect 24673 4131 24731 4137
rect 24673 4097 24685 4131
rect 24719 4097 24731 4131
rect 24964 4128 24992 4236
rect 40586 4224 40592 4236
rect 40644 4224 40650 4276
rect 45278 4264 45284 4276
rect 40972 4236 45284 4264
rect 40972 4196 41000 4236
rect 38626 4168 41000 4196
rect 28442 4128 28448 4140
rect 24964 4100 28448 4128
rect 24673 4091 24731 4097
rect 23216 4032 24624 4060
rect 17543 4029 17555 4032
rect 17497 4023 17555 4029
rect 22186 3992 22192 4004
rect 17512 3964 22192 3992
rect 17512 3924 17540 3964
rect 22186 3952 22192 3964
rect 22244 3952 22250 4004
rect 22830 3952 22836 4004
rect 22888 3992 22894 4004
rect 24688 3992 24716 4091
rect 28442 4088 28448 4100
rect 28500 4088 28506 4140
rect 35894 4128 35900 4140
rect 28966 4100 35900 4128
rect 24946 4020 24952 4072
rect 25004 4060 25010 4072
rect 28966 4060 28994 4100
rect 35894 4088 35900 4100
rect 35952 4128 35958 4140
rect 38470 4128 38476 4140
rect 35952 4100 38476 4128
rect 35952 4088 35958 4100
rect 38470 4088 38476 4100
rect 38528 4128 38534 4140
rect 38626 4128 38654 4168
rect 39850 4128 39856 4140
rect 38528 4100 38654 4128
rect 39811 4100 39856 4128
rect 38528 4088 38534 4100
rect 39850 4088 39856 4100
rect 39908 4088 39914 4140
rect 40494 4128 40500 4140
rect 40455 4100 40500 4128
rect 40494 4088 40500 4100
rect 40552 4088 40558 4140
rect 40972 4128 41000 4168
rect 41046 4156 41052 4208
rect 41104 4196 41110 4208
rect 41104 4168 42932 4196
rect 41104 4156 41110 4168
rect 42904 4137 42932 4168
rect 43548 4137 43576 4236
rect 45278 4224 45284 4236
rect 45336 4224 45342 4276
rect 43714 4196 43720 4208
rect 43675 4168 43720 4196
rect 43714 4156 43720 4168
rect 43772 4156 43778 4208
rect 46382 4156 46388 4208
rect 46440 4196 46446 4208
rect 46569 4199 46627 4205
rect 46569 4196 46581 4199
rect 46440 4168 46581 4196
rect 46440 4156 46446 4168
rect 46569 4165 46581 4168
rect 46615 4165 46627 4199
rect 47762 4196 47768 4208
rect 47723 4168 47768 4196
rect 46569 4159 46627 4165
rect 47762 4156 47768 4168
rect 47820 4156 47826 4208
rect 41141 4131 41199 4137
rect 41141 4128 41153 4131
rect 40972 4100 41153 4128
rect 41141 4097 41153 4100
rect 41187 4097 41199 4131
rect 41141 4091 41199 4097
rect 42889 4131 42947 4137
rect 42889 4097 42901 4131
rect 42935 4097 42947 4131
rect 42889 4091 42947 4097
rect 43533 4131 43591 4137
rect 43533 4097 43545 4131
rect 43579 4097 43591 4131
rect 43533 4091 43591 4097
rect 25004 4032 28994 4060
rect 25004 4020 25010 4032
rect 33778 4020 33784 4072
rect 33836 4060 33842 4072
rect 41325 4063 41383 4069
rect 33836 4032 40724 4060
rect 33836 4020 33842 4032
rect 22888 3964 24716 3992
rect 22888 3952 22894 3964
rect 24854 3952 24860 4004
rect 24912 3992 24918 4004
rect 40696 3992 40724 4032
rect 41325 4029 41337 4063
rect 41371 4060 41383 4063
rect 41690 4060 41696 4072
rect 41371 4032 41696 4060
rect 41371 4029 41383 4032
rect 41325 4023 41383 4029
rect 41690 4020 41696 4032
rect 41748 4020 41754 4072
rect 42904 4060 42932 4091
rect 44910 4088 44916 4140
rect 44968 4128 44974 4140
rect 44968 4100 45140 4128
rect 44968 4088 44974 4100
rect 45002 4060 45008 4072
rect 42904 4032 45008 4060
rect 45002 4020 45008 4032
rect 45060 4020 45066 4072
rect 45112 4069 45140 4100
rect 45097 4063 45155 4069
rect 45097 4029 45109 4063
rect 45143 4029 45155 4063
rect 45097 4023 45155 4029
rect 41046 3992 41052 4004
rect 24912 3964 26234 3992
rect 24912 3952 24918 3964
rect 17236 3896 17540 3924
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 20717 3927 20775 3933
rect 20717 3924 20729 3927
rect 20220 3896 20729 3924
rect 20220 3884 20226 3896
rect 20717 3893 20729 3896
rect 20763 3893 20775 3927
rect 20717 3887 20775 3893
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 22557 3927 22615 3933
rect 22557 3924 22569 3927
rect 21416 3896 22569 3924
rect 21416 3884 21422 3896
rect 22557 3893 22569 3896
rect 22603 3893 22615 3927
rect 22557 3887 22615 3893
rect 22738 3884 22744 3936
rect 22796 3924 22802 3936
rect 23293 3927 23351 3933
rect 23293 3924 23305 3927
rect 22796 3896 23305 3924
rect 22796 3884 22802 3896
rect 23293 3893 23305 3896
rect 23339 3893 23351 3927
rect 23934 3924 23940 3936
rect 23895 3896 23940 3924
rect 23293 3887 23351 3893
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 24762 3924 24768 3936
rect 24723 3896 24768 3924
rect 24762 3884 24768 3896
rect 24820 3884 24826 3936
rect 25498 3924 25504 3936
rect 25459 3896 25504 3924
rect 25498 3884 25504 3896
rect 25556 3884 25562 3936
rect 26206 3924 26234 3964
rect 38626 3964 40632 3992
rect 40696 3964 41052 3992
rect 38626 3924 38654 3964
rect 26206 3896 38654 3924
rect 39574 3884 39580 3936
rect 39632 3924 39638 3936
rect 39945 3927 40003 3933
rect 39945 3924 39957 3927
rect 39632 3896 39957 3924
rect 39632 3884 39638 3896
rect 39945 3893 39957 3896
rect 39991 3893 40003 3927
rect 40604 3924 40632 3964
rect 41046 3952 41052 3964
rect 41104 3952 41110 4004
rect 47949 3995 48007 4001
rect 47949 3992 47961 3995
rect 41432 3964 47961 3992
rect 41432 3924 41460 3964
rect 47949 3961 47961 3964
rect 47995 3961 48007 3995
rect 47949 3955 48007 3961
rect 40604 3896 41460 3924
rect 39945 3887 40003 3893
rect 41506 3884 41512 3936
rect 41564 3924 41570 3936
rect 41564 3896 41609 3924
rect 41564 3884 41570 3896
rect 42886 3884 42892 3936
rect 42944 3924 42950 3936
rect 42981 3927 43039 3933
rect 42981 3924 42993 3927
rect 42944 3896 42993 3924
rect 42944 3884 42950 3896
rect 42981 3893 42993 3896
rect 43027 3893 43039 3927
rect 42981 3887 43039 3893
rect 46017 3927 46075 3933
rect 46017 3893 46029 3927
rect 46063 3924 46075 3927
rect 46290 3924 46296 3936
rect 46063 3896 46296 3924
rect 46063 3893 46075 3896
rect 46017 3887 46075 3893
rect 46290 3884 46296 3896
rect 46348 3884 46354 3936
rect 46658 3924 46664 3936
rect 46619 3896 46664 3924
rect 46658 3884 46664 3896
rect 46716 3884 46722 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 17678 3720 17684 3732
rect 9723 3692 17264 3720
rect 17639 3692 17684 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 6638 3612 6644 3664
rect 6696 3652 6702 3664
rect 17236 3652 17264 3692
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 19429 3723 19487 3729
rect 19429 3689 19441 3723
rect 19475 3720 19487 3723
rect 20714 3720 20720 3732
rect 19475 3692 20720 3720
rect 19475 3689 19487 3692
rect 19429 3683 19487 3689
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 23014 3720 23020 3732
rect 22066 3692 23020 3720
rect 6696 3624 14136 3652
rect 17236 3624 18552 3652
rect 6696 3612 6702 3624
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1360 3488 1409 3516
rect 1360 3476 1366 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 2130 3516 2136 3528
rect 2091 3488 2136 3516
rect 1397 3479 1455 3485
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3516 6699 3519
rect 6886 3516 6914 3624
rect 7006 3544 7012 3596
rect 7064 3584 7070 3596
rect 10318 3584 10324 3596
rect 7064 3556 10180 3584
rect 10279 3556 10324 3584
rect 7064 3544 7070 3556
rect 7466 3516 7472 3528
rect 6687 3488 6914 3516
rect 7427 3488 7472 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 1762 3408 1768 3460
rect 1820 3448 1826 3460
rect 2976 3448 3004 3479
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7984 3488 8217 3516
rect 7984 3476 7990 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 1820 3420 3004 3448
rect 1820 3408 1826 3420
rect 8386 3408 8392 3460
rect 8444 3448 8450 3460
rect 9401 3451 9459 3457
rect 9401 3448 9413 3451
rect 8444 3420 9413 3448
rect 8444 3408 8450 3420
rect 9401 3417 9413 3420
rect 9447 3417 9459 3451
rect 10152 3448 10180 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 10502 3584 10508 3596
rect 10463 3556 10508 3584
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 13538 3516 13544 3528
rect 13499 3488 13544 3516
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 14108 3525 14136 3624
rect 17494 3544 17500 3596
rect 17552 3584 17558 3596
rect 17552 3556 18460 3584
rect 17552 3544 17558 3556
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 15289 3519 15347 3525
rect 15289 3485 15301 3519
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 17589 3519 17647 3525
rect 17589 3485 17601 3519
rect 17635 3516 17647 3519
rect 17954 3516 17960 3528
rect 17635 3488 17960 3516
rect 17635 3485 17647 3488
rect 17589 3479 17647 3485
rect 15304 3448 15332 3479
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18230 3516 18236 3528
rect 18191 3488 18236 3516
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 15470 3448 15476 3460
rect 10152 3420 15332 3448
rect 15431 3420 15476 3448
rect 9401 3411 9459 3417
rect 15470 3408 15476 3420
rect 15528 3408 15534 3460
rect 17126 3448 17132 3460
rect 17087 3420 17132 3448
rect 17126 3408 17132 3420
rect 17184 3408 17190 3460
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 1946 3340 1952 3392
rect 2004 3380 2010 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 2004 3352 2237 3380
rect 2004 3340 2010 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 6730 3380 6736 3392
rect 6691 3352 6736 3380
rect 2225 3343 2283 3349
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 13780 3352 14197 3380
rect 13780 3340 13786 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 18322 3380 18328 3392
rect 18283 3352 18328 3380
rect 14185 3343 14243 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 18432 3380 18460 3556
rect 18524 3448 18552 3624
rect 20070 3612 20076 3664
rect 20128 3652 20134 3664
rect 20128 3624 20484 3652
rect 20128 3612 20134 3624
rect 20162 3584 20168 3596
rect 20123 3556 20168 3584
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 20456 3593 20484 3624
rect 20530 3612 20536 3664
rect 20588 3652 20594 3664
rect 22066 3652 22094 3692
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 23106 3680 23112 3732
rect 23164 3720 23170 3732
rect 24857 3723 24915 3729
rect 24857 3720 24869 3723
rect 23164 3692 24869 3720
rect 23164 3680 23170 3692
rect 24857 3689 24869 3692
rect 24903 3689 24915 3723
rect 24857 3683 24915 3689
rect 25866 3680 25872 3732
rect 25924 3720 25930 3732
rect 39114 3720 39120 3732
rect 25924 3692 39120 3720
rect 25924 3680 25930 3692
rect 39114 3680 39120 3692
rect 39172 3680 39178 3732
rect 39209 3723 39267 3729
rect 39209 3689 39221 3723
rect 39255 3720 39267 3723
rect 40494 3720 40500 3732
rect 39255 3692 40500 3720
rect 39255 3689 39267 3692
rect 39209 3683 39267 3689
rect 40494 3680 40500 3692
rect 40552 3680 40558 3732
rect 45830 3720 45836 3732
rect 41248 3692 45836 3720
rect 20588 3624 22094 3652
rect 20588 3612 20594 3624
rect 22370 3612 22376 3664
rect 22428 3652 22434 3664
rect 23293 3655 23351 3661
rect 23293 3652 23305 3655
rect 22428 3624 23305 3652
rect 22428 3612 22434 3624
rect 23293 3621 23305 3624
rect 23339 3621 23351 3655
rect 23293 3615 23351 3621
rect 23382 3612 23388 3664
rect 23440 3652 23446 3664
rect 23440 3624 26234 3652
rect 23440 3612 23446 3624
rect 20441 3587 20499 3593
rect 20441 3553 20453 3587
rect 20487 3553 20499 3587
rect 20441 3547 20499 3553
rect 20990 3544 20996 3596
rect 21048 3584 21054 3596
rect 23934 3584 23940 3596
rect 21048 3556 23940 3584
rect 21048 3544 21054 3556
rect 23934 3544 23940 3556
rect 23992 3544 23998 3596
rect 25406 3584 25412 3596
rect 25367 3556 25412 3584
rect 25406 3544 25412 3556
rect 25464 3544 25470 3596
rect 26206 3584 26234 3624
rect 28902 3612 28908 3664
rect 28960 3652 28966 3664
rect 41248 3652 41276 3692
rect 45830 3680 45836 3692
rect 45888 3680 45894 3732
rect 47486 3652 47492 3664
rect 28960 3624 30972 3652
rect 28960 3612 28966 3624
rect 29546 3584 29552 3596
rect 26206 3556 29408 3584
rect 29507 3556 29552 3584
rect 19334 3516 19340 3528
rect 19295 3488 19340 3516
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19978 3516 19984 3528
rect 19939 3488 19984 3516
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 22554 3476 22560 3528
rect 22612 3516 22618 3528
rect 22741 3519 22799 3525
rect 22741 3516 22753 3519
rect 22612 3488 22753 3516
rect 22612 3476 22618 3488
rect 22741 3485 22753 3488
rect 22787 3485 22799 3519
rect 23198 3516 23204 3528
rect 23159 3488 23204 3516
rect 22741 3479 22799 3485
rect 23198 3476 23204 3488
rect 23256 3476 23262 3528
rect 24854 3516 24860 3528
rect 23308 3488 24860 3516
rect 18524 3420 22094 3448
rect 20806 3380 20812 3392
rect 18432 3352 20812 3380
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 22066 3380 22094 3420
rect 22646 3408 22652 3460
rect 22704 3448 22710 3460
rect 23308 3448 23336 3488
rect 24854 3476 24860 3488
rect 24912 3476 24918 3528
rect 22704 3420 23336 3448
rect 22704 3408 22710 3420
rect 24486 3408 24492 3460
rect 24544 3448 24550 3460
rect 24765 3451 24823 3457
rect 24765 3448 24777 3451
rect 24544 3420 24777 3448
rect 24544 3408 24550 3420
rect 24765 3417 24777 3420
rect 24811 3417 24823 3451
rect 25590 3448 25596 3460
rect 25551 3420 25596 3448
rect 24765 3411 24823 3417
rect 25590 3408 25596 3420
rect 25648 3408 25654 3460
rect 27246 3448 27252 3460
rect 27207 3420 27252 3448
rect 27246 3408 27252 3420
rect 27304 3408 27310 3460
rect 24578 3380 24584 3392
rect 22066 3352 24584 3380
rect 24578 3340 24584 3352
rect 24636 3340 24642 3392
rect 29380 3380 29408 3556
rect 29546 3544 29552 3556
rect 29604 3544 29610 3596
rect 30944 3516 30972 3624
rect 31404 3624 41276 3652
rect 41386 3624 44128 3652
rect 31404 3593 31432 3624
rect 31389 3587 31447 3593
rect 31389 3553 31401 3587
rect 31435 3553 31447 3587
rect 39942 3584 39948 3596
rect 31389 3547 31447 3553
rect 31496 3556 39948 3584
rect 31496 3516 31524 3556
rect 39942 3544 39948 3556
rect 40000 3544 40006 3596
rect 40034 3544 40040 3596
rect 40092 3584 40098 3596
rect 40092 3556 40137 3584
rect 40092 3544 40098 3556
rect 40678 3544 40684 3596
rect 40736 3584 40742 3596
rect 41386 3584 41414 3624
rect 40736 3556 41414 3584
rect 40736 3544 40742 3556
rect 41506 3544 41512 3596
rect 41564 3584 41570 3596
rect 41564 3556 41609 3584
rect 41564 3544 41570 3556
rect 30944 3488 31524 3516
rect 33045 3519 33103 3525
rect 33045 3485 33057 3519
rect 33091 3516 33103 3519
rect 33778 3516 33784 3528
rect 33091 3488 33784 3516
rect 33091 3485 33103 3488
rect 33045 3479 33103 3485
rect 33778 3476 33784 3488
rect 33836 3476 33842 3528
rect 33873 3519 33931 3525
rect 33873 3485 33885 3519
rect 33919 3485 33931 3519
rect 35894 3516 35900 3528
rect 35855 3488 35900 3516
rect 33873 3479 33931 3485
rect 29730 3448 29736 3460
rect 29691 3420 29736 3448
rect 29730 3408 29736 3420
rect 29788 3408 29794 3460
rect 32950 3408 32956 3460
rect 33008 3448 33014 3460
rect 33888 3448 33916 3479
rect 35894 3476 35900 3488
rect 35952 3476 35958 3528
rect 37734 3516 37740 3528
rect 37695 3488 37740 3516
rect 37734 3476 37740 3488
rect 37792 3476 37798 3528
rect 39117 3519 39175 3525
rect 39117 3485 39129 3519
rect 39163 3516 39175 3519
rect 39206 3516 39212 3528
rect 39163 3488 39212 3516
rect 39163 3485 39175 3488
rect 39117 3479 39175 3485
rect 39206 3476 39212 3488
rect 39264 3476 39270 3528
rect 40313 3519 40371 3525
rect 40313 3485 40325 3519
rect 40359 3485 40371 3519
rect 43993 3519 44051 3525
rect 43993 3516 44005 3519
rect 40313 3479 40371 3485
rect 42904 3488 44005 3516
rect 33008 3420 33916 3448
rect 36081 3451 36139 3457
rect 33008 3408 33014 3420
rect 36081 3417 36093 3451
rect 36127 3448 36139 3451
rect 36170 3448 36176 3460
rect 36127 3420 36176 3448
rect 36127 3417 36139 3420
rect 36081 3411 36139 3417
rect 36170 3408 36176 3420
rect 36228 3408 36234 3460
rect 37752 3448 37780 3476
rect 39666 3448 39672 3460
rect 37752 3420 39672 3448
rect 39666 3408 39672 3420
rect 39724 3408 39730 3460
rect 39758 3408 39764 3460
rect 39816 3448 39822 3460
rect 40328 3448 40356 3479
rect 41690 3448 41696 3460
rect 39816 3420 40356 3448
rect 41651 3420 41696 3448
rect 39816 3408 39822 3420
rect 41690 3408 41696 3420
rect 41748 3408 41754 3460
rect 42702 3408 42708 3460
rect 42760 3448 42766 3460
rect 42904 3448 42932 3488
rect 43993 3485 44005 3488
rect 44039 3485 44051 3519
rect 43993 3479 44051 3485
rect 42760 3420 42932 3448
rect 43349 3451 43407 3457
rect 42760 3408 42766 3420
rect 43349 3417 43361 3451
rect 43395 3448 43407 3451
rect 44100 3448 44128 3624
rect 45664 3624 47492 3652
rect 45186 3516 45192 3528
rect 45147 3488 45192 3516
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 45664 3525 45692 3624
rect 47486 3612 47492 3624
rect 47544 3612 47550 3664
rect 46290 3584 46296 3596
rect 46251 3556 46296 3584
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 46474 3584 46480 3596
rect 46435 3556 46480 3584
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 45649 3519 45707 3525
rect 45649 3485 45661 3519
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 47670 3448 47676 3460
rect 43395 3420 47676 3448
rect 43395 3417 43407 3420
rect 43349 3411 43407 3417
rect 47670 3408 47676 3420
rect 47728 3408 47734 3460
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 32214 3380 32220 3392
rect 29380 3352 32220 3380
rect 32214 3340 32220 3352
rect 32272 3340 32278 3392
rect 33134 3380 33140 3392
rect 33095 3352 33140 3380
rect 33134 3340 33140 3352
rect 33192 3340 33198 3392
rect 33870 3340 33876 3392
rect 33928 3380 33934 3392
rect 42518 3380 42524 3392
rect 33928 3352 42524 3380
rect 33928 3340 33934 3352
rect 42518 3340 42524 3352
rect 42576 3340 42582 3392
rect 45370 3340 45376 3392
rect 45428 3380 45434 3392
rect 45741 3383 45799 3389
rect 45741 3380 45753 3383
rect 45428 3352 45753 3380
rect 45428 3340 45434 3352
rect 45741 3349 45753 3352
rect 45787 3349 45799 3383
rect 45741 3343 45799 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 18230 3176 18236 3188
rect 1636 3148 14688 3176
rect 18191 3148 18236 3176
rect 1636 3136 1642 3148
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 8110 3108 8116 3120
rect 8071 3080 8116 3108
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 13722 3108 13728 3120
rect 13683 3080 13728 3108
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 14660 3108 14688 3148
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 18874 3176 18880 3188
rect 18835 3148 18880 3176
rect 18874 3136 18880 3148
rect 18932 3136 18938 3188
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 20530 3176 20536 3188
rect 19392 3148 20536 3176
rect 19392 3136 19398 3148
rect 20530 3136 20536 3148
rect 20588 3136 20594 3188
rect 20809 3179 20867 3185
rect 20809 3145 20821 3179
rect 20855 3176 20867 3179
rect 22002 3176 22008 3188
rect 20855 3148 22008 3176
rect 20855 3145 20867 3148
rect 20809 3139 20867 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 35802 3176 35808 3188
rect 22244 3148 23980 3176
rect 22244 3136 22250 3148
rect 22094 3108 22100 3120
rect 14660 3080 22100 3108
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 22738 3108 22744 3120
rect 22699 3080 22744 3108
rect 22738 3068 22744 3080
rect 22796 3068 22802 3120
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 7926 3040 7932 3052
rect 7887 3012 7932 3040
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3009 10287 3043
rect 13538 3040 13544 3052
rect 13499 3012 13544 3040
rect 10229 3003 10287 3009
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 716 2944 2237 2972
rect 716 2932 722 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 7800 2944 8401 2972
rect 7800 2932 7806 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 10244 2904 10272 3003
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 17313 3043 17371 3049
rect 17313 3009 17325 3043
rect 17359 3009 17371 3043
rect 18141 3043 18199 3049
rect 18141 3040 18153 3043
rect 17313 3003 17371 3009
rect 17696 3012 18153 3040
rect 14182 2972 14188 2984
rect 14143 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 15194 2932 15200 2984
rect 15252 2972 15258 2984
rect 17221 2975 17279 2981
rect 17221 2972 17233 2975
rect 15252 2944 17233 2972
rect 15252 2932 15258 2944
rect 17221 2941 17233 2944
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 17328 2904 17356 3003
rect 17696 2981 17724 3012
rect 18141 3009 18153 3012
rect 18187 3009 18199 3043
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 18141 3003 18199 3009
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3009 19487 3043
rect 19429 3003 19487 3009
rect 17681 2975 17739 2981
rect 17681 2941 17693 2975
rect 17727 2941 17739 2975
rect 19444 2972 19472 3003
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 20036 3012 20269 3040
rect 20036 3000 20042 3012
rect 20257 3009 20269 3012
rect 20303 3009 20315 3043
rect 20257 3003 20315 3009
rect 20717 3043 20775 3049
rect 20717 3009 20729 3043
rect 20763 3040 20775 3043
rect 21358 3040 21364 3052
rect 20763 3012 21364 3040
rect 20763 3009 20775 3012
rect 20717 3003 20775 3009
rect 21358 3000 21364 3012
rect 21416 3000 21422 3052
rect 21910 3040 21916 3052
rect 21871 3012 21916 3040
rect 21910 3000 21916 3012
rect 21968 3000 21974 3052
rect 22554 3040 22560 3052
rect 22515 3012 22560 3040
rect 22554 3000 22560 3012
rect 22612 3000 22618 3052
rect 20622 2972 20628 2984
rect 19444 2944 20628 2972
rect 17681 2935 17739 2941
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 20864 2944 22232 2972
rect 20864 2932 20870 2944
rect 22094 2904 22100 2916
rect 10244 2876 12434 2904
rect 17328 2876 20852 2904
rect 22055 2876 22100 2904
rect 10318 2836 10324 2848
rect 10279 2808 10324 2836
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 12406 2836 12434 2876
rect 18690 2836 18696 2848
rect 12406 2808 18696 2836
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 19521 2839 19579 2845
rect 19521 2805 19533 2839
rect 19567 2836 19579 2839
rect 20714 2836 20720 2848
rect 19567 2808 20720 2836
rect 19567 2805 19579 2808
rect 19521 2799 19579 2805
rect 20714 2796 20720 2808
rect 20772 2796 20778 2848
rect 20824 2836 20852 2876
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 22204 2904 22232 2944
rect 22462 2932 22468 2984
rect 22520 2972 22526 2984
rect 23017 2975 23075 2981
rect 23017 2972 23029 2975
rect 22520 2944 23029 2972
rect 22520 2932 22526 2944
rect 23017 2941 23029 2944
rect 23063 2941 23075 2975
rect 23017 2935 23075 2941
rect 23106 2932 23112 2984
rect 23164 2972 23170 2984
rect 23952 2972 23980 3148
rect 25056 3148 35808 3176
rect 24670 3068 24676 3120
rect 24728 3108 24734 3120
rect 25056 3117 25084 3148
rect 35802 3136 35808 3148
rect 35860 3136 35866 3188
rect 36170 3176 36176 3188
rect 36131 3148 36176 3176
rect 36170 3136 36176 3148
rect 36228 3136 36234 3188
rect 39117 3179 39175 3185
rect 39117 3145 39129 3179
rect 39163 3176 39175 3179
rect 39850 3176 39856 3188
rect 39163 3148 39856 3176
rect 39163 3145 39175 3148
rect 39117 3139 39175 3145
rect 39850 3136 39856 3148
rect 39908 3136 39914 3188
rect 40126 3136 40132 3188
rect 40184 3176 40190 3188
rect 47857 3179 47915 3185
rect 47857 3176 47869 3179
rect 40184 3148 47869 3176
rect 40184 3136 40190 3148
rect 47857 3145 47869 3148
rect 47903 3145 47915 3179
rect 47857 3139 47915 3145
rect 24949 3111 25007 3117
rect 24949 3108 24961 3111
rect 24728 3080 24961 3108
rect 24728 3068 24734 3080
rect 24949 3077 24961 3080
rect 24995 3077 25007 3111
rect 24949 3071 25007 3077
rect 25041 3111 25099 3117
rect 25041 3077 25053 3111
rect 25087 3077 25099 3111
rect 25958 3108 25964 3120
rect 25919 3080 25964 3108
rect 25041 3071 25099 3077
rect 25958 3068 25964 3080
rect 26016 3068 26022 3120
rect 27614 3108 27620 3120
rect 27575 3080 27620 3108
rect 27614 3068 27620 3080
rect 27672 3068 27678 3120
rect 33134 3108 33140 3120
rect 33095 3080 33140 3108
rect 33134 3068 33140 3080
rect 33192 3068 33198 3120
rect 40586 3108 40592 3120
rect 39592 3080 40592 3108
rect 27062 3000 27068 3052
rect 27120 3040 27126 3052
rect 27433 3043 27491 3049
rect 27433 3040 27445 3043
rect 27120 3012 27445 3040
rect 27120 3000 27126 3012
rect 27433 3009 27445 3012
rect 27479 3009 27491 3043
rect 32950 3040 32956 3052
rect 32911 3012 32956 3040
rect 27433 3003 27491 3009
rect 32950 3000 32956 3012
rect 33008 3000 33014 3052
rect 36078 3000 36084 3052
rect 36136 3040 36142 3052
rect 36357 3043 36415 3049
rect 36357 3040 36369 3043
rect 36136 3012 36369 3040
rect 36136 3000 36142 3012
rect 36357 3009 36369 3012
rect 36403 3009 36415 3043
rect 38470 3040 38476 3052
rect 38431 3012 38476 3040
rect 36357 3003 36415 3009
rect 38470 3000 38476 3012
rect 38528 3000 38534 3052
rect 39592 3049 39620 3080
rect 40586 3068 40592 3080
rect 40644 3068 40650 3120
rect 42886 3108 42892 3120
rect 42847 3080 42892 3108
rect 42886 3068 42892 3080
rect 42944 3068 42950 3120
rect 43162 3068 43168 3120
rect 43220 3108 43226 3120
rect 44545 3111 44603 3117
rect 44545 3108 44557 3111
rect 43220 3080 44557 3108
rect 43220 3068 43226 3080
rect 44545 3077 44557 3080
rect 44591 3077 44603 3111
rect 45370 3108 45376 3120
rect 45331 3080 45376 3108
rect 44545 3071 44603 3077
rect 45370 3068 45376 3080
rect 45428 3068 45434 3120
rect 39577 3043 39635 3049
rect 39577 3009 39589 3043
rect 39623 3009 39635 3043
rect 42702 3040 42708 3052
rect 39577 3003 39635 3009
rect 41386 3012 41644 3040
rect 42663 3012 42708 3040
rect 33502 2972 33508 2984
rect 23164 2944 23520 2972
rect 23952 2944 26234 2972
rect 33463 2944 33508 2972
rect 23164 2932 23170 2944
rect 23382 2904 23388 2916
rect 22204 2876 23388 2904
rect 23382 2864 23388 2876
rect 23440 2864 23446 2916
rect 23492 2904 23520 2944
rect 26050 2904 26056 2916
rect 23492 2876 26056 2904
rect 26050 2864 26056 2876
rect 26108 2864 26114 2916
rect 26206 2904 26234 2944
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 38657 2975 38715 2981
rect 38657 2941 38669 2975
rect 38703 2972 38715 2975
rect 39758 2972 39764 2984
rect 38703 2944 39764 2972
rect 38703 2941 38715 2944
rect 38657 2935 38715 2941
rect 39758 2932 39764 2944
rect 39816 2932 39822 2984
rect 39850 2932 39856 2984
rect 39908 2972 39914 2984
rect 40037 2975 40095 2981
rect 40037 2972 40049 2975
rect 39908 2944 40049 2972
rect 39908 2932 39914 2944
rect 40037 2941 40049 2944
rect 40083 2972 40095 2975
rect 40678 2972 40684 2984
rect 40083 2944 40684 2972
rect 40083 2941 40095 2944
rect 40037 2935 40095 2941
rect 40678 2932 40684 2944
rect 40736 2932 40742 2984
rect 41386 2904 41414 3012
rect 41616 2972 41644 3012
rect 42702 3000 42708 3012
rect 42760 3000 42766 3052
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 47762 3040 47768 3052
rect 47723 3012 47768 3040
rect 47762 3000 47768 3012
rect 47820 3000 47826 3052
rect 46934 2972 46940 2984
rect 41616 2944 46940 2972
rect 46934 2932 46940 2944
rect 46992 2932 46998 2984
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 26206 2876 39804 2904
rect 27246 2836 27252 2848
rect 20824 2808 27252 2836
rect 27246 2796 27252 2808
rect 27304 2836 27310 2848
rect 39666 2836 39672 2848
rect 27304 2808 39672 2836
rect 27304 2796 27310 2808
rect 39666 2796 39672 2808
rect 39724 2796 39730 2848
rect 39776 2836 39804 2876
rect 40052 2876 41414 2904
rect 40052 2836 40080 2876
rect 39776 2808 40080 2836
rect 40126 2796 40132 2848
rect 40184 2836 40190 2848
rect 45002 2836 45008 2848
rect 40184 2808 45008 2836
rect 40184 2796 40190 2808
rect 45002 2796 45008 2808
rect 45060 2796 45066 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 15470 2592 15476 2644
rect 15528 2632 15534 2644
rect 15565 2635 15623 2641
rect 15565 2632 15577 2635
rect 15528 2604 15577 2632
rect 15528 2592 15534 2604
rect 15565 2601 15577 2604
rect 15611 2601 15623 2635
rect 17954 2632 17960 2644
rect 17915 2604 17960 2632
rect 15565 2595 15623 2601
rect 17954 2592 17960 2604
rect 18012 2592 18018 2644
rect 18506 2592 18512 2644
rect 18564 2632 18570 2644
rect 18601 2635 18659 2641
rect 18601 2632 18613 2635
rect 18564 2604 18613 2632
rect 18564 2592 18570 2604
rect 18601 2601 18613 2604
rect 18647 2601 18659 2635
rect 20898 2632 20904 2644
rect 20859 2604 20904 2632
rect 18601 2595 18659 2601
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 21174 2592 21180 2644
rect 21232 2632 21238 2644
rect 22005 2635 22063 2641
rect 22005 2632 22017 2635
rect 21232 2604 22017 2632
rect 21232 2592 21238 2604
rect 22005 2601 22017 2604
rect 22051 2632 22063 2635
rect 24946 2632 24952 2644
rect 22051 2604 24952 2632
rect 22051 2601 22063 2604
rect 22005 2595 22063 2601
rect 24946 2592 24952 2604
rect 25004 2592 25010 2644
rect 26786 2592 26792 2644
rect 26844 2632 26850 2644
rect 28629 2635 28687 2641
rect 28629 2632 28641 2635
rect 26844 2604 28641 2632
rect 26844 2592 26850 2604
rect 28629 2601 28641 2604
rect 28675 2601 28687 2635
rect 29730 2632 29736 2644
rect 29691 2604 29736 2632
rect 28629 2595 28687 2601
rect 29730 2592 29736 2604
rect 29788 2592 29794 2644
rect 39206 2632 39212 2644
rect 39167 2604 39212 2632
rect 39206 2592 39212 2604
rect 39264 2592 39270 2644
rect 40402 2632 40408 2644
rect 40363 2604 40408 2632
rect 40402 2592 40408 2604
rect 40460 2592 40466 2644
rect 2774 2564 2780 2576
rect 1412 2536 2780 2564
rect 1412 2505 1440 2536
rect 2774 2524 2780 2536
rect 2832 2524 2838 2576
rect 15194 2564 15200 2576
rect 5276 2536 15200 2564
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2496 1639 2499
rect 1670 2496 1676 2508
rect 1627 2468 1676 2496
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 2866 2496 2872 2508
rect 2827 2468 2872 2496
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 5276 2505 5304 2536
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 17313 2567 17371 2573
rect 17313 2533 17325 2567
rect 17359 2564 17371 2567
rect 17586 2564 17592 2576
rect 17359 2536 17592 2564
rect 17359 2533 17371 2536
rect 17313 2527 17371 2533
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 20165 2567 20223 2573
rect 20165 2533 20177 2567
rect 20211 2564 20223 2567
rect 21082 2564 21088 2576
rect 20211 2536 21088 2564
rect 20211 2533 20223 2536
rect 20165 2527 20223 2533
rect 21082 2524 21088 2536
rect 21140 2524 21146 2576
rect 25498 2564 25504 2576
rect 24596 2536 25504 2564
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2465 5319 2499
rect 6730 2496 6736 2508
rect 6691 2468 6736 2496
rect 5261 2459 5319 2465
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 7098 2496 7104 2508
rect 7059 2468 7104 2496
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 9122 2496 9128 2508
rect 9083 2468 9128 2496
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 9309 2499 9367 2505
rect 9309 2465 9321 2499
rect 9355 2496 9367 2499
rect 10318 2496 10324 2508
rect 9355 2468 10324 2496
rect 9355 2465 9367 2468
rect 9309 2459 9367 2465
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10505 2499 10563 2505
rect 10505 2465 10517 2499
rect 10551 2465 10563 2499
rect 10505 2459 10563 2465
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 2792 2400 3801 2428
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 2792 2360 2820 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5166 2428 5172 2440
rect 5031 2400 5172 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 2648 2332 2820 2360
rect 6564 2360 6592 2391
rect 7466 2360 7472 2372
rect 6564 2332 7472 2360
rect 2648 2320 2654 2332
rect 7466 2320 7472 2332
rect 7524 2320 7530 2372
rect 9030 2320 9036 2372
rect 9088 2360 9094 2372
rect 10520 2360 10548 2459
rect 20714 2456 20720 2508
rect 20772 2496 20778 2508
rect 24596 2505 24624 2536
rect 25498 2524 25504 2536
rect 25556 2524 25562 2576
rect 25590 2524 25596 2576
rect 25648 2564 25654 2576
rect 44361 2567 44419 2573
rect 44361 2564 44373 2567
rect 25648 2536 44373 2564
rect 25648 2524 25654 2536
rect 44361 2533 44373 2536
rect 44407 2533 44419 2567
rect 44361 2527 44419 2533
rect 45278 2524 45284 2576
rect 45336 2524 45342 2576
rect 24581 2499 24639 2505
rect 20772 2468 22876 2496
rect 20772 2456 20778 2468
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15528 2400 15761 2428
rect 15528 2388 15534 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 17865 2431 17923 2437
rect 17865 2397 17877 2431
rect 17911 2428 17923 2431
rect 18322 2428 18328 2440
rect 17911 2400 18328 2428
rect 17911 2397 17923 2400
rect 17865 2391 17923 2397
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 18509 2431 18567 2437
rect 18509 2397 18521 2431
rect 18555 2428 18567 2431
rect 18598 2428 18604 2440
rect 18555 2400 18604 2428
rect 18555 2397 18567 2400
rect 18509 2391 18567 2397
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2428 20131 2431
rect 20990 2428 20996 2440
rect 20119 2400 20996 2428
rect 20119 2397 20131 2400
rect 20073 2391 20131 2397
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 22094 2428 22100 2440
rect 22055 2400 22100 2428
rect 22094 2388 22100 2400
rect 22152 2388 22158 2440
rect 22848 2437 22876 2468
rect 24581 2465 24593 2499
rect 24627 2465 24639 2499
rect 24762 2496 24768 2508
rect 24723 2468 24768 2496
rect 24581 2459 24639 2465
rect 24762 2456 24768 2468
rect 24820 2456 24826 2508
rect 25130 2496 25136 2508
rect 25091 2468 25136 2496
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 35802 2496 35808 2508
rect 35763 2468 35808 2496
rect 35802 2456 35808 2468
rect 35860 2456 35866 2508
rect 41325 2499 41383 2505
rect 41325 2465 41337 2499
rect 41371 2496 41383 2499
rect 41690 2496 41696 2508
rect 41371 2468 41696 2496
rect 41371 2465 41383 2468
rect 41325 2459 41383 2465
rect 41690 2456 41696 2468
rect 41748 2456 41754 2508
rect 42705 2499 42763 2505
rect 42705 2465 42717 2499
rect 42751 2496 42763 2499
rect 45094 2496 45100 2508
rect 42751 2468 45100 2496
rect 42751 2465 42763 2468
rect 42705 2459 42763 2465
rect 45094 2456 45100 2468
rect 45152 2456 45158 2508
rect 45189 2499 45247 2505
rect 45189 2465 45201 2499
rect 45235 2496 45247 2499
rect 45296 2496 45324 2524
rect 45235 2468 45324 2496
rect 45373 2499 45431 2505
rect 45235 2465 45247 2468
rect 45189 2459 45247 2465
rect 45373 2465 45385 2499
rect 45419 2496 45431 2499
rect 45738 2496 45744 2508
rect 45419 2468 45744 2496
rect 45419 2465 45431 2468
rect 45373 2459 45431 2465
rect 45738 2456 45744 2468
rect 45796 2456 45802 2508
rect 45830 2456 45836 2508
rect 45888 2496 45894 2508
rect 45888 2468 45933 2496
rect 45888 2456 45894 2468
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26476 2400 26985 2428
rect 26476 2388 26482 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 27249 2431 27307 2437
rect 27249 2397 27261 2431
rect 27295 2397 27307 2431
rect 27249 2391 27307 2397
rect 9088 2332 10548 2360
rect 9088 2320 9094 2332
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16172 2332 17141 2360
rect 16172 2320 16178 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 17129 2323 17187 2329
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 20809 2363 20867 2369
rect 20809 2360 20821 2363
rect 20680 2332 20821 2360
rect 20680 2320 20686 2332
rect 20809 2329 20821 2332
rect 20855 2329 20867 2363
rect 20809 2323 20867 2329
rect 24026 2320 24032 2372
rect 24084 2360 24090 2372
rect 27264 2360 27292 2391
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29696 2400 29929 2428
rect 29696 2388 29702 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35492 2400 35541 2428
rect 35492 2388 35498 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 38010 2388 38016 2440
rect 38068 2428 38074 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 38068 2400 38117 2428
rect 38068 2388 38074 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 39117 2431 39175 2437
rect 39117 2397 39129 2431
rect 39163 2428 39175 2431
rect 39574 2428 39580 2440
rect 39163 2400 39580 2428
rect 39163 2397 39175 2400
rect 39117 2391 39175 2397
rect 39574 2388 39580 2400
rect 39632 2388 39638 2440
rect 41049 2431 41107 2437
rect 41049 2397 41061 2431
rect 41095 2428 41107 2431
rect 41230 2428 41236 2440
rect 41095 2400 41236 2428
rect 41095 2397 41107 2400
rect 41049 2391 41107 2397
rect 41230 2388 41236 2400
rect 41288 2388 41294 2440
rect 42429 2431 42487 2437
rect 42429 2397 42441 2431
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 44177 2431 44235 2437
rect 44177 2397 44189 2431
rect 44223 2397 44235 2431
rect 44177 2391 44235 2397
rect 24084 2332 27292 2360
rect 24084 2320 24090 2332
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28537 2363 28595 2369
rect 28537 2360 28549 2363
rect 28408 2332 28549 2360
rect 28408 2320 28414 2332
rect 28537 2329 28549 2332
rect 28583 2329 28595 2363
rect 28537 2323 28595 2329
rect 29822 2320 29828 2372
rect 29880 2360 29886 2372
rect 29880 2332 38424 2360
rect 29880 2320 29886 2332
rect 3973 2295 4031 2301
rect 3973 2261 3985 2295
rect 4019 2292 4031 2295
rect 16850 2292 16856 2304
rect 4019 2264 16856 2292
rect 4019 2261 4031 2264
rect 3973 2255 4031 2261
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 29454 2252 29460 2304
rect 29512 2292 29518 2304
rect 38289 2295 38347 2301
rect 38289 2292 38301 2295
rect 29512 2264 38301 2292
rect 29512 2252 29518 2264
rect 38289 2261 38301 2264
rect 38335 2261 38347 2295
rect 38396 2292 38424 2332
rect 39298 2320 39304 2372
rect 39356 2360 39362 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39356 2332 40325 2360
rect 39356 2320 39362 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 42444 2360 42472 2391
rect 40644 2332 42472 2360
rect 44192 2360 44220 2391
rect 45462 2360 45468 2372
rect 44192 2332 45468 2360
rect 40644 2320 40650 2332
rect 45462 2320 45468 2332
rect 45520 2320 45526 2372
rect 47765 2363 47823 2369
rect 47765 2329 47777 2363
rect 47811 2360 47823 2363
rect 47946 2360 47952 2372
rect 47811 2332 47952 2360
rect 47811 2329 47823 2332
rect 47765 2323 47823 2329
rect 47946 2320 47952 2332
rect 48004 2320 48010 2372
rect 47857 2295 47915 2301
rect 47857 2292 47869 2295
rect 38396 2264 47869 2292
rect 38289 2255 38347 2261
rect 47857 2261 47869 2264
rect 47903 2261 47915 2295
rect 47857 2255 47915 2261
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 29276 47200 29328 47252
rect 19984 47132 20036 47184
rect 12256 47064 12308 47116
rect 13820 47064 13872 47116
rect 20076 47107 20128 47116
rect 20076 47073 20085 47107
rect 20085 47073 20119 47107
rect 20119 47073 20128 47107
rect 20076 47064 20128 47073
rect 20536 47064 20588 47116
rect 30748 47107 30800 47116
rect 30748 47073 30757 47107
rect 30757 47073 30791 47107
rect 30791 47073 30800 47107
rect 30748 47064 30800 47073
rect 45100 47064 45152 47116
rect 48320 47064 48372 47116
rect 1952 47039 2004 47048
rect 1952 47005 1961 47039
rect 1961 47005 1995 47039
rect 1995 47005 2004 47039
rect 1952 46996 2004 47005
rect 2596 46996 2648 47048
rect 3240 46996 3292 47048
rect 4804 47039 4856 47048
rect 4804 47005 4813 47039
rect 4813 47005 4847 47039
rect 4847 47005 4856 47039
rect 4804 46996 4856 47005
rect 5816 46996 5868 47048
rect 7104 46996 7156 47048
rect 9036 46996 9088 47048
rect 12624 47039 12676 47048
rect 12624 47005 12633 47039
rect 12633 47005 12667 47039
rect 12667 47005 12676 47039
rect 12624 46996 12676 47005
rect 14464 46996 14516 47048
rect 16488 46996 16540 47048
rect 4068 46971 4120 46980
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 5080 46928 5132 46980
rect 7840 46928 7892 46980
rect 9496 46928 9548 46980
rect 18696 46996 18748 47048
rect 20352 47039 20404 47048
rect 20352 47005 20361 47039
rect 20361 47005 20395 47039
rect 20395 47005 20404 47039
rect 20352 46996 20404 47005
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 30104 46996 30156 47048
rect 38108 46996 38160 47048
rect 42616 47039 42668 47048
rect 42616 47005 42625 47039
rect 42625 47005 42659 47039
rect 42659 47005 42668 47039
rect 42616 46996 42668 47005
rect 45192 47039 45244 47048
rect 45192 47005 45201 47039
rect 45201 47005 45235 47039
rect 45235 47005 45244 47039
rect 45192 46996 45244 47005
rect 47676 46996 47728 47048
rect 20168 46928 20220 46980
rect 2136 46903 2188 46912
rect 2136 46869 2145 46903
rect 2145 46869 2179 46903
rect 2179 46869 2188 46903
rect 2136 46860 2188 46869
rect 2872 46903 2924 46912
rect 2872 46869 2881 46903
rect 2881 46869 2915 46903
rect 2915 46869 2924 46903
rect 2872 46860 2924 46869
rect 6920 46903 6972 46912
rect 6920 46869 6929 46903
rect 6929 46869 6963 46903
rect 6963 46869 6972 46903
rect 29920 46903 29972 46912
rect 6920 46860 6972 46869
rect 29920 46869 29929 46903
rect 29929 46869 29963 46903
rect 29963 46869 29972 46903
rect 29920 46860 29972 46869
rect 39304 46860 39356 46912
rect 40408 46928 40460 46980
rect 43260 46928 43312 46980
rect 45468 46928 45520 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 2872 46588 2924 46640
rect 1400 46563 1452 46572
rect 1400 46529 1409 46563
rect 1409 46529 1443 46563
rect 1443 46529 1452 46563
rect 1400 46520 1452 46529
rect 11612 46520 11664 46572
rect 29276 46563 29328 46572
rect 29276 46529 29285 46563
rect 29285 46529 29319 46563
rect 29319 46529 29328 46563
rect 29276 46520 29328 46529
rect 38108 46563 38160 46572
rect 38108 46529 38117 46563
rect 38117 46529 38151 46563
rect 38151 46529 38160 46563
rect 38108 46520 38160 46529
rect 47860 46563 47912 46572
rect 47860 46529 47869 46563
rect 47869 46529 47903 46563
rect 47903 46529 47912 46563
rect 47860 46520 47912 46529
rect 3976 46495 4028 46504
rect 3976 46461 3985 46495
rect 3985 46461 4019 46495
rect 4019 46461 4028 46495
rect 3976 46452 4028 46461
rect 4988 46452 5040 46504
rect 3884 46384 3936 46436
rect 1676 46316 1728 46368
rect 2320 46359 2372 46368
rect 2320 46325 2329 46359
rect 2329 46325 2363 46359
rect 2363 46325 2372 46359
rect 2320 46316 2372 46325
rect 10600 46316 10652 46368
rect 14188 46452 14240 46504
rect 14280 46495 14332 46504
rect 14280 46461 14289 46495
rect 14289 46461 14323 46495
rect 14323 46461 14332 46495
rect 14280 46452 14332 46461
rect 19616 46495 19668 46504
rect 19616 46461 19625 46495
rect 19625 46461 19659 46495
rect 19659 46461 19668 46495
rect 19616 46452 19668 46461
rect 20628 46495 20680 46504
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 27620 46452 27672 46504
rect 20076 46384 20128 46436
rect 25780 46384 25832 46436
rect 37740 46452 37792 46504
rect 38384 46452 38436 46504
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 42616 46495 42668 46504
rect 42616 46461 42625 46495
rect 42625 46461 42659 46495
rect 42659 46461 42668 46495
rect 42616 46452 42668 46461
rect 45192 46495 45244 46504
rect 42524 46384 42576 46436
rect 45192 46461 45201 46495
rect 45201 46461 45235 46495
rect 45235 46461 45244 46495
rect 45192 46452 45244 46461
rect 45376 46495 45428 46504
rect 45376 46461 45385 46495
rect 45385 46461 45419 46495
rect 45419 46461 45428 46495
rect 45376 46452 45428 46461
rect 46848 46495 46900 46504
rect 46848 46461 46857 46495
rect 46857 46461 46891 46495
rect 46891 46461 46900 46495
rect 46848 46452 46900 46461
rect 17224 46316 17276 46368
rect 25228 46316 25280 46368
rect 31668 46316 31720 46368
rect 34520 46316 34572 46368
rect 39948 46316 40000 46368
rect 41328 46316 41380 46368
rect 44916 46316 44968 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3976 46112 4028 46164
rect 4988 46155 5040 46164
rect 4988 46121 4997 46155
rect 4997 46121 5031 46155
rect 5031 46121 5040 46155
rect 4988 46112 5040 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 19616 46112 19668 46164
rect 20076 46155 20128 46164
rect 20076 46121 20085 46155
rect 20085 46121 20119 46155
rect 20119 46121 20128 46155
rect 20076 46112 20128 46121
rect 27620 46155 27672 46164
rect 27620 46121 27629 46155
rect 27629 46121 27663 46155
rect 27663 46121 27672 46155
rect 27620 46112 27672 46121
rect 38384 46155 38436 46164
rect 38384 46121 38393 46155
rect 38393 46121 38427 46155
rect 38427 46121 38436 46155
rect 38384 46112 38436 46121
rect 38292 46044 38344 46096
rect 44180 46044 44232 46096
rect 2320 45976 2372 46028
rect 2780 46019 2832 46028
rect 2780 45985 2789 46019
rect 2789 45985 2823 46019
rect 2823 45985 2832 46019
rect 2780 45976 2832 45985
rect 10600 46019 10652 46028
rect 10600 45985 10609 46019
rect 10609 45985 10643 46019
rect 10643 45985 10652 46019
rect 10600 45976 10652 45985
rect 10968 45976 11020 46028
rect 21272 45976 21324 46028
rect 25228 46019 25280 46028
rect 25228 45985 25237 46019
rect 25237 45985 25271 46019
rect 25271 45985 25280 46019
rect 25228 45976 25280 45985
rect 25412 45976 25464 46028
rect 27068 45976 27120 46028
rect 27620 45976 27672 46028
rect 31668 46019 31720 46028
rect 31668 45985 31677 46019
rect 31677 45985 31711 46019
rect 31711 45985 31720 46019
rect 31668 45976 31720 45985
rect 32220 46019 32272 46028
rect 32220 45985 32229 46019
rect 32229 45985 32263 46019
rect 32263 45985 32272 46019
rect 32220 45976 32272 45985
rect 41328 46019 41380 46028
rect 41328 45985 41337 46019
rect 41337 45985 41371 46019
rect 41371 45985 41380 46019
rect 41328 45976 41380 45985
rect 41880 46019 41932 46028
rect 41880 45985 41889 46019
rect 41889 45985 41923 46019
rect 41923 45985 41932 46019
rect 41880 45976 41932 45985
rect 47032 46019 47084 46028
rect 47032 45985 47041 46019
rect 47041 45985 47075 46019
rect 47075 45985 47084 46019
rect 47032 45976 47084 45985
rect 4896 45951 4948 45960
rect 4896 45917 4905 45951
rect 4905 45917 4939 45951
rect 4939 45917 4948 45951
rect 4896 45908 4948 45917
rect 12900 45908 12952 45960
rect 14096 45951 14148 45960
rect 14096 45917 14105 45951
rect 14105 45917 14139 45951
rect 14139 45917 14148 45951
rect 14096 45908 14148 45917
rect 18972 45908 19024 45960
rect 20904 45951 20956 45960
rect 20904 45917 20913 45951
rect 20913 45917 20947 45951
rect 20947 45917 20956 45951
rect 20904 45908 20956 45917
rect 38292 45951 38344 45960
rect 2228 45840 2280 45892
rect 10784 45883 10836 45892
rect 10784 45849 10793 45883
rect 10793 45849 10827 45883
rect 10827 45849 10836 45883
rect 10784 45840 10836 45849
rect 21088 45883 21140 45892
rect 21088 45849 21097 45883
rect 21097 45849 21131 45883
rect 21131 45849 21140 45883
rect 21088 45840 21140 45849
rect 25412 45883 25464 45892
rect 25412 45849 25421 45883
rect 25421 45849 25455 45883
rect 25455 45849 25464 45883
rect 25412 45840 25464 45849
rect 20996 45772 21048 45824
rect 38292 45917 38301 45951
rect 38301 45917 38335 45951
rect 38335 45917 38344 45951
rect 38292 45908 38344 45917
rect 43812 45908 43864 45960
rect 45744 45908 45796 45960
rect 46296 45951 46348 45960
rect 46296 45917 46305 45951
rect 46305 45917 46339 45951
rect 46339 45917 46348 45951
rect 46296 45908 46348 45917
rect 32220 45840 32272 45892
rect 41512 45883 41564 45892
rect 41512 45849 41521 45883
rect 41521 45849 41555 45883
rect 41555 45849 41564 45883
rect 41512 45840 41564 45849
rect 46480 45883 46532 45892
rect 46480 45849 46489 45883
rect 46489 45849 46523 45883
rect 46523 45849 46532 45883
rect 46480 45840 46532 45849
rect 41696 45772 41748 45824
rect 43996 45772 44048 45824
rect 45744 45815 45796 45824
rect 45744 45781 45753 45815
rect 45753 45781 45787 45815
rect 45787 45781 45796 45815
rect 45744 45772 45796 45781
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 2228 45611 2280 45620
rect 2228 45577 2237 45611
rect 2237 45577 2271 45611
rect 2271 45577 2280 45611
rect 2228 45568 2280 45577
rect 10784 45611 10836 45620
rect 10784 45577 10793 45611
rect 10793 45577 10827 45611
rect 10827 45577 10836 45611
rect 10784 45568 10836 45577
rect 32220 45611 32272 45620
rect 32220 45577 32229 45611
rect 32229 45577 32263 45611
rect 32263 45577 32272 45611
rect 32220 45568 32272 45577
rect 42616 45568 42668 45620
rect 46480 45568 46532 45620
rect 41512 45500 41564 45552
rect 2412 45432 2464 45484
rect 20904 45432 20956 45484
rect 32128 45475 32180 45484
rect 25780 45364 25832 45416
rect 32128 45441 32137 45475
rect 32137 45441 32171 45475
rect 32171 45441 32180 45475
rect 32128 45432 32180 45441
rect 41052 45475 41104 45484
rect 41052 45441 41061 45475
rect 41061 45441 41095 45475
rect 41095 45441 41104 45475
rect 41696 45475 41748 45484
rect 41052 45432 41104 45441
rect 41696 45441 41705 45475
rect 41705 45441 41739 45475
rect 41739 45441 41748 45475
rect 41696 45432 41748 45441
rect 45836 45475 45888 45484
rect 4896 45296 4948 45348
rect 42432 45364 42484 45416
rect 42616 45407 42668 45416
rect 42616 45373 42625 45407
rect 42625 45373 42659 45407
rect 42659 45373 42668 45407
rect 42616 45364 42668 45373
rect 42800 45407 42852 45416
rect 42800 45373 42809 45407
rect 42809 45373 42843 45407
rect 42843 45373 42852 45407
rect 42800 45364 42852 45373
rect 43168 45407 43220 45416
rect 43168 45373 43177 45407
rect 43177 45373 43211 45407
rect 43211 45373 43220 45407
rect 43168 45364 43220 45373
rect 45836 45441 45845 45475
rect 45845 45441 45879 45475
rect 45879 45441 45888 45475
rect 45836 45432 45888 45441
rect 46388 45500 46440 45552
rect 46480 45432 46532 45484
rect 47308 45432 47360 45484
rect 46940 45364 46992 45416
rect 41052 45296 41104 45348
rect 46756 45296 46808 45348
rect 45100 45271 45152 45280
rect 45100 45237 45109 45271
rect 45109 45237 45143 45271
rect 45143 45237 45152 45271
rect 45100 45228 45152 45237
rect 45928 45228 45980 45280
rect 47676 45271 47728 45280
rect 47676 45237 47685 45271
rect 47685 45237 47719 45271
rect 47719 45237 47728 45271
rect 47676 45228 47728 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 21088 45024 21140 45076
rect 42800 45024 42852 45076
rect 43260 45067 43312 45076
rect 43260 45033 43269 45067
rect 43269 45033 43303 45067
rect 43303 45033 43312 45067
rect 43260 45024 43312 45033
rect 45192 45024 45244 45076
rect 45836 45024 45888 45076
rect 47400 45024 47452 45076
rect 25412 44956 25464 45008
rect 45100 44956 45152 45008
rect 42432 44888 42484 44940
rect 47676 44888 47728 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 21824 44820 21876 44872
rect 25780 44820 25832 44872
rect 43168 44863 43220 44872
rect 24676 44684 24728 44736
rect 43168 44829 43177 44863
rect 43177 44829 43211 44863
rect 43211 44829 43220 44863
rect 43168 44820 43220 44829
rect 44456 44820 44508 44872
rect 46020 44752 46072 44804
rect 47032 44752 47084 44804
rect 47584 44684 47636 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 45376 44480 45428 44532
rect 45468 44480 45520 44532
rect 24676 44455 24728 44464
rect 24676 44421 24685 44455
rect 24685 44421 24719 44455
rect 24719 44421 24728 44455
rect 24676 44412 24728 44421
rect 21824 44344 21876 44396
rect 42616 44344 42668 44396
rect 44180 44344 44232 44396
rect 46296 44344 46348 44396
rect 47308 44344 47360 44396
rect 24492 44319 24544 44328
rect 24492 44285 24501 44319
rect 24501 44285 24535 44319
rect 24535 44285 24544 44319
rect 24492 44276 24544 44285
rect 2964 44208 3016 44260
rect 42708 44276 42760 44328
rect 24584 44140 24636 44192
rect 47676 44183 47728 44192
rect 47676 44149 47685 44183
rect 47685 44149 47719 44183
rect 47719 44149 47728 44183
rect 47676 44140 47728 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 24584 43843 24636 43852
rect 24584 43809 24593 43843
rect 24593 43809 24627 43843
rect 24627 43809 24636 43843
rect 24584 43800 24636 43809
rect 34520 43800 34572 43852
rect 47676 43800 47728 43852
rect 48228 43800 48280 43852
rect 23480 43732 23532 43784
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1860 43299 1912 43308
rect 1860 43265 1869 43299
rect 1869 43265 1903 43299
rect 1903 43265 1912 43299
rect 1860 43256 1912 43265
rect 45284 43256 45336 43308
rect 47032 43299 47084 43308
rect 47032 43265 47041 43299
rect 47041 43265 47075 43299
rect 47075 43265 47084 43299
rect 47032 43256 47084 43265
rect 1952 43095 2004 43104
rect 1952 43061 1961 43095
rect 1961 43061 1995 43095
rect 1995 43061 2004 43095
rect 1952 43052 2004 43061
rect 47768 43095 47820 43104
rect 47768 43061 47777 43095
rect 47777 43061 47811 43095
rect 47811 43061 47820 43095
rect 47768 43052 47820 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 47768 42712 47820 42764
rect 47676 42576 47728 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 47676 42347 47728 42356
rect 47676 42313 47685 42347
rect 47685 42313 47719 42347
rect 47719 42313 47728 42347
rect 47676 42304 47728 42313
rect 47124 42168 47176 42220
rect 47584 42211 47636 42220
rect 47584 42177 47593 42211
rect 47593 42177 47627 42211
rect 47627 42177 47636 42211
rect 47584 42168 47636 42177
rect 1400 41964 1452 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 27620 41667 27672 41676
rect 27620 41633 27629 41667
rect 27629 41633 27663 41667
rect 27663 41633 27672 41667
rect 27620 41624 27672 41633
rect 47768 41624 47820 41676
rect 25780 41599 25832 41608
rect 25780 41565 25789 41599
rect 25789 41565 25823 41599
rect 25823 41565 25832 41599
rect 25780 41556 25832 41565
rect 26424 41599 26476 41608
rect 26424 41565 26433 41599
rect 26433 41565 26467 41599
rect 26467 41565 26476 41599
rect 26424 41556 26476 41565
rect 48136 41599 48188 41608
rect 48136 41565 48145 41599
rect 48145 41565 48179 41599
rect 48179 41565 48188 41599
rect 48136 41556 48188 41565
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 46940 41488 46992 41540
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 46940 41259 46992 41268
rect 46940 41225 46949 41259
rect 46949 41225 46983 41259
rect 46983 41225 46992 41259
rect 46940 41216 46992 41225
rect 14096 41080 14148 41132
rect 46572 41080 46624 41132
rect 47768 41123 47820 41132
rect 47768 41089 47777 41123
rect 47777 41089 47811 41123
rect 47811 41089 47820 41123
rect 47768 41080 47820 41089
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 26424 40604 26476 40656
rect 1400 40511 1452 40520
rect 1400 40477 1409 40511
rect 1409 40477 1443 40511
rect 1443 40477 1452 40511
rect 1400 40468 1452 40477
rect 46112 40511 46164 40520
rect 2136 40400 2188 40452
rect 27436 40443 27488 40452
rect 27436 40409 27445 40443
rect 27445 40409 27479 40443
rect 27479 40409 27488 40443
rect 27436 40400 27488 40409
rect 46112 40477 46121 40511
rect 46121 40477 46155 40511
rect 46155 40477 46164 40511
rect 46112 40468 46164 40477
rect 47676 40511 47728 40520
rect 47676 40477 47685 40511
rect 47685 40477 47719 40511
rect 47719 40477 47728 40511
rect 47676 40468 47728 40477
rect 46204 40400 46256 40452
rect 10968 40332 11020 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 48044 40060 48096 40112
rect 46112 39992 46164 40044
rect 46756 40035 46808 40044
rect 46756 40001 46765 40035
rect 46765 40001 46799 40035
rect 46799 40001 46808 40035
rect 46756 39992 46808 40001
rect 44732 39967 44784 39976
rect 44732 39933 44741 39967
rect 44741 39933 44775 39967
rect 44775 39933 44784 39967
rect 44732 39924 44784 39933
rect 46480 39788 46532 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 47676 39516 47728 39568
rect 46480 39491 46532 39500
rect 46480 39457 46489 39491
rect 46489 39457 46523 39491
rect 46523 39457 46532 39491
rect 46480 39448 46532 39457
rect 48228 39448 48280 39500
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 20536 39083 20588 39092
rect 20536 39049 20545 39083
rect 20545 39049 20579 39083
rect 20579 39049 20588 39083
rect 20536 39040 20588 39049
rect 20628 38879 20680 38888
rect 20628 38845 20637 38879
rect 20637 38845 20671 38879
rect 20671 38845 20680 38879
rect 20628 38836 20680 38845
rect 45744 38904 45796 38956
rect 47032 38904 47084 38956
rect 47308 38904 47360 38956
rect 47768 38947 47820 38956
rect 47768 38913 47777 38947
rect 47777 38913 47811 38947
rect 47811 38913 47820 38947
rect 47768 38904 47820 38913
rect 25044 38879 25096 38888
rect 25044 38845 25053 38879
rect 25053 38845 25087 38879
rect 25087 38845 25096 38879
rect 25044 38836 25096 38845
rect 22008 38768 22060 38820
rect 45652 38768 45704 38820
rect 19524 38700 19576 38752
rect 23756 38743 23808 38752
rect 23756 38709 23765 38743
rect 23765 38709 23799 38743
rect 23799 38709 23808 38743
rect 23756 38700 23808 38709
rect 46940 38743 46992 38752
rect 46940 38709 46949 38743
rect 46949 38709 46983 38743
rect 46983 38709 46992 38743
rect 46940 38700 46992 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 25044 38496 25096 38548
rect 18328 38360 18380 38412
rect 21272 38360 21324 38412
rect 23940 38360 23992 38412
rect 46940 38360 46992 38412
rect 48136 38403 48188 38412
rect 48136 38369 48145 38403
rect 48145 38369 48179 38403
rect 48179 38369 48188 38403
rect 48136 38360 48188 38369
rect 23204 38335 23256 38344
rect 23204 38301 23213 38335
rect 23213 38301 23247 38335
rect 23247 38301 23256 38335
rect 23204 38292 23256 38301
rect 19524 38267 19576 38276
rect 19524 38233 19533 38267
rect 19533 38233 19567 38267
rect 19567 38233 19576 38267
rect 19524 38224 19576 38233
rect 20260 38224 20312 38276
rect 45836 38292 45888 38344
rect 24676 38224 24728 38276
rect 16856 38156 16908 38208
rect 17500 38199 17552 38208
rect 17500 38165 17509 38199
rect 17509 38165 17543 38199
rect 17543 38165 17552 38199
rect 17500 38156 17552 38165
rect 17592 38199 17644 38208
rect 17592 38165 17601 38199
rect 17601 38165 17635 38199
rect 17635 38165 17644 38199
rect 17592 38156 17644 38165
rect 19248 38156 19300 38208
rect 23296 38199 23348 38208
rect 23296 38165 23305 38199
rect 23305 38165 23339 38199
rect 23339 38165 23348 38199
rect 23296 38156 23348 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 17592 37995 17644 38004
rect 17592 37961 17601 37995
rect 17601 37961 17635 37995
rect 17635 37961 17644 37995
rect 17592 37952 17644 37961
rect 20260 37995 20312 38004
rect 20260 37961 20269 37995
rect 20269 37961 20303 37995
rect 20303 37961 20312 37995
rect 20260 37952 20312 37961
rect 22376 37952 22428 38004
rect 23204 37952 23256 38004
rect 17224 37884 17276 37936
rect 15292 37816 15344 37868
rect 16856 37859 16908 37868
rect 16856 37825 16865 37859
rect 16865 37825 16899 37859
rect 16899 37825 16908 37859
rect 16856 37816 16908 37825
rect 18052 37791 18104 37800
rect 18052 37757 18061 37791
rect 18061 37757 18095 37791
rect 18095 37757 18104 37791
rect 18052 37748 18104 37757
rect 18696 37816 18748 37868
rect 19248 37816 19300 37868
rect 20536 37816 20588 37868
rect 20996 37859 21048 37868
rect 20996 37825 21005 37859
rect 21005 37825 21039 37859
rect 21039 37825 21048 37859
rect 20996 37816 21048 37825
rect 21548 37816 21600 37868
rect 23296 37884 23348 37936
rect 22284 37816 22336 37868
rect 47584 37859 47636 37868
rect 47584 37825 47593 37859
rect 47593 37825 47627 37859
rect 47627 37825 47636 37859
rect 47584 37816 47636 37825
rect 15844 37680 15896 37732
rect 19340 37680 19392 37732
rect 20628 37748 20680 37800
rect 21272 37748 21324 37800
rect 23756 37748 23808 37800
rect 16580 37612 16632 37664
rect 21364 37612 21416 37664
rect 22008 37655 22060 37664
rect 22008 37621 22017 37655
rect 22017 37621 22051 37655
rect 22051 37621 22060 37655
rect 22008 37612 22060 37621
rect 24676 37655 24728 37664
rect 24676 37621 24685 37655
rect 24685 37621 24719 37655
rect 24719 37621 24728 37655
rect 24676 37612 24728 37621
rect 47032 37655 47084 37664
rect 47032 37621 47041 37655
rect 47041 37621 47075 37655
rect 47075 37621 47084 37655
rect 47032 37612 47084 37621
rect 47676 37655 47728 37664
rect 47676 37621 47685 37655
rect 47685 37621 47719 37655
rect 47719 37621 47728 37655
rect 47676 37612 47728 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 17500 37408 17552 37460
rect 18052 37408 18104 37460
rect 15844 37315 15896 37324
rect 15844 37281 15853 37315
rect 15853 37281 15887 37315
rect 15887 37281 15896 37315
rect 15844 37272 15896 37281
rect 18052 37315 18104 37324
rect 18052 37281 18061 37315
rect 18061 37281 18095 37315
rect 18095 37281 18104 37315
rect 18052 37272 18104 37281
rect 48136 37315 48188 37324
rect 48136 37281 48145 37315
rect 48145 37281 48179 37315
rect 48179 37281 48188 37315
rect 48136 37272 48188 37281
rect 1768 37204 1820 37256
rect 14188 37204 14240 37256
rect 17500 37204 17552 37256
rect 20536 37247 20588 37256
rect 20536 37213 20545 37247
rect 20545 37213 20579 37247
rect 20579 37213 20588 37247
rect 20536 37204 20588 37213
rect 16580 37136 16632 37188
rect 20904 37204 20956 37256
rect 21272 37247 21324 37256
rect 21272 37213 21281 37247
rect 21281 37213 21315 37247
rect 21315 37213 21324 37247
rect 21272 37204 21324 37213
rect 22652 37204 22704 37256
rect 12624 37068 12676 37120
rect 20536 37068 20588 37120
rect 22928 37068 22980 37120
rect 23112 37068 23164 37120
rect 28448 37204 28500 37256
rect 25780 37179 25832 37188
rect 25780 37145 25789 37179
rect 25789 37145 25823 37179
rect 25823 37145 25832 37179
rect 25780 37136 25832 37145
rect 27068 37136 27120 37188
rect 27896 37136 27948 37188
rect 27252 37111 27304 37120
rect 27252 37077 27261 37111
rect 27261 37077 27295 37111
rect 27295 37077 27304 37111
rect 28632 37111 28684 37120
rect 27252 37068 27304 37077
rect 28632 37077 28641 37111
rect 28641 37077 28675 37111
rect 28675 37077 28684 37111
rect 28632 37068 28684 37077
rect 47676 37136 47728 37188
rect 47032 37068 47084 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 9496 36864 9548 36916
rect 15200 36796 15252 36848
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 2228 36660 2280 36712
rect 2780 36703 2832 36712
rect 2780 36669 2789 36703
rect 2789 36669 2823 36703
rect 2823 36669 2832 36703
rect 2780 36660 2832 36669
rect 14188 36660 14240 36712
rect 16488 36660 16540 36712
rect 16028 36592 16080 36644
rect 17500 36728 17552 36780
rect 18052 36660 18104 36712
rect 18604 36660 18656 36712
rect 22652 36907 22704 36916
rect 21548 36728 21600 36780
rect 22652 36873 22661 36907
rect 22661 36873 22695 36907
rect 22695 36873 22704 36907
rect 22652 36864 22704 36873
rect 22928 36864 22980 36916
rect 23388 36864 23440 36916
rect 25320 36864 25372 36916
rect 25780 36907 25832 36916
rect 25780 36873 25789 36907
rect 25789 36873 25823 36907
rect 25823 36873 25832 36907
rect 25780 36864 25832 36873
rect 27068 36907 27120 36916
rect 27068 36873 27077 36907
rect 27077 36873 27111 36907
rect 27111 36873 27120 36907
rect 27068 36864 27120 36873
rect 25688 36796 25740 36848
rect 23112 36728 23164 36780
rect 23664 36660 23716 36712
rect 23940 36660 23992 36712
rect 24860 36728 24912 36780
rect 24952 36771 25004 36780
rect 24952 36737 24961 36771
rect 24961 36737 24995 36771
rect 24995 36737 25004 36771
rect 24952 36728 25004 36737
rect 26148 36728 26200 36780
rect 28448 36796 28500 36848
rect 28632 36796 28684 36848
rect 27896 36771 27948 36780
rect 27896 36737 27905 36771
rect 27905 36737 27939 36771
rect 27939 36737 27948 36771
rect 27896 36728 27948 36737
rect 26056 36660 26108 36712
rect 28172 36703 28224 36712
rect 25044 36592 25096 36644
rect 28172 36669 28181 36703
rect 28181 36669 28215 36703
rect 28215 36669 28224 36703
rect 28172 36660 28224 36669
rect 17408 36524 17460 36576
rect 18420 36524 18472 36576
rect 18604 36524 18656 36576
rect 23388 36524 23440 36576
rect 23572 36524 23624 36576
rect 23940 36524 23992 36576
rect 27712 36592 27764 36644
rect 25964 36524 26016 36576
rect 27988 36524 28040 36576
rect 28816 36524 28868 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2228 36363 2280 36372
rect 2228 36329 2237 36363
rect 2237 36329 2271 36363
rect 2271 36329 2280 36363
rect 2228 36320 2280 36329
rect 15200 36363 15252 36372
rect 15200 36329 15209 36363
rect 15209 36329 15243 36363
rect 15243 36329 15252 36363
rect 15200 36320 15252 36329
rect 15568 36320 15620 36372
rect 16488 36363 16540 36372
rect 10968 36252 11020 36304
rect 16488 36329 16497 36363
rect 16497 36329 16531 36363
rect 16531 36329 16540 36363
rect 16488 36320 16540 36329
rect 15568 36184 15620 36236
rect 16028 36227 16080 36236
rect 2228 36116 2280 36168
rect 15292 36116 15344 36168
rect 16028 36193 16037 36227
rect 16037 36193 16071 36227
rect 16071 36193 16080 36227
rect 16028 36184 16080 36193
rect 22560 36252 22612 36304
rect 23664 36320 23716 36372
rect 25780 36320 25832 36372
rect 25964 36363 26016 36372
rect 25964 36329 25973 36363
rect 25973 36329 26007 36363
rect 26007 36329 26016 36363
rect 25964 36320 26016 36329
rect 28172 36320 28224 36372
rect 23572 36252 23624 36304
rect 27804 36252 27856 36304
rect 29184 36252 29236 36304
rect 16488 36184 16540 36236
rect 17408 36227 17460 36236
rect 16212 36116 16264 36168
rect 17040 36116 17092 36168
rect 17408 36193 17417 36227
rect 17417 36193 17451 36227
rect 17451 36193 17460 36227
rect 17408 36184 17460 36193
rect 23112 36227 23164 36236
rect 18328 36116 18380 36168
rect 19064 36116 19116 36168
rect 23112 36193 23121 36227
rect 23121 36193 23155 36227
rect 23155 36193 23164 36227
rect 23112 36184 23164 36193
rect 20260 36159 20312 36168
rect 15292 35980 15344 36032
rect 16488 35980 16540 36032
rect 19984 36048 20036 36100
rect 20260 36125 20269 36159
rect 20269 36125 20303 36159
rect 20303 36125 20312 36159
rect 20260 36116 20312 36125
rect 23572 36159 23624 36168
rect 23572 36125 23581 36159
rect 23581 36125 23615 36159
rect 23615 36125 23624 36159
rect 23572 36116 23624 36125
rect 25044 36184 25096 36236
rect 24860 36116 24912 36168
rect 20536 36048 20588 36100
rect 21916 36048 21968 36100
rect 19432 35980 19484 36032
rect 24952 36048 25004 36100
rect 23388 35980 23440 36032
rect 23756 35980 23808 36032
rect 24768 36023 24820 36032
rect 24768 35989 24777 36023
rect 24777 35989 24811 36023
rect 24811 35989 24820 36023
rect 24768 35980 24820 35989
rect 25872 36159 25924 36168
rect 25872 36125 25881 36159
rect 25881 36125 25915 36159
rect 25915 36125 25924 36159
rect 26056 36159 26108 36168
rect 25872 36116 25924 36125
rect 26056 36125 26065 36159
rect 26065 36125 26099 36159
rect 26099 36125 26108 36159
rect 26056 36116 26108 36125
rect 27804 36116 27856 36168
rect 27988 36159 28040 36168
rect 27988 36125 27997 36159
rect 27997 36125 28031 36159
rect 28031 36125 28040 36159
rect 27988 36116 28040 36125
rect 28172 36048 28224 36100
rect 27252 35980 27304 36032
rect 28080 35980 28132 36032
rect 28448 36116 28500 36168
rect 29644 36023 29696 36032
rect 29644 35989 29653 36023
rect 29653 35989 29687 36023
rect 29687 35989 29696 36023
rect 29644 35980 29696 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 20628 35776 20680 35828
rect 24124 35819 24176 35828
rect 19432 35708 19484 35760
rect 19984 35708 20036 35760
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 16396 35640 16448 35692
rect 24124 35785 24133 35819
rect 24133 35785 24167 35819
rect 24167 35785 24176 35819
rect 24124 35776 24176 35785
rect 23756 35751 23808 35760
rect 23756 35717 23765 35751
rect 23765 35717 23799 35751
rect 23799 35717 23808 35751
rect 23756 35708 23808 35717
rect 26424 35708 26476 35760
rect 24768 35683 24820 35692
rect 14188 35572 14240 35624
rect 20720 35572 20772 35624
rect 21272 35572 21324 35624
rect 24768 35649 24777 35683
rect 24777 35649 24811 35683
rect 24811 35649 24820 35683
rect 24768 35640 24820 35649
rect 25688 35640 25740 35692
rect 27896 35708 27948 35760
rect 29644 35708 29696 35760
rect 31300 35640 31352 35692
rect 24860 35572 24912 35624
rect 28356 35572 28408 35624
rect 1492 35436 1544 35488
rect 15476 35436 15528 35488
rect 20812 35479 20864 35488
rect 20812 35445 20821 35479
rect 20821 35445 20855 35479
rect 20855 35445 20864 35479
rect 23940 35479 23992 35488
rect 20812 35436 20864 35445
rect 23940 35445 23949 35479
rect 23949 35445 23983 35479
rect 23983 35445 23992 35479
rect 23940 35436 23992 35445
rect 25964 35436 26016 35488
rect 27712 35436 27764 35488
rect 28264 35436 28316 35488
rect 28908 35436 28960 35488
rect 31208 35436 31260 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 18880 35232 18932 35284
rect 20536 35275 20588 35284
rect 20260 35164 20312 35216
rect 20536 35241 20545 35275
rect 20545 35241 20579 35275
rect 20579 35241 20588 35275
rect 20536 35232 20588 35241
rect 20904 35164 20956 35216
rect 27528 35232 27580 35284
rect 28172 35232 28224 35284
rect 18328 35096 18380 35148
rect 14188 35071 14240 35080
rect 14188 35037 14197 35071
rect 14197 35037 14231 35071
rect 14231 35037 14240 35071
rect 14188 35028 14240 35037
rect 20996 35096 21048 35148
rect 27896 35096 27948 35148
rect 43996 35096 44048 35148
rect 14464 35003 14516 35012
rect 14464 34969 14473 35003
rect 14473 34969 14507 35003
rect 14507 34969 14516 35003
rect 14464 34960 14516 34969
rect 15476 34960 15528 35012
rect 15844 34892 15896 34944
rect 18512 34960 18564 35012
rect 19340 34960 19392 35012
rect 20812 35071 20864 35080
rect 20812 35037 20821 35071
rect 20821 35037 20855 35071
rect 20855 35037 20864 35071
rect 20812 35028 20864 35037
rect 21180 35028 21232 35080
rect 22376 35071 22428 35080
rect 22376 35037 22385 35071
rect 22385 35037 22419 35071
rect 22419 35037 22428 35071
rect 22376 35028 22428 35037
rect 27804 35071 27856 35080
rect 27804 35037 27813 35071
rect 27813 35037 27847 35071
rect 27847 35037 27856 35071
rect 27804 35028 27856 35037
rect 28172 35071 28224 35080
rect 28172 35037 28181 35071
rect 28181 35037 28215 35071
rect 28215 35037 28224 35071
rect 28172 35028 28224 35037
rect 48136 35071 48188 35080
rect 48136 35037 48145 35071
rect 48145 35037 48179 35071
rect 48179 35037 48188 35071
rect 48136 35028 48188 35037
rect 22652 34960 22704 35012
rect 25228 34960 25280 35012
rect 25964 34960 26016 35012
rect 26240 34960 26292 35012
rect 29092 34960 29144 35012
rect 30472 35003 30524 35012
rect 30472 34969 30481 35003
rect 30481 34969 30515 35003
rect 30515 34969 30524 35003
rect 30472 34960 30524 34969
rect 31208 34960 31260 35012
rect 17684 34892 17736 34944
rect 22560 34892 22612 34944
rect 25596 34892 25648 34944
rect 27252 34935 27304 34944
rect 27252 34901 27261 34935
rect 27261 34901 27295 34935
rect 27295 34901 27304 34935
rect 27252 34892 27304 34901
rect 28080 34892 28132 34944
rect 28264 34892 28316 34944
rect 30012 34892 30064 34944
rect 30196 34892 30248 34944
rect 47124 34892 47176 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 14464 34688 14516 34740
rect 18512 34688 18564 34740
rect 15476 34552 15528 34604
rect 15844 34552 15896 34604
rect 16120 34552 16172 34604
rect 15752 34527 15804 34536
rect 15752 34493 15761 34527
rect 15761 34493 15795 34527
rect 15795 34493 15804 34527
rect 17960 34620 18012 34672
rect 17408 34595 17460 34604
rect 17408 34561 17417 34595
rect 17417 34561 17451 34595
rect 17451 34561 17460 34595
rect 17408 34552 17460 34561
rect 17684 34595 17736 34604
rect 17684 34561 17693 34595
rect 17693 34561 17727 34595
rect 17727 34561 17736 34595
rect 17684 34552 17736 34561
rect 18512 34527 18564 34536
rect 15752 34484 15804 34493
rect 18512 34493 18521 34527
rect 18521 34493 18555 34527
rect 18555 34493 18564 34527
rect 18512 34484 18564 34493
rect 18696 34595 18748 34604
rect 18696 34561 18705 34595
rect 18705 34561 18739 34595
rect 18739 34561 18748 34595
rect 19340 34595 19392 34604
rect 18696 34552 18748 34561
rect 19340 34561 19349 34595
rect 19349 34561 19383 34595
rect 19383 34561 19392 34595
rect 19340 34552 19392 34561
rect 20904 34688 20956 34740
rect 23572 34688 23624 34740
rect 24860 34688 24912 34740
rect 25044 34688 25096 34740
rect 26884 34688 26936 34740
rect 30472 34688 30524 34740
rect 22560 34620 22612 34672
rect 24768 34620 24820 34672
rect 20720 34552 20772 34604
rect 24676 34595 24728 34604
rect 24676 34561 24685 34595
rect 24685 34561 24719 34595
rect 24719 34561 24728 34595
rect 24676 34552 24728 34561
rect 25596 34595 25648 34604
rect 22100 34527 22152 34536
rect 22100 34493 22109 34527
rect 22109 34493 22143 34527
rect 22143 34493 22152 34527
rect 22100 34484 22152 34493
rect 25596 34561 25605 34595
rect 25605 34561 25639 34595
rect 25639 34561 25648 34595
rect 25596 34552 25648 34561
rect 27620 34595 27672 34604
rect 27620 34561 27629 34595
rect 27629 34561 27663 34595
rect 27663 34561 27672 34595
rect 27620 34552 27672 34561
rect 27712 34552 27764 34604
rect 27988 34620 28040 34672
rect 28908 34620 28960 34672
rect 28080 34552 28132 34604
rect 28356 34595 28408 34604
rect 28356 34561 28365 34595
rect 28365 34561 28399 34595
rect 28399 34561 28408 34595
rect 28356 34552 28408 34561
rect 30012 34620 30064 34672
rect 25412 34527 25464 34536
rect 25412 34493 25421 34527
rect 25421 34493 25455 34527
rect 25455 34493 25464 34527
rect 25412 34484 25464 34493
rect 28724 34484 28776 34536
rect 18052 34416 18104 34468
rect 19064 34416 19116 34468
rect 20996 34416 21048 34468
rect 17868 34348 17920 34400
rect 18144 34348 18196 34400
rect 23572 34391 23624 34400
rect 23572 34357 23581 34391
rect 23581 34357 23615 34391
rect 23615 34357 23624 34391
rect 23572 34348 23624 34357
rect 25596 34416 25648 34468
rect 30196 34552 30248 34604
rect 31116 34595 31168 34604
rect 31116 34561 31125 34595
rect 31125 34561 31159 34595
rect 31159 34561 31168 34595
rect 31116 34552 31168 34561
rect 48136 34595 48188 34604
rect 48136 34561 48145 34595
rect 48145 34561 48179 34595
rect 48179 34561 48188 34595
rect 48136 34552 48188 34561
rect 29000 34527 29052 34536
rect 29000 34493 29009 34527
rect 29009 34493 29043 34527
rect 29043 34493 29052 34527
rect 29000 34484 29052 34493
rect 30012 34527 30064 34536
rect 30012 34493 30021 34527
rect 30021 34493 30055 34527
rect 30055 34493 30064 34527
rect 30012 34484 30064 34493
rect 29368 34416 29420 34468
rect 24860 34391 24912 34400
rect 24860 34357 24869 34391
rect 24869 34357 24903 34391
rect 24903 34357 24912 34391
rect 24860 34348 24912 34357
rect 25320 34391 25372 34400
rect 25320 34357 25329 34391
rect 25329 34357 25363 34391
rect 25363 34357 25372 34391
rect 25320 34348 25372 34357
rect 28816 34391 28868 34400
rect 28816 34357 28825 34391
rect 28825 34357 28859 34391
rect 28859 34357 28868 34391
rect 28816 34348 28868 34357
rect 47216 34348 47268 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 17408 34144 17460 34196
rect 18236 34187 18288 34196
rect 18236 34153 18245 34187
rect 18245 34153 18279 34187
rect 18279 34153 18288 34187
rect 18236 34144 18288 34153
rect 22100 34144 22152 34196
rect 22652 34187 22704 34196
rect 22652 34153 22661 34187
rect 22661 34153 22695 34187
rect 22695 34153 22704 34187
rect 22652 34144 22704 34153
rect 24860 34144 24912 34196
rect 25228 34144 25280 34196
rect 27620 34144 27672 34196
rect 28172 34144 28224 34196
rect 31116 34144 31168 34196
rect 16212 34008 16264 34060
rect 1308 33940 1360 33992
rect 14188 33983 14240 33992
rect 14188 33949 14197 33983
rect 14197 33949 14231 33983
rect 14231 33949 14240 33983
rect 14188 33940 14240 33949
rect 16396 33983 16448 33992
rect 16396 33949 16405 33983
rect 16405 33949 16439 33983
rect 16439 33949 16448 33983
rect 16396 33940 16448 33949
rect 14464 33915 14516 33924
rect 14464 33881 14473 33915
rect 14473 33881 14507 33915
rect 14507 33881 14516 33915
rect 14464 33872 14516 33881
rect 1584 33804 1636 33856
rect 16396 33804 16448 33856
rect 17960 34008 18012 34060
rect 18420 34008 18472 34060
rect 18972 34008 19024 34060
rect 17040 33940 17092 33992
rect 17224 33940 17276 33992
rect 18052 33983 18104 33992
rect 18052 33949 18061 33983
rect 18061 33949 18095 33983
rect 18095 33949 18104 33983
rect 18052 33940 18104 33949
rect 19064 33940 19116 33992
rect 20168 34008 20220 34060
rect 25044 34076 25096 34128
rect 27252 34076 27304 34128
rect 27988 34076 28040 34128
rect 29092 34076 29144 34128
rect 21272 33983 21324 33992
rect 21272 33949 21281 33983
rect 21281 33949 21315 33983
rect 21315 33949 21324 33983
rect 21272 33940 21324 33949
rect 21456 33983 21508 33992
rect 19340 33804 19392 33856
rect 20260 33872 20312 33924
rect 21456 33949 21465 33983
rect 21465 33949 21499 33983
rect 21499 33949 21508 33983
rect 21456 33940 21508 33949
rect 25596 34008 25648 34060
rect 22284 33940 22336 33992
rect 22744 33940 22796 33992
rect 23572 33983 23624 33992
rect 23572 33949 23581 33983
rect 23581 33949 23615 33983
rect 23615 33949 23624 33983
rect 23572 33940 23624 33949
rect 24400 33940 24452 33992
rect 24768 33940 24820 33992
rect 25044 33983 25096 33992
rect 25044 33949 25053 33983
rect 25053 33949 25087 33983
rect 25087 33949 25096 33983
rect 25044 33940 25096 33949
rect 20996 33804 21048 33856
rect 22468 33804 22520 33856
rect 22560 33804 22612 33856
rect 25964 33983 26016 33992
rect 25964 33949 25973 33983
rect 25973 33949 26007 33983
rect 26007 33949 26016 33983
rect 25964 33940 26016 33949
rect 27528 34008 27580 34060
rect 26884 33983 26936 33992
rect 26884 33949 26893 33983
rect 26893 33949 26927 33983
rect 26927 33949 26936 33983
rect 26884 33940 26936 33949
rect 26976 33940 27028 33992
rect 27620 33940 27672 33992
rect 29276 34008 29328 34060
rect 30012 34008 30064 34060
rect 30196 34008 30248 34060
rect 28264 33940 28316 33992
rect 28816 33940 28868 33992
rect 29000 33983 29052 33992
rect 29000 33949 29009 33983
rect 29009 33949 29043 33983
rect 29043 33949 29052 33983
rect 29000 33940 29052 33949
rect 45560 34076 45612 34128
rect 44180 34008 44232 34060
rect 47124 34051 47176 34060
rect 47124 34017 47133 34051
rect 47133 34017 47167 34051
rect 47167 34017 47176 34051
rect 47124 34008 47176 34017
rect 24676 33804 24728 33856
rect 27068 33804 27120 33856
rect 27252 33804 27304 33856
rect 47216 33915 47268 33924
rect 47216 33881 47225 33915
rect 47225 33881 47259 33915
rect 47259 33881 47268 33915
rect 47216 33872 47268 33881
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 14464 33600 14516 33652
rect 16396 33600 16448 33652
rect 18144 33600 18196 33652
rect 16948 33532 17000 33584
rect 17408 33532 17460 33584
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 2504 33396 2556 33448
rect 17776 33507 17828 33516
rect 17776 33473 17785 33507
rect 17785 33473 17819 33507
rect 17819 33473 17828 33507
rect 17776 33464 17828 33473
rect 19432 33600 19484 33652
rect 20720 33600 20772 33652
rect 21272 33600 21324 33652
rect 22468 33600 22520 33652
rect 18696 33532 18748 33584
rect 19340 33532 19392 33584
rect 19708 33464 19760 33516
rect 19984 33464 20036 33516
rect 20536 33464 20588 33516
rect 24952 33532 25004 33584
rect 25320 33532 25372 33584
rect 25964 33600 26016 33652
rect 27620 33600 27672 33652
rect 27804 33600 27856 33652
rect 30012 33600 30064 33652
rect 18880 33396 18932 33448
rect 23388 33396 23440 33448
rect 23572 33464 23624 33516
rect 25596 33464 25648 33516
rect 27068 33507 27120 33516
rect 27068 33473 27077 33507
rect 27077 33473 27111 33507
rect 27111 33473 27120 33507
rect 29276 33532 29328 33584
rect 29368 33575 29420 33584
rect 29368 33541 29377 33575
rect 29377 33541 29411 33575
rect 29411 33541 29420 33575
rect 29368 33532 29420 33541
rect 27068 33464 27120 33473
rect 28816 33464 28868 33516
rect 25412 33396 25464 33448
rect 26884 33396 26936 33448
rect 27252 33439 27304 33448
rect 27252 33405 27261 33439
rect 27261 33405 27295 33439
rect 27295 33405 27304 33439
rect 27252 33396 27304 33405
rect 21088 33328 21140 33380
rect 24400 33328 24452 33380
rect 26976 33328 27028 33380
rect 30288 33464 30340 33516
rect 47860 33507 47912 33516
rect 47860 33473 47869 33507
rect 47869 33473 47903 33507
rect 47903 33473 47912 33507
rect 47860 33464 47912 33473
rect 21824 33260 21876 33312
rect 22560 33260 22612 33312
rect 24952 33260 25004 33312
rect 29000 33260 29052 33312
rect 29644 33260 29696 33312
rect 41420 33260 41472 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 16948 33099 17000 33108
rect 16948 33065 16957 33099
rect 16957 33065 16991 33099
rect 16991 33065 17000 33099
rect 16948 33056 17000 33065
rect 18696 33056 18748 33108
rect 19248 33056 19300 33108
rect 1492 32988 1544 33040
rect 1584 32963 1636 32972
rect 1584 32929 1593 32963
rect 1593 32929 1627 32963
rect 1627 32929 1636 32963
rect 1584 32920 1636 32929
rect 22284 32988 22336 33040
rect 22468 33056 22520 33108
rect 26148 33056 26200 33108
rect 27896 33099 27948 33108
rect 27896 33065 27905 33099
rect 27905 33065 27939 33099
rect 27939 33065 27948 33099
rect 27896 33056 27948 33065
rect 23848 32988 23900 33040
rect 24768 32988 24820 33040
rect 16396 32895 16448 32904
rect 16396 32861 16405 32895
rect 16405 32861 16439 32895
rect 16439 32861 16448 32895
rect 16396 32852 16448 32861
rect 16672 32895 16724 32904
rect 16672 32861 16681 32895
rect 16681 32861 16715 32895
rect 16715 32861 16724 32895
rect 16672 32852 16724 32861
rect 17684 32852 17736 32904
rect 17776 32852 17828 32904
rect 18144 32895 18196 32904
rect 18144 32861 18153 32895
rect 18153 32861 18187 32895
rect 18187 32861 18196 32895
rect 18144 32852 18196 32861
rect 3976 32784 4028 32836
rect 16948 32784 17000 32836
rect 18052 32784 18104 32836
rect 19708 32827 19760 32836
rect 19708 32793 19717 32827
rect 19717 32793 19751 32827
rect 19751 32793 19760 32827
rect 19708 32784 19760 32793
rect 20168 32784 20220 32836
rect 19340 32716 19392 32768
rect 21364 32784 21416 32836
rect 21732 32920 21784 32972
rect 24308 32920 24360 32972
rect 26792 32920 26844 32972
rect 27896 32920 27948 32972
rect 21824 32852 21876 32904
rect 22560 32852 22612 32904
rect 23940 32852 23992 32904
rect 26608 32852 26660 32904
rect 26884 32895 26936 32904
rect 26884 32861 26893 32895
rect 26893 32861 26927 32895
rect 26927 32861 26936 32895
rect 26884 32852 26936 32861
rect 27068 32852 27120 32904
rect 27252 32895 27304 32904
rect 27252 32861 27261 32895
rect 27261 32861 27295 32895
rect 27295 32861 27304 32895
rect 27252 32852 27304 32861
rect 29644 32852 29696 32904
rect 30012 32852 30064 32904
rect 46296 32895 46348 32904
rect 46296 32861 46305 32895
rect 46305 32861 46339 32895
rect 46339 32861 46348 32895
rect 46296 32852 46348 32861
rect 20444 32716 20496 32768
rect 22192 32716 22244 32768
rect 22744 32759 22796 32768
rect 22744 32725 22753 32759
rect 22753 32725 22787 32759
rect 22787 32725 22796 32759
rect 22744 32716 22796 32725
rect 25136 32784 25188 32836
rect 27344 32784 27396 32836
rect 30564 32784 30616 32836
rect 31392 32784 31444 32836
rect 47676 32784 47728 32836
rect 48136 32827 48188 32836
rect 48136 32793 48145 32827
rect 48145 32793 48179 32827
rect 48179 32793 48188 32827
rect 48136 32784 48188 32793
rect 23756 32759 23808 32768
rect 23756 32725 23765 32759
rect 23765 32725 23799 32759
rect 23799 32725 23808 32759
rect 23756 32716 23808 32725
rect 24584 32716 24636 32768
rect 24768 32716 24820 32768
rect 28172 32716 28224 32768
rect 30012 32716 30064 32768
rect 30288 32716 30340 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 20168 32512 20220 32564
rect 2504 32487 2556 32496
rect 2504 32453 2513 32487
rect 2513 32453 2547 32487
rect 2547 32453 2556 32487
rect 2504 32444 2556 32453
rect 17040 32444 17092 32496
rect 15292 32376 15344 32428
rect 17132 32419 17184 32428
rect 17132 32385 17141 32419
rect 17141 32385 17175 32419
rect 17175 32385 17184 32419
rect 17132 32376 17184 32385
rect 19984 32444 20036 32496
rect 22560 32512 22612 32564
rect 24308 32555 24360 32564
rect 24308 32521 24317 32555
rect 24317 32521 24351 32555
rect 24351 32521 24360 32555
rect 24308 32512 24360 32521
rect 28356 32512 28408 32564
rect 30564 32555 30616 32564
rect 30564 32521 30573 32555
rect 30573 32521 30607 32555
rect 30607 32521 30616 32555
rect 30564 32512 30616 32521
rect 31392 32555 31444 32564
rect 31392 32521 31401 32555
rect 31401 32521 31435 32555
rect 31435 32521 31444 32555
rect 31392 32512 31444 32521
rect 47676 32555 47728 32564
rect 47676 32521 47685 32555
rect 47685 32521 47719 32555
rect 47719 32521 47728 32555
rect 47676 32512 47728 32521
rect 23204 32487 23256 32496
rect 23204 32453 23213 32487
rect 23213 32453 23247 32487
rect 23247 32453 23256 32487
rect 23204 32444 23256 32453
rect 26424 32487 26476 32496
rect 26424 32453 26433 32487
rect 26433 32453 26467 32487
rect 26467 32453 26476 32487
rect 26424 32444 26476 32453
rect 30288 32487 30340 32496
rect 30288 32453 30297 32487
rect 30297 32453 30331 32487
rect 30331 32453 30340 32487
rect 30288 32444 30340 32453
rect 17868 32376 17920 32428
rect 18236 32376 18288 32428
rect 20444 32419 20496 32428
rect 20444 32385 20453 32419
rect 20453 32385 20487 32419
rect 20487 32385 20496 32419
rect 20444 32376 20496 32385
rect 20536 32419 20588 32428
rect 20536 32385 20545 32419
rect 20545 32385 20579 32419
rect 20579 32385 20588 32419
rect 20536 32376 20588 32385
rect 21180 32376 21232 32428
rect 2320 32351 2372 32360
rect 2320 32317 2329 32351
rect 2329 32317 2363 32351
rect 2363 32317 2372 32351
rect 2320 32308 2372 32317
rect 3976 32351 4028 32360
rect 3976 32317 3985 32351
rect 3985 32317 4019 32351
rect 4019 32317 4028 32351
rect 3976 32308 4028 32317
rect 20628 32351 20680 32360
rect 20628 32317 20637 32351
rect 20637 32317 20671 32351
rect 20671 32317 20680 32351
rect 20628 32308 20680 32317
rect 20720 32351 20772 32360
rect 20720 32317 20729 32351
rect 20729 32317 20763 32351
rect 20763 32317 20772 32351
rect 20720 32308 20772 32317
rect 17960 32240 18012 32292
rect 18052 32240 18104 32292
rect 21732 32308 21784 32360
rect 22376 32376 22428 32428
rect 23388 32376 23440 32428
rect 24216 32419 24268 32428
rect 24216 32385 24225 32419
rect 24225 32385 24259 32419
rect 24259 32385 24268 32419
rect 24216 32376 24268 32385
rect 24952 32419 25004 32428
rect 24952 32385 24961 32419
rect 24961 32385 24995 32419
rect 24995 32385 25004 32419
rect 24952 32376 25004 32385
rect 27988 32376 28040 32428
rect 29920 32419 29972 32428
rect 29920 32385 29929 32419
rect 29929 32385 29963 32419
rect 29963 32385 29972 32419
rect 29920 32376 29972 32385
rect 30012 32419 30064 32428
rect 30012 32385 30022 32419
rect 30022 32385 30056 32419
rect 30056 32385 30064 32419
rect 30196 32419 30248 32428
rect 30012 32376 30064 32385
rect 30196 32385 30205 32419
rect 30205 32385 30239 32419
rect 30239 32385 30248 32419
rect 30196 32376 30248 32385
rect 25320 32308 25372 32360
rect 26424 32308 26476 32360
rect 28264 32308 28316 32360
rect 29736 32308 29788 32360
rect 31300 32419 31352 32428
rect 31300 32385 31309 32419
rect 31309 32385 31343 32419
rect 31343 32385 31352 32419
rect 31300 32376 31352 32385
rect 21456 32240 21508 32292
rect 1400 32172 1452 32224
rect 15660 32172 15712 32224
rect 17224 32215 17276 32224
rect 17224 32181 17233 32215
rect 17233 32181 17267 32215
rect 17267 32181 17276 32215
rect 17224 32172 17276 32181
rect 18512 32172 18564 32224
rect 21824 32172 21876 32224
rect 23204 32240 23256 32292
rect 46296 32376 46348 32428
rect 47492 32376 47544 32428
rect 47676 32376 47728 32428
rect 41420 32240 41472 32292
rect 22744 32172 22796 32224
rect 23572 32215 23624 32224
rect 23572 32181 23581 32215
rect 23581 32181 23615 32215
rect 23615 32181 23624 32215
rect 23572 32172 23624 32181
rect 25228 32172 25280 32224
rect 25688 32172 25740 32224
rect 28172 32215 28224 32224
rect 28172 32181 28181 32215
rect 28181 32181 28215 32215
rect 28215 32181 28224 32215
rect 28172 32172 28224 32181
rect 29644 32172 29696 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 17132 31968 17184 32020
rect 18328 31968 18380 32020
rect 21364 32011 21416 32020
rect 21364 31977 21373 32011
rect 21373 31977 21407 32011
rect 21407 31977 21416 32011
rect 21364 31968 21416 31977
rect 21732 31968 21784 32020
rect 23388 31968 23440 32020
rect 27528 31968 27580 32020
rect 29276 31968 29328 32020
rect 29920 31968 29972 32020
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 1860 31875 1912 31884
rect 1860 31841 1869 31875
rect 1869 31841 1903 31875
rect 1903 31841 1912 31875
rect 1860 31832 1912 31841
rect 14188 31832 14240 31884
rect 16764 31875 16816 31884
rect 16764 31841 16773 31875
rect 16773 31841 16807 31875
rect 16807 31841 16816 31875
rect 16764 31832 16816 31841
rect 15660 31764 15712 31816
rect 17224 31832 17276 31884
rect 17960 31832 18012 31884
rect 1584 31739 1636 31748
rect 1584 31705 1593 31739
rect 1593 31705 1627 31739
rect 1627 31705 1636 31739
rect 1584 31696 1636 31705
rect 18512 31807 18564 31816
rect 18512 31773 18521 31807
rect 18521 31773 18555 31807
rect 18555 31773 18564 31807
rect 18512 31764 18564 31773
rect 25596 31900 25648 31952
rect 28172 31900 28224 31952
rect 28356 31900 28408 31952
rect 29736 31900 29788 31952
rect 30196 31900 30248 31952
rect 21824 31875 21876 31884
rect 19432 31764 19484 31816
rect 21824 31841 21833 31875
rect 21833 31841 21867 31875
rect 21867 31841 21876 31875
rect 21824 31832 21876 31841
rect 24768 31832 24820 31884
rect 22192 31807 22244 31816
rect 22192 31773 22201 31807
rect 22201 31773 22235 31807
rect 22235 31773 22244 31807
rect 22192 31764 22244 31773
rect 18328 31696 18380 31748
rect 19248 31696 19300 31748
rect 21456 31696 21508 31748
rect 22100 31696 22152 31748
rect 23204 31764 23256 31816
rect 24032 31764 24084 31816
rect 24584 31807 24636 31816
rect 24584 31773 24593 31807
rect 24593 31773 24627 31807
rect 24627 31773 24636 31807
rect 24584 31764 24636 31773
rect 24860 31764 24912 31816
rect 26148 31764 26200 31816
rect 46020 31832 46072 31884
rect 28172 31807 28224 31816
rect 28172 31773 28181 31807
rect 28181 31773 28215 31807
rect 28215 31773 28224 31807
rect 28356 31807 28408 31816
rect 28172 31764 28224 31773
rect 28356 31773 28365 31807
rect 28365 31773 28399 31807
rect 28399 31773 28408 31807
rect 28356 31764 28408 31773
rect 28816 31764 28868 31816
rect 29644 31807 29696 31816
rect 29644 31773 29653 31807
rect 29653 31773 29687 31807
rect 29687 31773 29696 31807
rect 29644 31764 29696 31773
rect 29828 31807 29880 31816
rect 29828 31773 29837 31807
rect 29837 31773 29871 31807
rect 29871 31773 29880 31807
rect 29828 31764 29880 31773
rect 44180 31764 44232 31816
rect 47308 31807 47360 31816
rect 47308 31773 47317 31807
rect 47317 31773 47351 31807
rect 47351 31773 47360 31807
rect 47308 31764 47360 31773
rect 27988 31696 28040 31748
rect 17408 31628 17460 31680
rect 17868 31628 17920 31680
rect 18236 31628 18288 31680
rect 21180 31628 21232 31680
rect 23480 31628 23532 31680
rect 24216 31628 24268 31680
rect 26424 31671 26476 31680
rect 26424 31637 26433 31671
rect 26433 31637 26467 31671
rect 26467 31637 26476 31671
rect 26424 31628 26476 31637
rect 27712 31628 27764 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1584 31424 1636 31476
rect 15476 31424 15528 31476
rect 15660 31356 15712 31408
rect 2136 31331 2188 31340
rect 2136 31297 2145 31331
rect 2145 31297 2179 31331
rect 2179 31297 2188 31331
rect 2136 31288 2188 31297
rect 2412 31288 2464 31340
rect 16764 31288 16816 31340
rect 17132 31288 17184 31340
rect 18880 31356 18932 31408
rect 22008 31356 22060 31408
rect 24584 31424 24636 31476
rect 24768 31424 24820 31476
rect 30196 31424 30248 31476
rect 22744 31356 22796 31408
rect 27988 31356 28040 31408
rect 18512 31288 18564 31340
rect 20628 31331 20680 31340
rect 18052 31263 18104 31272
rect 18052 31229 18061 31263
rect 18061 31229 18095 31263
rect 18095 31229 18104 31263
rect 18052 31220 18104 31229
rect 17960 31152 18012 31204
rect 18328 31220 18380 31272
rect 19340 31220 19392 31272
rect 20628 31297 20637 31331
rect 20637 31297 20671 31331
rect 20671 31297 20680 31331
rect 20628 31288 20680 31297
rect 20720 31331 20772 31340
rect 20720 31297 20730 31331
rect 20730 31297 20764 31331
rect 20764 31297 20772 31331
rect 20996 31331 21048 31340
rect 20720 31288 20772 31297
rect 20996 31297 21005 31331
rect 21005 31297 21039 31331
rect 21039 31297 21048 31331
rect 20996 31288 21048 31297
rect 20352 31220 20404 31272
rect 24768 31288 24820 31340
rect 27712 31288 27764 31340
rect 28080 31331 28132 31340
rect 28080 31297 28089 31331
rect 28089 31297 28123 31331
rect 28123 31297 28132 31331
rect 28080 31288 28132 31297
rect 28908 31288 28960 31340
rect 29276 31356 29328 31408
rect 21732 31152 21784 31204
rect 16028 31084 16080 31136
rect 16764 31084 16816 31136
rect 18052 31084 18104 31136
rect 20904 31084 20956 31136
rect 25320 31220 25372 31272
rect 25780 31263 25832 31272
rect 25780 31229 25789 31263
rect 25789 31229 25823 31263
rect 25823 31229 25832 31263
rect 25780 31220 25832 31229
rect 28172 31220 28224 31272
rect 27068 31152 27120 31204
rect 28816 31195 28868 31204
rect 28816 31161 28825 31195
rect 28825 31161 28859 31195
rect 28859 31161 28868 31195
rect 28816 31152 28868 31161
rect 30104 31220 30156 31272
rect 23572 31127 23624 31136
rect 23572 31093 23581 31127
rect 23581 31093 23615 31127
rect 23615 31093 23624 31127
rect 23572 31084 23624 31093
rect 26700 31084 26752 31136
rect 27620 31084 27672 31136
rect 28632 31084 28684 31136
rect 30104 31084 30156 31136
rect 31024 31084 31076 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 15660 30880 15712 30932
rect 17132 30880 17184 30932
rect 20996 30880 21048 30932
rect 22744 30923 22796 30932
rect 20628 30812 20680 30864
rect 21916 30812 21968 30864
rect 22744 30889 22753 30923
rect 22753 30889 22787 30923
rect 22787 30889 22796 30923
rect 22744 30880 22796 30889
rect 27068 30880 27120 30932
rect 28172 30923 28224 30932
rect 23112 30812 23164 30864
rect 14556 30744 14608 30796
rect 15476 30719 15528 30728
rect 15476 30685 15485 30719
rect 15485 30685 15519 30719
rect 15519 30685 15528 30719
rect 15476 30676 15528 30685
rect 16856 30719 16908 30728
rect 16856 30685 16865 30719
rect 16865 30685 16899 30719
rect 16899 30685 16908 30719
rect 16856 30676 16908 30685
rect 16948 30676 17000 30728
rect 22100 30744 22152 30796
rect 17960 30676 18012 30728
rect 18236 30719 18288 30728
rect 18236 30685 18245 30719
rect 18245 30685 18279 30719
rect 18279 30685 18288 30719
rect 18236 30676 18288 30685
rect 21180 30676 21232 30728
rect 21916 30676 21968 30728
rect 22376 30676 22428 30728
rect 24860 30744 24912 30796
rect 27896 30744 27948 30796
rect 28172 30889 28181 30923
rect 28181 30889 28215 30923
rect 28215 30889 28224 30923
rect 28172 30880 28224 30889
rect 28816 30923 28868 30932
rect 28816 30889 28825 30923
rect 28825 30889 28859 30923
rect 28859 30889 28868 30923
rect 28816 30880 28868 30889
rect 28080 30812 28132 30864
rect 25136 30676 25188 30728
rect 28632 30719 28684 30728
rect 28632 30685 28641 30719
rect 28641 30685 28675 30719
rect 28675 30685 28684 30719
rect 28632 30676 28684 30685
rect 16672 30608 16724 30660
rect 20720 30608 20772 30660
rect 22008 30651 22060 30660
rect 22008 30617 22017 30651
rect 22017 30617 22051 30651
rect 22051 30617 22060 30651
rect 22008 30608 22060 30617
rect 23572 30608 23624 30660
rect 26700 30651 26752 30660
rect 26700 30617 26709 30651
rect 26709 30617 26743 30651
rect 26743 30617 26752 30651
rect 26700 30608 26752 30617
rect 27712 30608 27764 30660
rect 28172 30608 28224 30660
rect 30472 30651 30524 30660
rect 30472 30617 30481 30651
rect 30481 30617 30515 30651
rect 30515 30617 30524 30651
rect 30472 30608 30524 30617
rect 31116 30608 31168 30660
rect 17316 30540 17368 30592
rect 21272 30540 21324 30592
rect 28356 30540 28408 30592
rect 28908 30540 28960 30592
rect 30104 30540 30156 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 19984 30268 20036 30320
rect 20536 30311 20588 30320
rect 20536 30277 20545 30311
rect 20545 30277 20579 30311
rect 20579 30277 20588 30311
rect 20536 30268 20588 30277
rect 20720 30268 20772 30320
rect 21916 30268 21968 30320
rect 23848 30268 23900 30320
rect 20352 30243 20404 30252
rect 20352 30209 20361 30243
rect 20361 30209 20395 30243
rect 20395 30209 20404 30243
rect 20352 30200 20404 30209
rect 25596 30268 25648 30320
rect 26148 30336 26200 30388
rect 25780 30268 25832 30320
rect 27344 30268 27396 30320
rect 12992 30175 13044 30184
rect 12992 30141 13001 30175
rect 13001 30141 13035 30175
rect 13035 30141 13044 30175
rect 12992 30132 13044 30141
rect 13452 30132 13504 30184
rect 8300 30064 8352 30116
rect 18236 30132 18288 30184
rect 21272 30132 21324 30184
rect 21364 30132 21416 30184
rect 24584 30200 24636 30252
rect 18972 30064 19024 30116
rect 19432 29996 19484 30048
rect 20444 29996 20496 30048
rect 21548 30064 21600 30116
rect 22560 30064 22612 30116
rect 25504 30200 25556 30252
rect 28632 30336 28684 30388
rect 30472 30336 30524 30388
rect 28172 30268 28224 30320
rect 30380 30268 30432 30320
rect 28540 30200 28592 30252
rect 28816 30200 28868 30252
rect 30104 30200 30156 30252
rect 30288 30200 30340 30252
rect 31024 30243 31076 30252
rect 31024 30209 31033 30243
rect 31033 30209 31067 30243
rect 31067 30209 31076 30243
rect 31024 30200 31076 30209
rect 26056 30132 26108 30184
rect 23848 30039 23900 30048
rect 23848 30005 23857 30039
rect 23857 30005 23891 30039
rect 23891 30005 23900 30039
rect 23848 29996 23900 30005
rect 25136 29996 25188 30048
rect 26148 30064 26200 30116
rect 28632 30064 28684 30116
rect 25872 30039 25924 30048
rect 25872 30005 25881 30039
rect 25881 30005 25915 30039
rect 25915 30005 25924 30039
rect 25872 29996 25924 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 21916 29835 21968 29844
rect 21916 29801 21925 29835
rect 21925 29801 21959 29835
rect 21959 29801 21968 29835
rect 21916 29792 21968 29801
rect 25504 29835 25556 29844
rect 25504 29801 25513 29835
rect 25513 29801 25547 29835
rect 25547 29801 25556 29835
rect 25504 29792 25556 29801
rect 26148 29835 26200 29844
rect 26148 29801 26157 29835
rect 26157 29801 26191 29835
rect 26191 29801 26200 29835
rect 26148 29792 26200 29801
rect 27068 29835 27120 29844
rect 27068 29801 27077 29835
rect 27077 29801 27111 29835
rect 27111 29801 27120 29835
rect 27068 29792 27120 29801
rect 27712 29835 27764 29844
rect 27712 29801 27721 29835
rect 27721 29801 27755 29835
rect 27755 29801 27764 29835
rect 27712 29792 27764 29801
rect 31116 29835 31168 29844
rect 31116 29801 31125 29835
rect 31125 29801 31159 29835
rect 31159 29801 31168 29835
rect 31116 29792 31168 29801
rect 24216 29724 24268 29776
rect 24952 29724 25004 29776
rect 13820 29588 13872 29640
rect 17316 29631 17368 29640
rect 17316 29597 17325 29631
rect 17325 29597 17359 29631
rect 17359 29597 17368 29631
rect 17316 29588 17368 29597
rect 17592 29631 17644 29640
rect 17592 29597 17601 29631
rect 17601 29597 17635 29631
rect 17635 29597 17644 29631
rect 17592 29588 17644 29597
rect 18236 29588 18288 29640
rect 20260 29588 20312 29640
rect 20444 29588 20496 29640
rect 20720 29588 20772 29640
rect 22008 29631 22060 29640
rect 14280 29495 14332 29504
rect 14280 29461 14289 29495
rect 14289 29461 14323 29495
rect 14323 29461 14332 29495
rect 14280 29452 14332 29461
rect 14924 29495 14976 29504
rect 14924 29461 14933 29495
rect 14933 29461 14967 29495
rect 14967 29461 14976 29495
rect 14924 29452 14976 29461
rect 16672 29452 16724 29504
rect 18604 29452 18656 29504
rect 18880 29452 18932 29504
rect 21180 29520 21232 29572
rect 22008 29597 22017 29631
rect 22017 29597 22051 29631
rect 22051 29597 22060 29631
rect 22008 29588 22060 29597
rect 22376 29588 22428 29640
rect 23664 29588 23716 29640
rect 22100 29520 22152 29572
rect 25872 29588 25924 29640
rect 26056 29631 26108 29640
rect 26056 29597 26065 29631
rect 26065 29597 26099 29631
rect 26099 29597 26108 29631
rect 26056 29588 26108 29597
rect 26148 29631 26200 29640
rect 26148 29597 26157 29631
rect 26157 29597 26191 29631
rect 26191 29597 26200 29631
rect 26148 29588 26200 29597
rect 27344 29588 27396 29640
rect 28356 29588 28408 29640
rect 28632 29631 28684 29640
rect 28632 29597 28641 29631
rect 28641 29597 28675 29631
rect 28675 29597 28684 29631
rect 28632 29588 28684 29597
rect 29000 29588 29052 29640
rect 30288 29588 30340 29640
rect 30840 29588 30892 29640
rect 47308 29631 47360 29640
rect 47308 29597 47317 29631
rect 47317 29597 47351 29631
rect 47351 29597 47360 29631
rect 47308 29588 47360 29597
rect 47400 29588 47452 29640
rect 20536 29452 20588 29504
rect 21272 29452 21324 29504
rect 22560 29495 22612 29504
rect 22560 29461 22569 29495
rect 22569 29461 22603 29495
rect 22603 29461 22612 29495
rect 22560 29452 22612 29461
rect 24216 29452 24268 29504
rect 29000 29452 29052 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 13452 29291 13504 29300
rect 13452 29257 13461 29291
rect 13461 29257 13495 29291
rect 13495 29257 13504 29291
rect 13452 29248 13504 29257
rect 17592 29291 17644 29300
rect 17592 29257 17601 29291
rect 17601 29257 17635 29291
rect 17635 29257 17644 29291
rect 17592 29248 17644 29257
rect 14280 29223 14332 29232
rect 14280 29189 14289 29223
rect 14289 29189 14323 29223
rect 14323 29189 14332 29223
rect 14280 29180 14332 29189
rect 15936 29223 15988 29232
rect 15936 29189 15945 29223
rect 15945 29189 15979 29223
rect 15979 29189 15988 29223
rect 15936 29180 15988 29189
rect 13820 29112 13872 29164
rect 11704 29044 11756 29096
rect 16856 29112 16908 29164
rect 17960 29112 18012 29164
rect 19800 29180 19852 29232
rect 18236 29155 18288 29164
rect 18236 29121 18245 29155
rect 18245 29121 18279 29155
rect 18279 29121 18288 29155
rect 18236 29112 18288 29121
rect 18604 29155 18656 29164
rect 18604 29121 18613 29155
rect 18613 29121 18647 29155
rect 18647 29121 18656 29155
rect 18604 29112 18656 29121
rect 20444 29248 20496 29300
rect 20260 29180 20312 29232
rect 20536 29155 20588 29164
rect 7840 28976 7892 29028
rect 19156 29044 19208 29096
rect 20536 29121 20545 29155
rect 20545 29121 20579 29155
rect 20579 29121 20588 29155
rect 20536 29112 20588 29121
rect 21180 29112 21232 29164
rect 21364 29112 21416 29164
rect 22100 29112 22152 29164
rect 22652 29112 22704 29164
rect 25504 29112 25556 29164
rect 19340 28976 19392 29028
rect 18052 28908 18104 28960
rect 19064 28908 19116 28960
rect 23848 29044 23900 29096
rect 25688 29044 25740 29096
rect 29184 29112 29236 29164
rect 28908 29044 28960 29096
rect 29460 29087 29512 29096
rect 29460 29053 29469 29087
rect 29469 29053 29503 29087
rect 29503 29053 29512 29087
rect 29460 29044 29512 29053
rect 21732 28976 21784 29028
rect 21824 28976 21876 29028
rect 26424 28976 26476 29028
rect 27252 28976 27304 29028
rect 21180 28908 21232 28960
rect 22008 28951 22060 28960
rect 22008 28917 22017 28951
rect 22017 28917 22051 28951
rect 22051 28917 22060 28951
rect 22008 28908 22060 28917
rect 25412 28951 25464 28960
rect 25412 28917 25421 28951
rect 25421 28917 25455 28951
rect 25455 28917 25464 28951
rect 25412 28908 25464 28917
rect 29000 28976 29052 29028
rect 30380 29112 30432 29164
rect 31668 29112 31720 29164
rect 30196 28908 30248 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 11980 28704 12032 28756
rect 11612 28568 11664 28620
rect 17960 28704 18012 28756
rect 19064 28704 19116 28756
rect 19340 28747 19392 28756
rect 19340 28713 19349 28747
rect 19349 28713 19383 28747
rect 19383 28713 19392 28747
rect 19340 28704 19392 28713
rect 19800 28747 19852 28756
rect 19800 28713 19809 28747
rect 19809 28713 19843 28747
rect 19843 28713 19852 28747
rect 19800 28704 19852 28713
rect 20352 28704 20404 28756
rect 21824 28704 21876 28756
rect 22652 28747 22704 28756
rect 22652 28713 22661 28747
rect 22661 28713 22695 28747
rect 22695 28713 22704 28747
rect 22652 28704 22704 28713
rect 25412 28747 25464 28756
rect 25412 28713 25421 28747
rect 25421 28713 25455 28747
rect 25455 28713 25464 28747
rect 25412 28704 25464 28713
rect 13268 28568 13320 28620
rect 14924 28568 14976 28620
rect 16028 28568 16080 28620
rect 16672 28611 16724 28620
rect 16672 28577 16681 28611
rect 16681 28577 16715 28611
rect 16715 28577 16724 28611
rect 16672 28568 16724 28577
rect 19432 28568 19484 28620
rect 20904 28611 20956 28620
rect 20904 28577 20913 28611
rect 20913 28577 20947 28611
rect 20947 28577 20956 28611
rect 20904 28568 20956 28577
rect 21180 28611 21232 28620
rect 21180 28577 21189 28611
rect 21189 28577 21223 28611
rect 21223 28577 21232 28611
rect 21180 28568 21232 28577
rect 23480 28568 23532 28620
rect 23756 28611 23808 28620
rect 23756 28577 23765 28611
rect 23765 28577 23799 28611
rect 23799 28577 23808 28611
rect 23756 28568 23808 28577
rect 10876 28500 10928 28552
rect 12532 28432 12584 28484
rect 16580 28432 16632 28484
rect 17408 28432 17460 28484
rect 20720 28500 20772 28552
rect 24400 28543 24452 28552
rect 24400 28509 24409 28543
rect 24409 28509 24443 28543
rect 24443 28509 24452 28543
rect 24400 28500 24452 28509
rect 31668 28679 31720 28688
rect 31668 28645 31677 28679
rect 31677 28645 31711 28679
rect 31711 28645 31720 28679
rect 31668 28636 31720 28645
rect 30196 28611 30248 28620
rect 30196 28577 30205 28611
rect 30205 28577 30239 28611
rect 30239 28577 30248 28611
rect 30196 28568 30248 28577
rect 40408 28568 40460 28620
rect 47400 28568 47452 28620
rect 47860 28611 47912 28620
rect 47860 28577 47869 28611
rect 47869 28577 47903 28611
rect 47903 28577 47912 28611
rect 47860 28568 47912 28577
rect 25780 28543 25832 28552
rect 22560 28432 22612 28484
rect 23664 28432 23716 28484
rect 24216 28432 24268 28484
rect 25228 28432 25280 28484
rect 25780 28509 25789 28543
rect 25789 28509 25823 28543
rect 25823 28509 25832 28543
rect 25780 28500 25832 28509
rect 26424 28543 26476 28552
rect 26424 28509 26433 28543
rect 26433 28509 26467 28543
rect 26467 28509 26476 28543
rect 26424 28500 26476 28509
rect 26608 28543 26660 28552
rect 26608 28509 26617 28543
rect 26617 28509 26651 28543
rect 26651 28509 26660 28543
rect 26608 28500 26660 28509
rect 26700 28543 26752 28552
rect 26700 28509 26709 28543
rect 26709 28509 26743 28543
rect 26743 28509 26752 28543
rect 26700 28500 26752 28509
rect 20720 28364 20772 28416
rect 22928 28364 22980 28416
rect 24492 28364 24544 28416
rect 26240 28364 26292 28416
rect 27252 28500 27304 28552
rect 28356 28543 28408 28552
rect 28356 28509 28365 28543
rect 28365 28509 28399 28543
rect 28399 28509 28408 28543
rect 28356 28500 28408 28509
rect 29092 28500 29144 28552
rect 46296 28543 46348 28552
rect 46296 28509 46305 28543
rect 46305 28509 46339 28543
rect 46339 28509 46348 28543
rect 46296 28500 46348 28509
rect 28632 28432 28684 28484
rect 30932 28432 30984 28484
rect 27252 28364 27304 28416
rect 29184 28364 29236 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 1676 28160 1728 28212
rect 10876 28203 10928 28212
rect 10876 28169 10885 28203
rect 10885 28169 10919 28203
rect 10919 28169 10928 28203
rect 10876 28160 10928 28169
rect 11612 28203 11664 28212
rect 11612 28169 11621 28203
rect 11621 28169 11655 28203
rect 11655 28169 11664 28203
rect 11612 28160 11664 28169
rect 12532 28203 12584 28212
rect 12532 28169 12541 28203
rect 12541 28169 12575 28203
rect 12575 28169 12584 28203
rect 12532 28160 12584 28169
rect 10508 28024 10560 28076
rect 11520 28067 11572 28076
rect 11520 28033 11529 28067
rect 11529 28033 11563 28067
rect 11563 28033 11572 28067
rect 11520 28024 11572 28033
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 12348 28024 12400 28076
rect 14096 27956 14148 28008
rect 14464 27999 14516 28008
rect 14464 27965 14473 27999
rect 14473 27965 14507 27999
rect 14507 27965 14516 27999
rect 14464 27956 14516 27965
rect 16028 28024 16080 28076
rect 19248 28160 19300 28212
rect 19432 28160 19484 28212
rect 20720 28160 20772 28212
rect 21916 28160 21968 28212
rect 22652 28160 22704 28212
rect 23112 28203 23164 28212
rect 23112 28169 23121 28203
rect 23121 28169 23155 28203
rect 23155 28169 23164 28203
rect 23112 28160 23164 28169
rect 24400 28160 24452 28212
rect 26148 28160 26200 28212
rect 26700 28160 26752 28212
rect 30932 28203 30984 28212
rect 30932 28169 30941 28203
rect 30941 28169 30975 28203
rect 30975 28169 30984 28203
rect 30932 28160 30984 28169
rect 18052 28092 18104 28144
rect 18512 28092 18564 28144
rect 19064 28092 19116 28144
rect 20536 28067 20588 28076
rect 3332 27888 3384 27940
rect 14188 27888 14240 27940
rect 14372 27888 14424 27940
rect 19156 27956 19208 28008
rect 20536 28033 20545 28067
rect 20545 28033 20579 28067
rect 20579 28033 20588 28067
rect 20536 28024 20588 28033
rect 20628 28067 20680 28076
rect 20628 28033 20637 28067
rect 20637 28033 20671 28067
rect 20671 28033 20680 28067
rect 21824 28067 21876 28076
rect 20628 28024 20680 28033
rect 21824 28033 21833 28067
rect 21833 28033 21867 28067
rect 21867 28033 21876 28067
rect 21824 28024 21876 28033
rect 22928 28067 22980 28076
rect 22928 28033 22937 28067
rect 22937 28033 22971 28067
rect 22971 28033 22980 28067
rect 22928 28024 22980 28033
rect 25228 28024 25280 28076
rect 25412 28067 25464 28076
rect 25412 28033 25421 28067
rect 25421 28033 25455 28067
rect 25455 28033 25464 28067
rect 25412 28024 25464 28033
rect 27252 28135 27304 28144
rect 27252 28101 27261 28135
rect 27261 28101 27295 28135
rect 27295 28101 27304 28135
rect 27252 28092 27304 28101
rect 27988 28092 28040 28144
rect 26976 28067 27028 28076
rect 26976 28033 26985 28067
rect 26985 28033 27019 28067
rect 27019 28033 27028 28067
rect 26976 28024 27028 28033
rect 29184 28067 29236 28076
rect 29184 28033 29193 28067
rect 29193 28033 29227 28067
rect 29227 28033 29236 28067
rect 29184 28024 29236 28033
rect 30840 28067 30892 28076
rect 30840 28033 30849 28067
rect 30849 28033 30883 28067
rect 30883 28033 30892 28067
rect 30840 28024 30892 28033
rect 25596 27999 25648 28008
rect 25596 27965 25605 27999
rect 25605 27965 25639 27999
rect 25639 27965 25648 27999
rect 25596 27956 25648 27965
rect 25872 27956 25924 28008
rect 47860 28160 47912 28212
rect 47216 28024 47268 28076
rect 25780 27888 25832 27940
rect 28908 27888 28960 27940
rect 20352 27820 20404 27872
rect 21180 27820 21232 27872
rect 21548 27820 21600 27872
rect 22744 27863 22796 27872
rect 22744 27829 22753 27863
rect 22753 27829 22787 27863
rect 22787 27829 22796 27863
rect 22744 27820 22796 27829
rect 25228 27820 25280 27872
rect 29000 27820 29052 27872
rect 29552 27863 29604 27872
rect 29552 27829 29561 27863
rect 29561 27829 29595 27863
rect 29595 27829 29604 27863
rect 29552 27820 29604 27829
rect 47032 27863 47084 27872
rect 47032 27829 47041 27863
rect 47041 27829 47075 27863
rect 47075 27829 47084 27863
rect 47032 27820 47084 27829
rect 47676 27863 47728 27872
rect 47676 27829 47685 27863
rect 47685 27829 47719 27863
rect 47719 27829 47728 27863
rect 47676 27820 47728 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 14464 27616 14516 27668
rect 20352 27616 20404 27668
rect 22744 27616 22796 27668
rect 26516 27616 26568 27668
rect 26976 27616 27028 27668
rect 29092 27616 29144 27668
rect 32220 27616 32272 27668
rect 45560 27616 45612 27668
rect 17408 27548 17460 27600
rect 18512 27591 18564 27600
rect 18512 27557 18521 27591
rect 18521 27557 18555 27591
rect 18555 27557 18564 27591
rect 18512 27548 18564 27557
rect 21824 27548 21876 27600
rect 23388 27548 23440 27600
rect 13820 27480 13872 27532
rect 20536 27480 20588 27532
rect 20904 27480 20956 27532
rect 23756 27480 23808 27532
rect 11152 27455 11204 27464
rect 11152 27421 11161 27455
rect 11161 27421 11195 27455
rect 11195 27421 11204 27455
rect 11152 27412 11204 27421
rect 12348 27412 12400 27464
rect 13912 27412 13964 27464
rect 14740 27455 14792 27464
rect 14740 27421 14749 27455
rect 14749 27421 14783 27455
rect 14783 27421 14792 27455
rect 14740 27412 14792 27421
rect 19064 27412 19116 27464
rect 21088 27412 21140 27464
rect 25412 27480 25464 27532
rect 25780 27412 25832 27464
rect 25872 27455 25924 27464
rect 25872 27421 25881 27455
rect 25881 27421 25915 27455
rect 25915 27421 25924 27455
rect 25872 27412 25924 27421
rect 12440 27344 12492 27396
rect 20720 27344 20772 27396
rect 23664 27344 23716 27396
rect 26516 27480 26568 27532
rect 26700 27455 26752 27464
rect 26700 27421 26709 27455
rect 26709 27421 26743 27455
rect 26743 27421 26752 27455
rect 26700 27412 26752 27421
rect 28448 27548 28500 27600
rect 28540 27548 28592 27600
rect 28816 27548 28868 27600
rect 29276 27548 29328 27600
rect 28172 27412 28224 27464
rect 28954 27480 29006 27532
rect 29552 27480 29604 27532
rect 47032 27480 47084 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 28540 27455 28592 27464
rect 28540 27421 28549 27455
rect 28549 27421 28583 27455
rect 28583 27421 28592 27455
rect 28540 27412 28592 27421
rect 30840 27412 30892 27464
rect 10784 27276 10836 27328
rect 12072 27319 12124 27328
rect 12072 27285 12081 27319
rect 12081 27285 12115 27319
rect 12115 27285 12124 27319
rect 12072 27276 12124 27285
rect 14188 27319 14240 27328
rect 14188 27285 14197 27319
rect 14197 27285 14231 27319
rect 14231 27285 14240 27319
rect 14188 27276 14240 27285
rect 25596 27276 25648 27328
rect 25688 27276 25740 27328
rect 27896 27276 27948 27328
rect 28448 27276 28500 27328
rect 47676 27344 47728 27396
rect 28908 27276 28960 27328
rect 29368 27276 29420 27328
rect 30380 27276 30432 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 11520 27072 11572 27124
rect 11428 27004 11480 27056
rect 11704 27004 11756 27056
rect 12440 27072 12492 27124
rect 13084 27072 13136 27124
rect 13176 27072 13228 27124
rect 27988 27115 28040 27124
rect 13452 27004 13504 27056
rect 14188 27004 14240 27056
rect 10508 26979 10560 26988
rect 10508 26945 10517 26979
rect 10517 26945 10551 26979
rect 10551 26945 10560 26979
rect 10508 26936 10560 26945
rect 11980 26936 12032 26988
rect 21824 27004 21876 27056
rect 27988 27081 27997 27115
rect 27997 27081 28031 27115
rect 28031 27081 28040 27115
rect 27988 27072 28040 27081
rect 28540 27072 28592 27124
rect 45836 27072 45888 27124
rect 46204 27072 46256 27124
rect 24032 27004 24084 27056
rect 15844 26936 15896 26988
rect 20260 26979 20312 26988
rect 20260 26945 20269 26979
rect 20269 26945 20303 26979
rect 20303 26945 20312 26979
rect 20260 26936 20312 26945
rect 20536 26936 20588 26988
rect 21088 26936 21140 26988
rect 25688 26979 25740 26988
rect 25688 26945 25697 26979
rect 25697 26945 25731 26979
rect 25731 26945 25740 26979
rect 25688 26936 25740 26945
rect 26608 27004 26660 27056
rect 26240 26979 26292 26988
rect 26240 26945 26249 26979
rect 26249 26945 26283 26979
rect 26283 26945 26292 26979
rect 28448 27004 28500 27056
rect 29368 27047 29420 27056
rect 29368 27013 29377 27047
rect 29377 27013 29411 27047
rect 29411 27013 29420 27047
rect 29368 27004 29420 27013
rect 30380 27004 30432 27056
rect 26240 26936 26292 26945
rect 27896 26979 27948 26988
rect 27896 26945 27905 26979
rect 27905 26945 27939 26979
rect 27939 26945 27948 26979
rect 27896 26936 27948 26945
rect 28816 26936 28868 26988
rect 29092 26979 29144 26988
rect 29092 26945 29101 26979
rect 29101 26945 29135 26979
rect 29135 26945 29144 26979
rect 29092 26936 29144 26945
rect 45836 26936 45888 26988
rect 13176 26911 13228 26920
rect 11888 26800 11940 26852
rect 12256 26800 12308 26852
rect 10508 26775 10560 26784
rect 10508 26741 10517 26775
rect 10517 26741 10551 26775
rect 10551 26741 10560 26775
rect 10508 26732 10560 26741
rect 13176 26877 13185 26911
rect 13185 26877 13219 26911
rect 13219 26877 13228 26911
rect 13176 26868 13228 26877
rect 20812 26868 20864 26920
rect 25596 26868 25648 26920
rect 20720 26800 20772 26852
rect 21272 26800 21324 26852
rect 26056 26911 26108 26920
rect 26056 26877 26065 26911
rect 26065 26877 26099 26911
rect 26099 26877 26108 26911
rect 26056 26868 26108 26877
rect 32128 26868 32180 26920
rect 47492 26868 47544 26920
rect 26700 26800 26752 26852
rect 13820 26732 13872 26784
rect 16120 26775 16172 26784
rect 16120 26741 16129 26775
rect 16129 26741 16163 26775
rect 16163 26741 16172 26775
rect 16120 26732 16172 26741
rect 18236 26732 18288 26784
rect 20444 26732 20496 26784
rect 26424 26775 26476 26784
rect 26424 26741 26433 26775
rect 26433 26741 26467 26775
rect 26467 26741 26476 26775
rect 26424 26732 26476 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 12256 26571 12308 26580
rect 12256 26537 12265 26571
rect 12265 26537 12299 26571
rect 12299 26537 12308 26571
rect 12256 26528 12308 26537
rect 23664 26571 23716 26580
rect 10508 26435 10560 26444
rect 10508 26401 10517 26435
rect 10517 26401 10551 26435
rect 10551 26401 10560 26435
rect 10508 26392 10560 26401
rect 10784 26435 10836 26444
rect 10784 26401 10793 26435
rect 10793 26401 10827 26435
rect 10827 26401 10836 26435
rect 10784 26392 10836 26401
rect 13452 26392 13504 26444
rect 12072 26256 12124 26308
rect 12256 26256 12308 26308
rect 13268 26367 13320 26376
rect 13268 26333 13277 26367
rect 13277 26333 13311 26367
rect 13311 26333 13320 26367
rect 16120 26460 16172 26512
rect 13268 26324 13320 26333
rect 15752 26367 15804 26376
rect 12992 26299 13044 26308
rect 12992 26265 13001 26299
rect 13001 26265 13035 26299
rect 13035 26265 13044 26299
rect 12992 26256 13044 26265
rect 13452 26256 13504 26308
rect 11428 26188 11480 26240
rect 15752 26333 15761 26367
rect 15761 26333 15795 26367
rect 15795 26333 15804 26367
rect 15752 26324 15804 26333
rect 20812 26324 20864 26376
rect 21456 26324 21508 26376
rect 21916 26460 21968 26512
rect 23664 26537 23673 26571
rect 23673 26537 23707 26571
rect 23707 26537 23716 26571
rect 23664 26528 23716 26537
rect 26240 26503 26292 26512
rect 26240 26469 26249 26503
rect 26249 26469 26283 26503
rect 26283 26469 26292 26503
rect 26240 26460 26292 26469
rect 21640 26367 21692 26376
rect 21640 26333 21649 26367
rect 21649 26333 21683 26367
rect 21683 26333 21692 26367
rect 21640 26324 21692 26333
rect 21824 26367 21876 26376
rect 21824 26333 21833 26367
rect 21833 26333 21867 26367
rect 21867 26333 21876 26367
rect 21824 26324 21876 26333
rect 24584 26392 24636 26444
rect 45008 26392 45060 26444
rect 46388 26392 46440 26444
rect 48044 26435 48096 26444
rect 48044 26401 48053 26435
rect 48053 26401 48087 26435
rect 48087 26401 48096 26435
rect 48044 26392 48096 26401
rect 23204 26324 23256 26376
rect 45836 26324 45888 26376
rect 46020 26324 46072 26376
rect 16212 26299 16264 26308
rect 16212 26265 16221 26299
rect 16221 26265 16255 26299
rect 16255 26265 16264 26299
rect 16212 26256 16264 26265
rect 22284 26256 22336 26308
rect 15936 26188 15988 26240
rect 16396 26231 16448 26240
rect 16396 26197 16405 26231
rect 16405 26197 16439 26231
rect 16439 26197 16448 26231
rect 16396 26188 16448 26197
rect 17040 26231 17092 26240
rect 17040 26197 17049 26231
rect 17049 26197 17083 26231
rect 17083 26197 17092 26231
rect 17040 26188 17092 26197
rect 18880 26188 18932 26240
rect 20996 26188 21048 26240
rect 22192 26188 22244 26240
rect 46388 26299 46440 26308
rect 46388 26265 46397 26299
rect 46397 26265 46431 26299
rect 46431 26265 46440 26299
rect 46388 26256 46440 26265
rect 22836 26188 22888 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 11152 25984 11204 26036
rect 13176 25984 13228 26036
rect 13820 26027 13872 26036
rect 13820 25993 13829 26027
rect 13829 25993 13863 26027
rect 13863 25993 13872 26027
rect 13820 25984 13872 25993
rect 16396 25984 16448 26036
rect 11428 25916 11480 25968
rect 10416 25848 10468 25900
rect 10968 25848 11020 25900
rect 11888 25891 11940 25900
rect 11888 25857 11897 25891
rect 11897 25857 11931 25891
rect 11931 25857 11940 25891
rect 11888 25848 11940 25857
rect 12808 25848 12860 25900
rect 13452 25916 13504 25968
rect 15660 25916 15712 25968
rect 20260 25984 20312 26036
rect 21272 26027 21324 26036
rect 21272 25993 21281 26027
rect 21281 25993 21315 26027
rect 21315 25993 21324 26027
rect 21272 25984 21324 25993
rect 22284 26027 22336 26036
rect 22284 25993 22293 26027
rect 22293 25993 22327 26027
rect 22327 25993 22336 26027
rect 22284 25984 22336 25993
rect 22376 25984 22428 26036
rect 27436 25984 27488 26036
rect 46388 25984 46440 26036
rect 46664 25984 46716 26036
rect 47584 25984 47636 26036
rect 17040 25916 17092 25968
rect 17960 25916 18012 25968
rect 20996 25916 21048 25968
rect 21824 25916 21876 25968
rect 13084 25848 13136 25900
rect 14004 25848 14056 25900
rect 15568 25848 15620 25900
rect 18880 25891 18932 25900
rect 18880 25857 18889 25891
rect 18889 25857 18923 25891
rect 18923 25857 18932 25891
rect 18880 25848 18932 25857
rect 11980 25780 12032 25832
rect 12992 25712 13044 25764
rect 16580 25780 16632 25832
rect 19984 25848 20036 25900
rect 21456 25848 21508 25900
rect 21916 25848 21968 25900
rect 23112 25848 23164 25900
rect 23204 25848 23256 25900
rect 45836 25848 45888 25900
rect 14096 25712 14148 25764
rect 16212 25712 16264 25764
rect 19064 25755 19116 25764
rect 19064 25721 19073 25755
rect 19073 25721 19107 25755
rect 19107 25721 19116 25755
rect 19064 25712 19116 25721
rect 19984 25712 20036 25764
rect 22284 25780 22336 25832
rect 47216 25780 47268 25832
rect 9404 25644 9456 25696
rect 19524 25644 19576 25696
rect 20260 25644 20312 25696
rect 24860 25644 24912 25696
rect 26056 25644 26108 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 16580 25483 16632 25492
rect 16580 25449 16589 25483
rect 16589 25449 16623 25483
rect 16623 25449 16632 25483
rect 16580 25440 16632 25449
rect 20996 25483 21048 25492
rect 20996 25449 21005 25483
rect 21005 25449 21039 25483
rect 21039 25449 21048 25483
rect 20996 25440 21048 25449
rect 21640 25483 21692 25492
rect 21640 25449 21649 25483
rect 21649 25449 21683 25483
rect 21683 25449 21692 25483
rect 21640 25440 21692 25449
rect 26700 25440 26752 25492
rect 9404 25347 9456 25356
rect 9404 25313 9413 25347
rect 9413 25313 9447 25347
rect 9447 25313 9456 25347
rect 9404 25304 9456 25313
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 18880 25372 18932 25424
rect 22008 25372 22060 25424
rect 22192 25372 22244 25424
rect 45836 25415 45888 25424
rect 45836 25381 45845 25415
rect 45845 25381 45879 25415
rect 45879 25381 45888 25415
rect 45836 25372 45888 25381
rect 13636 25304 13688 25356
rect 15568 25347 15620 25356
rect 15568 25313 15577 25347
rect 15577 25313 15611 25347
rect 15611 25313 15620 25347
rect 15568 25304 15620 25313
rect 19248 25347 19300 25356
rect 19248 25313 19257 25347
rect 19257 25313 19291 25347
rect 19291 25313 19300 25347
rect 19248 25304 19300 25313
rect 19524 25347 19576 25356
rect 19524 25313 19533 25347
rect 19533 25313 19567 25347
rect 19567 25313 19576 25347
rect 19524 25304 19576 25313
rect 23480 25304 23532 25356
rect 26976 25304 27028 25356
rect 48136 25347 48188 25356
rect 48136 25313 48145 25347
rect 48145 25313 48179 25347
rect 48179 25313 48188 25347
rect 48136 25304 48188 25313
rect 13912 25236 13964 25288
rect 15660 25236 15712 25288
rect 1676 25211 1728 25220
rect 1676 25177 1685 25211
rect 1685 25177 1719 25211
rect 1719 25177 1728 25211
rect 1676 25168 1728 25177
rect 9680 25211 9732 25220
rect 9680 25177 9689 25211
rect 9689 25177 9723 25211
rect 9723 25177 9732 25211
rect 9680 25168 9732 25177
rect 10416 25168 10468 25220
rect 11428 25211 11480 25220
rect 11428 25177 11437 25211
rect 11437 25177 11471 25211
rect 11471 25177 11480 25211
rect 11428 25168 11480 25177
rect 13728 25168 13780 25220
rect 14004 25168 14056 25220
rect 20996 25236 21048 25288
rect 21916 25236 21968 25288
rect 16580 25168 16632 25220
rect 20260 25168 20312 25220
rect 14096 25100 14148 25152
rect 15844 25100 15896 25152
rect 24492 25236 24544 25288
rect 25044 25236 25096 25288
rect 45744 25236 45796 25288
rect 46296 25279 46348 25288
rect 46296 25245 46305 25279
rect 46305 25245 46339 25279
rect 46339 25245 46348 25279
rect 46296 25236 46348 25245
rect 22652 25211 22704 25220
rect 22652 25177 22661 25211
rect 22661 25177 22695 25211
rect 22695 25177 22704 25211
rect 22652 25168 22704 25177
rect 22836 25211 22888 25220
rect 22836 25177 22845 25211
rect 22845 25177 22879 25211
rect 22879 25177 22888 25211
rect 22836 25168 22888 25177
rect 23756 25100 23808 25152
rect 26056 25168 26108 25220
rect 47676 25168 47728 25220
rect 26424 25100 26476 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 22652 24896 22704 24948
rect 25228 24939 25280 24948
rect 25228 24905 25237 24939
rect 25237 24905 25271 24939
rect 25271 24905 25280 24939
rect 25228 24896 25280 24905
rect 46204 24896 46256 24948
rect 46756 24896 46808 24948
rect 14096 24828 14148 24880
rect 23756 24871 23808 24880
rect 23756 24837 23765 24871
rect 23765 24837 23799 24871
rect 23799 24837 23808 24871
rect 23756 24828 23808 24837
rect 11428 24760 11480 24812
rect 9956 24735 10008 24744
rect 9956 24701 9965 24735
rect 9965 24701 9999 24735
rect 9999 24701 10008 24735
rect 9956 24692 10008 24701
rect 10968 24692 11020 24744
rect 13084 24735 13136 24744
rect 13084 24701 13093 24735
rect 13093 24701 13127 24735
rect 13127 24701 13136 24735
rect 13084 24692 13136 24701
rect 13360 24735 13412 24744
rect 13360 24701 13369 24735
rect 13369 24701 13403 24735
rect 13403 24701 13412 24735
rect 13360 24692 13412 24701
rect 17960 24760 18012 24812
rect 18880 24760 18932 24812
rect 19984 24803 20036 24812
rect 19984 24769 19993 24803
rect 19993 24769 20027 24803
rect 20027 24769 20036 24803
rect 19984 24760 20036 24769
rect 22192 24803 22244 24812
rect 22192 24769 22201 24803
rect 22201 24769 22235 24803
rect 22235 24769 22244 24803
rect 22192 24760 22244 24769
rect 22468 24803 22520 24812
rect 22468 24769 22477 24803
rect 22477 24769 22511 24803
rect 22511 24769 22520 24803
rect 23480 24803 23532 24812
rect 22468 24760 22520 24769
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 24860 24760 24912 24812
rect 45560 24828 45612 24880
rect 24768 24692 24820 24744
rect 47492 24760 47544 24812
rect 47676 24803 47728 24812
rect 47676 24769 47685 24803
rect 47685 24769 47719 24803
rect 47719 24769 47728 24803
rect 47676 24760 47728 24769
rect 45376 24735 45428 24744
rect 9680 24624 9732 24676
rect 10968 24556 11020 24608
rect 15752 24624 15804 24676
rect 16488 24624 16540 24676
rect 17960 24624 18012 24676
rect 15476 24556 15528 24608
rect 19156 24556 19208 24608
rect 22836 24624 22888 24676
rect 23388 24624 23440 24676
rect 20352 24556 20404 24608
rect 22008 24599 22060 24608
rect 22008 24565 22017 24599
rect 22017 24565 22051 24599
rect 22051 24565 22060 24599
rect 22008 24556 22060 24565
rect 45376 24701 45385 24735
rect 45385 24701 45419 24735
rect 45419 24701 45428 24735
rect 45376 24692 45428 24701
rect 46848 24735 46900 24744
rect 46848 24701 46857 24735
rect 46857 24701 46891 24735
rect 46891 24701 46900 24735
rect 46848 24692 46900 24701
rect 46848 24556 46900 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 10416 24352 10468 24404
rect 13360 24352 13412 24404
rect 21916 24352 21968 24404
rect 24952 24352 25004 24404
rect 25136 24352 25188 24404
rect 10416 24191 10468 24200
rect 10416 24157 10425 24191
rect 10425 24157 10459 24191
rect 10459 24157 10468 24191
rect 10416 24148 10468 24157
rect 12992 24284 13044 24336
rect 13084 24284 13136 24336
rect 20996 24284 21048 24336
rect 40776 24284 40828 24336
rect 12808 24259 12860 24268
rect 12808 24225 12817 24259
rect 12817 24225 12851 24259
rect 12851 24225 12860 24259
rect 12808 24216 12860 24225
rect 15476 24216 15528 24268
rect 16580 24216 16632 24268
rect 12808 24080 12860 24132
rect 12992 24148 13044 24200
rect 12992 24012 13044 24064
rect 14004 24148 14056 24200
rect 15752 24148 15804 24200
rect 16028 24191 16080 24200
rect 16028 24157 16037 24191
rect 16037 24157 16071 24191
rect 16071 24157 16080 24191
rect 16028 24148 16080 24157
rect 16396 24191 16448 24200
rect 16396 24157 16405 24191
rect 16405 24157 16439 24191
rect 16439 24157 16448 24191
rect 16396 24148 16448 24157
rect 16488 24191 16540 24200
rect 16488 24157 16497 24191
rect 16497 24157 16531 24191
rect 16531 24157 16540 24191
rect 19248 24216 19300 24268
rect 22008 24216 22060 24268
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 16488 24148 16540 24157
rect 17960 24191 18012 24200
rect 17960 24157 17969 24191
rect 17969 24157 18003 24191
rect 18003 24157 18012 24191
rect 17960 24148 18012 24157
rect 13728 24080 13780 24132
rect 14740 24012 14792 24064
rect 16304 24055 16356 24064
rect 16304 24021 16313 24055
rect 16313 24021 16347 24055
rect 16347 24021 16356 24055
rect 16304 24012 16356 24021
rect 16672 24012 16724 24064
rect 18052 24055 18104 24064
rect 18052 24021 18061 24055
rect 18061 24021 18095 24055
rect 18095 24021 18104 24055
rect 18052 24012 18104 24021
rect 20352 24080 20404 24132
rect 24768 24148 24820 24200
rect 24860 24148 24912 24200
rect 22284 24012 22336 24064
rect 23664 24012 23716 24064
rect 25504 24080 25556 24132
rect 28816 24148 28868 24200
rect 29736 24123 29788 24132
rect 29736 24089 29745 24123
rect 29745 24089 29779 24123
rect 29779 24089 29788 24123
rect 29736 24080 29788 24089
rect 40040 24080 40092 24132
rect 47676 24080 47728 24132
rect 26976 24012 27028 24064
rect 27344 24055 27396 24064
rect 27344 24021 27353 24055
rect 27353 24021 27387 24055
rect 27387 24021 27396 24055
rect 27344 24012 27396 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 11888 23740 11940 23792
rect 10324 23715 10376 23724
rect 10324 23681 10333 23715
rect 10333 23681 10367 23715
rect 10367 23681 10376 23715
rect 10324 23672 10376 23681
rect 13728 23808 13780 23860
rect 15936 23851 15988 23860
rect 15936 23817 15945 23851
rect 15945 23817 15979 23851
rect 15979 23817 15988 23851
rect 15936 23808 15988 23817
rect 16396 23808 16448 23860
rect 17960 23808 18012 23860
rect 22284 23808 22336 23860
rect 12992 23783 13044 23792
rect 12992 23749 13001 23783
rect 13001 23749 13035 23783
rect 13035 23749 13044 23783
rect 12992 23740 13044 23749
rect 15476 23740 15528 23792
rect 16304 23740 16356 23792
rect 12808 23715 12860 23724
rect 7656 23647 7708 23656
rect 7656 23613 7665 23647
rect 7665 23613 7699 23647
rect 7699 23613 7708 23647
rect 7656 23604 7708 23613
rect 7932 23647 7984 23656
rect 7932 23613 7941 23647
rect 7941 23613 7975 23647
rect 7975 23613 7984 23647
rect 7932 23604 7984 23613
rect 11888 23604 11940 23656
rect 12808 23681 12817 23715
rect 12817 23681 12851 23715
rect 12851 23681 12860 23715
rect 12808 23672 12860 23681
rect 16672 23715 16724 23724
rect 13820 23647 13872 23656
rect 13820 23613 13829 23647
rect 13829 23613 13863 23647
rect 13863 23613 13872 23647
rect 13820 23604 13872 23613
rect 16672 23681 16681 23715
rect 16681 23681 16715 23715
rect 16715 23681 16724 23715
rect 16672 23672 16724 23681
rect 18052 23672 18104 23724
rect 22100 23715 22152 23724
rect 22100 23681 22109 23715
rect 22109 23681 22143 23715
rect 22143 23681 22152 23715
rect 22100 23672 22152 23681
rect 16120 23604 16172 23656
rect 15292 23536 15344 23588
rect 16672 23536 16724 23588
rect 10324 23511 10376 23520
rect 10324 23477 10333 23511
rect 10333 23477 10367 23511
rect 10367 23477 10376 23511
rect 10324 23468 10376 23477
rect 12256 23511 12308 23520
rect 12256 23477 12265 23511
rect 12265 23477 12299 23511
rect 12299 23477 12308 23511
rect 12256 23468 12308 23477
rect 19340 23647 19392 23656
rect 19340 23613 19349 23647
rect 19349 23613 19383 23647
rect 19383 23613 19392 23647
rect 19340 23604 19392 23613
rect 20812 23604 20864 23656
rect 23664 23715 23716 23724
rect 23020 23604 23072 23656
rect 23664 23681 23673 23715
rect 23673 23681 23707 23715
rect 23707 23681 23716 23715
rect 23664 23672 23716 23681
rect 24860 23672 24912 23724
rect 25688 23715 25740 23724
rect 25688 23681 25697 23715
rect 25697 23681 25731 23715
rect 25731 23681 25740 23715
rect 25688 23672 25740 23681
rect 26148 23715 26200 23724
rect 26148 23681 26157 23715
rect 26157 23681 26191 23715
rect 26191 23681 26200 23715
rect 26148 23672 26200 23681
rect 26240 23672 26292 23724
rect 27252 23740 27304 23792
rect 27344 23740 27396 23792
rect 37280 23740 37332 23792
rect 40776 23851 40828 23860
rect 40776 23817 40785 23851
rect 40785 23817 40819 23851
rect 40819 23817 40828 23851
rect 40776 23808 40828 23817
rect 45376 23808 45428 23860
rect 47676 23851 47728 23860
rect 47676 23817 47685 23851
rect 47685 23817 47719 23851
rect 47719 23817 47728 23851
rect 47676 23808 47728 23817
rect 46572 23740 46624 23792
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 40776 23672 40828 23724
rect 28816 23604 28868 23656
rect 29000 23604 29052 23656
rect 29920 23647 29972 23656
rect 29920 23613 29929 23647
rect 29929 23613 29963 23647
rect 29963 23613 29972 23647
rect 29920 23604 29972 23613
rect 41420 23672 41472 23724
rect 46756 23672 46808 23724
rect 47124 23672 47176 23724
rect 47584 23715 47636 23724
rect 47584 23681 47593 23715
rect 47593 23681 47627 23715
rect 47627 23681 47636 23715
rect 47584 23672 47636 23681
rect 45744 23536 45796 23588
rect 20812 23468 20864 23520
rect 21180 23468 21232 23520
rect 22284 23468 22336 23520
rect 22928 23511 22980 23520
rect 22928 23477 22937 23511
rect 22937 23477 22971 23511
rect 22971 23477 22980 23511
rect 22928 23468 22980 23477
rect 23572 23468 23624 23520
rect 24492 23511 24544 23520
rect 24492 23477 24501 23511
rect 24501 23477 24535 23511
rect 24535 23477 24544 23511
rect 24492 23468 24544 23477
rect 41328 23468 41380 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 7656 23264 7708 23316
rect 16028 23264 16080 23316
rect 16580 23264 16632 23316
rect 15476 23239 15528 23248
rect 15476 23205 15485 23239
rect 15485 23205 15519 23239
rect 15519 23205 15528 23239
rect 15476 23196 15528 23205
rect 15752 23196 15804 23248
rect 2136 23128 2188 23180
rect 16580 23128 16632 23180
rect 7656 23103 7708 23112
rect 7656 23069 7665 23103
rect 7665 23069 7699 23103
rect 7699 23069 7708 23103
rect 7656 23060 7708 23069
rect 9680 23103 9732 23112
rect 8944 22924 8996 22976
rect 9680 23069 9689 23103
rect 9689 23069 9723 23103
rect 9723 23069 9732 23103
rect 9680 23060 9732 23069
rect 9956 23060 10008 23112
rect 10324 23103 10376 23112
rect 10324 23069 10333 23103
rect 10333 23069 10367 23103
rect 10367 23069 10376 23103
rect 10324 23060 10376 23069
rect 11980 23060 12032 23112
rect 10232 22924 10284 22976
rect 11520 22924 11572 22976
rect 12256 22924 12308 22976
rect 13912 23060 13964 23112
rect 14004 23060 14056 23112
rect 15844 23103 15896 23112
rect 15844 23069 15853 23103
rect 15853 23069 15887 23103
rect 15887 23069 15896 23103
rect 15844 23060 15896 23069
rect 16672 23103 16724 23112
rect 16672 23069 16681 23103
rect 16681 23069 16715 23103
rect 16715 23069 16724 23103
rect 16672 23060 16724 23069
rect 16580 22992 16632 23044
rect 13452 22967 13504 22976
rect 13452 22933 13461 22967
rect 13461 22933 13495 22967
rect 13495 22933 13504 22967
rect 13452 22924 13504 22933
rect 14372 22924 14424 22976
rect 15844 22924 15896 22976
rect 16028 22967 16080 22976
rect 16028 22933 16037 22967
rect 16037 22933 16071 22967
rect 16071 22933 16080 22967
rect 21364 23171 21416 23180
rect 21364 23137 21373 23171
rect 21373 23137 21407 23171
rect 21407 23137 21416 23171
rect 21364 23128 21416 23137
rect 22928 23264 22980 23316
rect 29736 23264 29788 23316
rect 22284 23171 22336 23180
rect 22284 23137 22293 23171
rect 22293 23137 22327 23171
rect 22327 23137 22336 23171
rect 22284 23128 22336 23137
rect 24492 23128 24544 23180
rect 26240 23128 26292 23180
rect 20536 23060 20588 23112
rect 20720 23103 20772 23112
rect 20720 23069 20729 23103
rect 20729 23069 20763 23103
rect 20763 23069 20772 23103
rect 20720 23060 20772 23069
rect 26148 23060 26200 23112
rect 27344 23128 27396 23180
rect 38292 23196 38344 23248
rect 47308 23171 47360 23180
rect 47308 23137 47317 23171
rect 47317 23137 47351 23171
rect 47351 23137 47360 23171
rect 47308 23128 47360 23137
rect 18604 23035 18656 23044
rect 18604 23001 18613 23035
rect 18613 23001 18647 23035
rect 18647 23001 18656 23035
rect 18604 22992 18656 23001
rect 18972 22992 19024 23044
rect 19432 22992 19484 23044
rect 22192 22992 22244 23044
rect 16028 22924 16080 22933
rect 16856 22967 16908 22976
rect 16856 22933 16865 22967
rect 16865 22933 16899 22967
rect 16899 22933 16908 22967
rect 23572 22992 23624 23044
rect 24860 23035 24912 23044
rect 24860 23001 24869 23035
rect 24869 23001 24903 23035
rect 24903 23001 24912 23035
rect 24860 22992 24912 23001
rect 25596 22992 25648 23044
rect 16856 22924 16908 22933
rect 26240 22992 26292 23044
rect 26976 22992 27028 23044
rect 28632 23060 28684 23112
rect 28908 23060 28960 23112
rect 41328 23060 41380 23112
rect 46940 23060 46992 23112
rect 26332 22967 26384 22976
rect 26332 22933 26341 22967
rect 26341 22933 26375 22967
rect 26375 22933 26384 22967
rect 26332 22924 26384 22933
rect 27436 22967 27488 22976
rect 27436 22933 27445 22967
rect 27445 22933 27479 22967
rect 27479 22933 27488 22967
rect 27436 22924 27488 22933
rect 27528 22924 27580 22976
rect 28264 22967 28316 22976
rect 28264 22933 28273 22967
rect 28273 22933 28307 22967
rect 28307 22933 28316 22967
rect 28264 22924 28316 22933
rect 28816 22924 28868 22976
rect 29552 22924 29604 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 3700 22720 3752 22772
rect 7472 22584 7524 22636
rect 9312 22516 9364 22568
rect 3516 22448 3568 22500
rect 9956 22423 10008 22432
rect 9956 22389 9965 22423
rect 9965 22389 9999 22423
rect 9999 22389 10008 22423
rect 9956 22380 10008 22389
rect 10232 22720 10284 22772
rect 16120 22763 16172 22772
rect 16120 22729 16129 22763
rect 16129 22729 16163 22763
rect 16163 22729 16172 22763
rect 16120 22720 16172 22729
rect 16856 22720 16908 22772
rect 19340 22720 19392 22772
rect 13452 22652 13504 22704
rect 11428 22584 11480 22636
rect 14372 22627 14424 22636
rect 14372 22593 14381 22627
rect 14381 22593 14415 22627
rect 14415 22593 14424 22627
rect 14372 22584 14424 22593
rect 18604 22652 18656 22704
rect 46756 22720 46808 22772
rect 47768 22720 47820 22772
rect 25596 22695 25648 22704
rect 25596 22661 25605 22695
rect 25605 22661 25639 22695
rect 25639 22661 25648 22695
rect 25596 22652 25648 22661
rect 25688 22652 25740 22704
rect 19616 22584 19668 22636
rect 19984 22584 20036 22636
rect 20996 22627 21048 22636
rect 20996 22593 21005 22627
rect 21005 22593 21039 22627
rect 21039 22593 21048 22627
rect 20996 22584 21048 22593
rect 11520 22559 11572 22568
rect 11520 22525 11529 22559
rect 11529 22525 11563 22559
rect 11563 22525 11572 22559
rect 11520 22516 11572 22525
rect 11704 22559 11756 22568
rect 11704 22525 11713 22559
rect 11713 22525 11747 22559
rect 11747 22525 11756 22559
rect 11704 22516 11756 22525
rect 15936 22516 15988 22568
rect 17592 22559 17644 22568
rect 17592 22525 17601 22559
rect 17601 22525 17635 22559
rect 17635 22525 17644 22559
rect 17592 22516 17644 22525
rect 19156 22559 19208 22568
rect 19156 22525 19165 22559
rect 19165 22525 19199 22559
rect 19199 22525 19208 22559
rect 19156 22516 19208 22525
rect 10416 22380 10468 22432
rect 11980 22380 12032 22432
rect 20260 22423 20312 22432
rect 20260 22389 20269 22423
rect 20269 22389 20303 22423
rect 20303 22389 20312 22423
rect 20260 22380 20312 22389
rect 20720 22380 20772 22432
rect 22836 22584 22888 22636
rect 24216 22584 24268 22636
rect 22560 22516 22612 22568
rect 24860 22516 24912 22568
rect 25504 22627 25556 22636
rect 25504 22593 25513 22627
rect 25513 22593 25547 22627
rect 25547 22593 25556 22627
rect 25504 22584 25556 22593
rect 26148 22627 26200 22636
rect 26148 22593 26157 22627
rect 26157 22593 26191 22627
rect 26191 22593 26200 22627
rect 27436 22652 27488 22704
rect 27712 22652 27764 22704
rect 28356 22652 28408 22704
rect 29920 22652 29972 22704
rect 26148 22584 26200 22593
rect 26240 22516 26292 22568
rect 27252 22627 27304 22636
rect 27252 22593 27261 22627
rect 27261 22593 27295 22627
rect 27295 22593 27304 22627
rect 27252 22584 27304 22593
rect 27620 22584 27672 22636
rect 28448 22584 28500 22636
rect 28632 22584 28684 22636
rect 29552 22627 29604 22636
rect 29552 22593 29561 22627
rect 29561 22593 29595 22627
rect 29595 22593 29604 22627
rect 29552 22584 29604 22593
rect 28264 22516 28316 22568
rect 25688 22448 25740 22500
rect 26056 22448 26108 22500
rect 26976 22448 27028 22500
rect 29000 22448 29052 22500
rect 45836 22584 45888 22636
rect 46848 22584 46900 22636
rect 46572 22516 46624 22568
rect 23204 22423 23256 22432
rect 23204 22389 23213 22423
rect 23213 22389 23247 22423
rect 23247 22389 23256 22423
rect 23204 22380 23256 22389
rect 26608 22380 26660 22432
rect 26884 22380 26936 22432
rect 27528 22380 27580 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 11704 22176 11756 22228
rect 11796 22176 11848 22228
rect 14004 22176 14056 22228
rect 17592 22219 17644 22228
rect 17592 22185 17601 22219
rect 17601 22185 17635 22219
rect 17635 22185 17644 22219
rect 17592 22176 17644 22185
rect 22836 22219 22888 22228
rect 22836 22185 22845 22219
rect 22845 22185 22879 22219
rect 22879 22185 22888 22219
rect 22836 22176 22888 22185
rect 43168 22176 43220 22228
rect 8944 22083 8996 22092
rect 8944 22049 8953 22083
rect 8953 22049 8987 22083
rect 8987 22049 8996 22083
rect 8944 22040 8996 22049
rect 11428 22040 11480 22092
rect 12256 22040 12308 22092
rect 7564 22015 7616 22024
rect 7564 21981 7573 22015
rect 7573 21981 7607 22015
rect 7607 21981 7616 22015
rect 7564 21972 7616 21981
rect 11152 22015 11204 22024
rect 11152 21981 11161 22015
rect 11161 21981 11195 22015
rect 11195 21981 11204 22015
rect 11152 21972 11204 21981
rect 11888 21972 11940 22024
rect 16028 22108 16080 22160
rect 22560 22108 22612 22160
rect 27252 22108 27304 22160
rect 15936 22083 15988 22092
rect 15936 22049 15945 22083
rect 15945 22049 15979 22083
rect 15979 22049 15988 22083
rect 15936 22040 15988 22049
rect 16672 22040 16724 22092
rect 20812 22040 20864 22092
rect 23940 22040 23992 22092
rect 27620 22040 27672 22092
rect 29000 22083 29052 22092
rect 29000 22049 29009 22083
rect 29009 22049 29043 22083
rect 29043 22049 29052 22083
rect 29000 22040 29052 22049
rect 46940 22040 46992 22092
rect 47124 22083 47176 22092
rect 47124 22049 47133 22083
rect 47133 22049 47167 22083
rect 47167 22049 47176 22083
rect 47124 22040 47176 22049
rect 47768 22040 47820 22092
rect 16120 21972 16172 22024
rect 17500 22015 17552 22024
rect 17500 21981 17509 22015
rect 17509 21981 17543 22015
rect 17543 21981 17552 22015
rect 17500 21972 17552 21981
rect 19616 21972 19668 22024
rect 20168 21972 20220 22024
rect 24768 22015 24820 22024
rect 9220 21947 9272 21956
rect 9220 21913 9229 21947
rect 9229 21913 9263 21947
rect 9263 21913 9272 21947
rect 9220 21904 9272 21913
rect 9956 21904 10008 21956
rect 11520 21904 11572 21956
rect 14924 21904 14976 21956
rect 7472 21836 7524 21888
rect 9312 21836 9364 21888
rect 11704 21836 11756 21888
rect 11980 21879 12032 21888
rect 11980 21845 11989 21879
rect 11989 21845 12023 21879
rect 12023 21845 12032 21879
rect 11980 21836 12032 21845
rect 13636 21836 13688 21888
rect 24768 21981 24777 22015
rect 24777 21981 24811 22015
rect 24811 21981 24820 22015
rect 24768 21972 24820 21981
rect 26608 22015 26660 22024
rect 26608 21981 26617 22015
rect 26617 21981 26651 22015
rect 26651 21981 26660 22015
rect 26608 21972 26660 21981
rect 26884 21972 26936 22024
rect 27252 22015 27304 22024
rect 27252 21981 27261 22015
rect 27261 21981 27295 22015
rect 27295 21981 27304 22015
rect 27252 21972 27304 21981
rect 20812 21904 20864 21956
rect 21088 21904 21140 21956
rect 28540 21904 28592 21956
rect 46756 21904 46808 21956
rect 21548 21836 21600 21888
rect 26976 21836 27028 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 9128 21632 9180 21684
rect 9220 21632 9272 21684
rect 9772 21675 9824 21684
rect 9772 21641 9781 21675
rect 9781 21641 9815 21675
rect 9815 21641 9824 21675
rect 9772 21632 9824 21641
rect 7472 21607 7524 21616
rect 7472 21573 7481 21607
rect 7481 21573 7515 21607
rect 7515 21573 7524 21607
rect 7472 21564 7524 21573
rect 7564 21564 7616 21616
rect 17500 21632 17552 21684
rect 20168 21632 20220 21684
rect 11520 21564 11572 21616
rect 20 21360 72 21412
rect 9312 21428 9364 21480
rect 10232 21471 10284 21480
rect 10232 21437 10241 21471
rect 10241 21437 10275 21471
rect 10275 21437 10284 21471
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 11888 21496 11940 21548
rect 12348 21496 12400 21548
rect 14740 21496 14792 21548
rect 16672 21539 16724 21548
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 18972 21564 19024 21616
rect 20260 21564 20312 21616
rect 20996 21564 21048 21616
rect 26976 21632 27028 21684
rect 27252 21632 27304 21684
rect 28540 21675 28592 21684
rect 28540 21641 28549 21675
rect 28549 21641 28583 21675
rect 28583 21641 28592 21675
rect 28540 21632 28592 21641
rect 47952 21607 48004 21616
rect 23940 21539 23992 21548
rect 23940 21505 23949 21539
rect 23949 21505 23983 21539
rect 23983 21505 23992 21539
rect 23940 21496 23992 21505
rect 24860 21496 24912 21548
rect 26700 21496 26752 21548
rect 47952 21573 47961 21607
rect 47961 21573 47995 21607
rect 47995 21573 48004 21607
rect 47952 21564 48004 21573
rect 10232 21428 10284 21437
rect 11060 21428 11112 21480
rect 11796 21428 11848 21480
rect 16580 21428 16632 21480
rect 17408 21428 17460 21480
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 18972 21428 19024 21480
rect 22376 21428 22428 21480
rect 22560 21471 22612 21480
rect 22560 21437 22569 21471
rect 22569 21437 22603 21471
rect 22603 21437 22612 21471
rect 22560 21428 22612 21437
rect 27528 21428 27580 21480
rect 9680 21360 9732 21412
rect 46480 21360 46532 21412
rect 9772 21292 9824 21344
rect 10324 21292 10376 21344
rect 10968 21292 11020 21344
rect 11980 21292 12032 21344
rect 12256 21292 12308 21344
rect 20444 21292 20496 21344
rect 24768 21292 24820 21344
rect 25320 21335 25372 21344
rect 25320 21301 25329 21335
rect 25329 21301 25363 21335
rect 25363 21301 25372 21335
rect 25320 21292 25372 21301
rect 25964 21292 26016 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 10600 21088 10652 21140
rect 10784 21131 10836 21140
rect 10784 21097 10793 21131
rect 10793 21097 10827 21131
rect 10827 21097 10836 21131
rect 10784 21088 10836 21097
rect 10968 21088 11020 21140
rect 14924 21131 14976 21140
rect 14924 21097 14933 21131
rect 14933 21097 14967 21131
rect 14967 21097 14976 21131
rect 14924 21088 14976 21097
rect 18880 21088 18932 21140
rect 11060 21020 11112 21072
rect 11152 21020 11204 21072
rect 20352 21020 20404 21072
rect 3608 20952 3660 21004
rect 23020 21088 23072 21140
rect 26700 21088 26752 21140
rect 14096 20927 14148 20936
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 18420 20884 18472 20936
rect 19248 20927 19300 20936
rect 19248 20893 19257 20927
rect 19257 20893 19291 20927
rect 19291 20893 19300 20927
rect 19248 20884 19300 20893
rect 20168 20884 20220 20936
rect 9312 20816 9364 20868
rect 10600 20859 10652 20868
rect 10600 20825 10609 20859
rect 10609 20825 10643 20859
rect 10643 20825 10652 20859
rect 10600 20816 10652 20825
rect 14740 20859 14792 20868
rect 9680 20748 9732 20800
rect 10232 20748 10284 20800
rect 14188 20791 14240 20800
rect 14188 20757 14197 20791
rect 14197 20757 14231 20791
rect 14231 20757 14240 20791
rect 14188 20748 14240 20757
rect 14740 20825 14749 20859
rect 14749 20825 14783 20859
rect 14783 20825 14792 20859
rect 14740 20816 14792 20825
rect 15660 20816 15712 20868
rect 20444 20884 20496 20936
rect 21088 20927 21140 20936
rect 21088 20893 21097 20927
rect 21097 20893 21131 20927
rect 21131 20893 21140 20927
rect 21088 20884 21140 20893
rect 26884 20952 26936 21004
rect 27436 20995 27488 21004
rect 27436 20961 27445 20995
rect 27445 20961 27479 20995
rect 27479 20961 27488 20995
rect 27436 20952 27488 20961
rect 28080 20952 28132 21004
rect 32220 20995 32272 21004
rect 32220 20961 32229 20995
rect 32229 20961 32263 20995
rect 32263 20961 32272 20995
rect 32220 20952 32272 20961
rect 47768 20952 47820 21004
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 23388 20884 23440 20936
rect 26700 20927 26752 20936
rect 22192 20816 22244 20868
rect 26700 20893 26709 20927
rect 26709 20893 26743 20927
rect 26743 20893 26752 20927
rect 26700 20884 26752 20893
rect 27252 20884 27304 20936
rect 29552 20884 29604 20936
rect 18604 20748 18656 20800
rect 21180 20748 21232 20800
rect 24400 20748 24452 20800
rect 24768 20816 24820 20868
rect 30564 20859 30616 20868
rect 30564 20825 30573 20859
rect 30573 20825 30607 20859
rect 30607 20825 30616 20859
rect 30564 20816 30616 20825
rect 46480 20859 46532 20868
rect 46480 20825 46489 20859
rect 46489 20825 46523 20859
rect 46523 20825 46532 20859
rect 46480 20816 46532 20825
rect 24860 20748 24912 20800
rect 26148 20748 26200 20800
rect 27804 20748 27856 20800
rect 46296 20748 46348 20800
rect 47308 20748 47360 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 10600 20544 10652 20596
rect 13084 20544 13136 20596
rect 21364 20544 21416 20596
rect 29552 20587 29604 20596
rect 14188 20476 14240 20528
rect 9680 20340 9732 20392
rect 10324 20451 10376 20460
rect 10324 20417 10333 20451
rect 10333 20417 10367 20451
rect 10367 20417 10376 20451
rect 10324 20408 10376 20417
rect 10784 20340 10836 20392
rect 11612 20340 11664 20392
rect 12348 20383 12400 20392
rect 12348 20349 12357 20383
rect 12357 20349 12391 20383
rect 12391 20349 12400 20383
rect 12348 20340 12400 20349
rect 12440 20340 12492 20392
rect 15844 20408 15896 20460
rect 21180 20476 21232 20528
rect 18420 20408 18472 20460
rect 18604 20451 18656 20460
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 20168 20408 20220 20460
rect 22100 20476 22152 20528
rect 24400 20519 24452 20528
rect 24400 20485 24409 20519
rect 24409 20485 24443 20519
rect 24443 20485 24452 20519
rect 24400 20476 24452 20485
rect 28080 20519 28132 20528
rect 28080 20485 28089 20519
rect 28089 20485 28123 20519
rect 28123 20485 28132 20519
rect 28080 20476 28132 20485
rect 28632 20476 28684 20528
rect 29552 20553 29561 20587
rect 29561 20553 29595 20587
rect 29595 20553 29604 20587
rect 29552 20544 29604 20553
rect 30564 20587 30616 20596
rect 30564 20553 30573 20587
rect 30573 20553 30607 20587
rect 30607 20553 30616 20587
rect 30564 20544 30616 20553
rect 30104 20476 30156 20528
rect 24216 20451 24268 20460
rect 24216 20417 24225 20451
rect 24225 20417 24259 20451
rect 24259 20417 24268 20451
rect 24216 20408 24268 20417
rect 26976 20451 27028 20460
rect 26976 20417 26985 20451
rect 26985 20417 27019 20451
rect 27019 20417 27028 20451
rect 26976 20408 27028 20417
rect 27620 20408 27672 20460
rect 27804 20451 27856 20460
rect 27804 20417 27813 20451
rect 27813 20417 27847 20451
rect 27847 20417 27856 20451
rect 27804 20408 27856 20417
rect 30472 20451 30524 20460
rect 30472 20417 30481 20451
rect 30481 20417 30515 20451
rect 30515 20417 30524 20451
rect 46388 20544 46440 20596
rect 46480 20544 46532 20596
rect 46296 20476 46348 20528
rect 30472 20408 30524 20417
rect 45928 20451 45980 20460
rect 18512 20340 18564 20392
rect 21364 20340 21416 20392
rect 22284 20340 22336 20392
rect 26056 20383 26108 20392
rect 13912 20272 13964 20324
rect 26056 20349 26065 20383
rect 26065 20349 26099 20383
rect 26099 20349 26108 20383
rect 26056 20340 26108 20349
rect 45928 20417 45937 20451
rect 45937 20417 45971 20451
rect 45971 20417 45980 20451
rect 45928 20408 45980 20417
rect 46480 20408 46532 20460
rect 47768 20451 47820 20460
rect 47768 20417 47777 20451
rect 47777 20417 47811 20451
rect 47811 20417 47820 20451
rect 47768 20408 47820 20417
rect 9956 20204 10008 20256
rect 14096 20204 14148 20256
rect 14188 20204 14240 20256
rect 14464 20247 14516 20256
rect 14464 20213 14473 20247
rect 14473 20213 14507 20247
rect 14507 20213 14516 20247
rect 14464 20204 14516 20213
rect 15936 20204 15988 20256
rect 17224 20247 17276 20256
rect 17224 20213 17233 20247
rect 17233 20213 17267 20247
rect 17267 20213 17276 20247
rect 17224 20204 17276 20213
rect 17500 20204 17552 20256
rect 18788 20204 18840 20256
rect 23388 20204 23440 20256
rect 25780 20204 25832 20256
rect 27068 20247 27120 20256
rect 27068 20213 27077 20247
rect 27077 20213 27111 20247
rect 27111 20213 27120 20247
rect 27068 20204 27120 20213
rect 45192 20247 45244 20256
rect 45192 20213 45201 20247
rect 45201 20213 45235 20247
rect 45235 20213 45244 20247
rect 45192 20204 45244 20213
rect 45744 20247 45796 20256
rect 45744 20213 45753 20247
rect 45753 20213 45787 20247
rect 45787 20213 45796 20247
rect 45744 20204 45796 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 11612 20043 11664 20052
rect 11612 20009 11621 20043
rect 11621 20009 11655 20043
rect 11655 20009 11664 20043
rect 11612 20000 11664 20009
rect 12348 20000 12400 20052
rect 14924 20000 14976 20052
rect 26148 20043 26200 20052
rect 9956 19975 10008 19984
rect 9956 19941 9965 19975
rect 9965 19941 9999 19975
rect 9999 19941 10008 19975
rect 9956 19932 10008 19941
rect 3976 19864 4028 19916
rect 13912 19932 13964 19984
rect 14096 19975 14148 19984
rect 14096 19941 14105 19975
rect 14105 19941 14139 19975
rect 14139 19941 14148 19975
rect 14096 19932 14148 19941
rect 10324 19864 10376 19916
rect 1768 19796 1820 19848
rect 10232 19796 10284 19848
rect 10600 19796 10652 19848
rect 14004 19864 14056 19916
rect 15936 19907 15988 19916
rect 15936 19873 15945 19907
rect 15945 19873 15979 19907
rect 15979 19873 15988 19907
rect 15936 19864 15988 19873
rect 18420 19932 18472 19984
rect 20260 19932 20312 19984
rect 18328 19907 18380 19916
rect 18328 19873 18337 19907
rect 18337 19873 18371 19907
rect 18371 19873 18380 19907
rect 18328 19864 18380 19873
rect 23388 19907 23440 19916
rect 23388 19873 23397 19907
rect 23397 19873 23431 19907
rect 23431 19873 23440 19907
rect 23388 19864 23440 19873
rect 25320 19864 25372 19916
rect 26148 20009 26157 20043
rect 26157 20009 26191 20043
rect 26191 20009 26200 20043
rect 26148 20000 26200 20009
rect 27528 20043 27580 20052
rect 27528 20009 27537 20043
rect 27537 20009 27571 20043
rect 27571 20009 27580 20043
rect 27528 20000 27580 20009
rect 28632 20043 28684 20052
rect 28632 20009 28641 20043
rect 28641 20009 28675 20043
rect 28675 20009 28684 20043
rect 28632 20000 28684 20009
rect 25780 19932 25832 19984
rect 30472 19932 30524 19984
rect 46204 20000 46256 20052
rect 45192 19932 45244 19984
rect 45560 19864 45612 19916
rect 45744 19864 45796 19916
rect 47032 19864 47084 19916
rect 9128 19728 9180 19780
rect 10784 19660 10836 19712
rect 12072 19728 12124 19780
rect 13452 19660 13504 19712
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 18420 19839 18472 19848
rect 18420 19805 18429 19839
rect 18429 19805 18463 19839
rect 18463 19805 18472 19839
rect 18420 19796 18472 19805
rect 14740 19728 14792 19780
rect 17132 19728 17184 19780
rect 19984 19796 20036 19848
rect 20444 19839 20496 19848
rect 20444 19805 20453 19839
rect 20453 19805 20487 19839
rect 20487 19805 20496 19839
rect 20444 19796 20496 19805
rect 21180 19839 21232 19848
rect 21180 19805 21189 19839
rect 21189 19805 21223 19839
rect 21223 19805 21232 19839
rect 21180 19796 21232 19805
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 24400 19839 24452 19848
rect 24400 19805 24409 19839
rect 24409 19805 24443 19839
rect 24443 19805 24452 19839
rect 24400 19796 24452 19805
rect 27068 19796 27120 19848
rect 27252 19839 27304 19848
rect 27252 19805 27261 19839
rect 27261 19805 27295 19839
rect 27295 19805 27304 19839
rect 27252 19796 27304 19805
rect 27344 19796 27396 19848
rect 27620 19796 27672 19848
rect 14556 19660 14608 19712
rect 18052 19703 18104 19712
rect 18052 19669 18061 19703
rect 18061 19669 18095 19703
rect 18095 19669 18104 19703
rect 18052 19660 18104 19669
rect 22376 19728 22428 19780
rect 22652 19728 22704 19780
rect 26884 19728 26936 19780
rect 47676 19728 47728 19780
rect 48136 19771 48188 19780
rect 48136 19737 48145 19771
rect 48145 19737 48179 19771
rect 48179 19737 48188 19771
rect 48136 19728 48188 19737
rect 19248 19660 19300 19712
rect 19984 19660 20036 19712
rect 27436 19660 27488 19712
rect 46296 19660 46348 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 11612 19456 11664 19508
rect 3516 19388 3568 19440
rect 12072 19456 12124 19508
rect 22284 19499 22336 19508
rect 14740 19388 14792 19440
rect 17224 19388 17276 19440
rect 18788 19388 18840 19440
rect 22284 19465 22293 19499
rect 22293 19465 22327 19499
rect 22327 19465 22336 19499
rect 22284 19456 22336 19465
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 9680 19320 9732 19372
rect 9864 19363 9916 19372
rect 9864 19329 9873 19363
rect 9873 19329 9907 19363
rect 9907 19329 9916 19363
rect 9864 19320 9916 19329
rect 10600 19320 10652 19372
rect 10784 19363 10836 19372
rect 10784 19329 10793 19363
rect 10793 19329 10827 19363
rect 10827 19329 10836 19363
rect 10784 19320 10836 19329
rect 11980 19363 12032 19372
rect 11980 19329 11989 19363
rect 11989 19329 12023 19363
rect 12023 19329 12032 19363
rect 11980 19320 12032 19329
rect 12072 19320 12124 19372
rect 12440 19320 12492 19372
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 10324 19252 10376 19304
rect 13452 19227 13504 19236
rect 13452 19193 13461 19227
rect 13461 19193 13495 19227
rect 13495 19193 13504 19227
rect 13452 19184 13504 19193
rect 14280 19320 14332 19372
rect 17500 19363 17552 19372
rect 17500 19329 17509 19363
rect 17509 19329 17543 19363
rect 17543 19329 17552 19363
rect 17500 19320 17552 19329
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 26884 19456 26936 19508
rect 27252 19456 27304 19508
rect 45192 19388 45244 19440
rect 14004 19295 14056 19304
rect 14004 19261 14013 19295
rect 14013 19261 14047 19295
rect 14047 19261 14056 19295
rect 14004 19252 14056 19261
rect 17224 19252 17276 19304
rect 18420 19252 18472 19304
rect 22284 19252 22336 19304
rect 22560 19252 22612 19304
rect 13912 19184 13964 19236
rect 14556 19184 14608 19236
rect 16856 19184 16908 19236
rect 17316 19184 17368 19236
rect 27344 19320 27396 19372
rect 27528 19320 27580 19372
rect 45560 19363 45612 19372
rect 45560 19329 45569 19363
rect 45569 19329 45603 19363
rect 45603 19329 45612 19363
rect 45560 19320 45612 19329
rect 45744 19363 45796 19372
rect 45744 19329 45753 19363
rect 45753 19329 45787 19363
rect 45787 19329 45796 19363
rect 45744 19320 45796 19329
rect 23020 19295 23072 19304
rect 23020 19261 23029 19295
rect 23029 19261 23063 19295
rect 23063 19261 23072 19295
rect 23020 19252 23072 19261
rect 9312 19116 9364 19168
rect 11336 19116 11388 19168
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 12900 19116 12952 19125
rect 12992 19116 13044 19168
rect 19248 19159 19300 19168
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 20812 19116 20864 19168
rect 46112 19184 46164 19236
rect 46388 19320 46440 19372
rect 46388 19184 46440 19236
rect 22836 19116 22888 19168
rect 28172 19116 28224 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 3976 18912 4028 18964
rect 9312 18819 9364 18828
rect 9312 18785 9321 18819
rect 9321 18785 9355 18819
rect 9355 18785 9364 18819
rect 9312 18776 9364 18785
rect 9404 18776 9456 18828
rect 11336 18819 11388 18828
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 9036 18751 9088 18760
rect 2136 18708 2188 18717
rect 9036 18717 9045 18751
rect 9045 18717 9079 18751
rect 9079 18717 9088 18751
rect 9036 18708 9088 18717
rect 6644 18640 6696 18692
rect 9404 18640 9456 18692
rect 10324 18640 10376 18692
rect 9680 18572 9732 18624
rect 11336 18785 11345 18819
rect 11345 18785 11379 18819
rect 11379 18785 11388 18819
rect 11336 18776 11388 18785
rect 11612 18819 11664 18828
rect 11612 18785 11621 18819
rect 11621 18785 11655 18819
rect 11655 18785 11664 18819
rect 11612 18776 11664 18785
rect 12900 18776 12952 18828
rect 17132 18819 17184 18828
rect 17132 18785 17141 18819
rect 17141 18785 17175 18819
rect 17175 18785 17184 18819
rect 17132 18776 17184 18785
rect 18512 18912 18564 18964
rect 20536 18912 20588 18964
rect 21824 18912 21876 18964
rect 23020 18912 23072 18964
rect 24400 18955 24452 18964
rect 24400 18921 24409 18955
rect 24409 18921 24443 18955
rect 24443 18921 24452 18955
rect 24400 18912 24452 18921
rect 27252 18912 27304 18964
rect 18052 18844 18104 18896
rect 16672 18751 16724 18760
rect 16672 18717 16681 18751
rect 16681 18717 16715 18751
rect 16715 18717 16724 18751
rect 16672 18708 16724 18717
rect 17408 18708 17460 18760
rect 19340 18751 19392 18760
rect 19340 18717 19349 18751
rect 19349 18717 19383 18751
rect 19383 18717 19392 18751
rect 19340 18708 19392 18717
rect 19432 18708 19484 18760
rect 20536 18751 20588 18760
rect 20536 18717 20545 18751
rect 20545 18717 20579 18751
rect 20579 18717 20588 18751
rect 20536 18708 20588 18717
rect 22192 18708 22244 18760
rect 12072 18640 12124 18692
rect 13636 18640 13688 18692
rect 14832 18640 14884 18692
rect 16580 18640 16632 18692
rect 17224 18640 17276 18692
rect 12992 18572 13044 18624
rect 13084 18615 13136 18624
rect 13084 18581 13093 18615
rect 13093 18581 13127 18615
rect 13127 18581 13136 18615
rect 13084 18572 13136 18581
rect 13452 18572 13504 18624
rect 18420 18640 18472 18692
rect 20076 18640 20128 18692
rect 22652 18640 22704 18692
rect 47400 18844 47452 18896
rect 24400 18751 24452 18760
rect 24400 18717 24409 18751
rect 24409 18717 24443 18751
rect 24443 18717 24452 18751
rect 24400 18708 24452 18717
rect 24860 18640 24912 18692
rect 25596 18776 25648 18828
rect 26884 18776 26936 18828
rect 47308 18776 47360 18828
rect 26976 18708 27028 18760
rect 28172 18751 28224 18760
rect 27344 18683 27396 18692
rect 27344 18649 27353 18683
rect 27353 18649 27387 18683
rect 27387 18649 27396 18683
rect 28172 18717 28181 18751
rect 28181 18717 28215 18751
rect 28215 18717 28224 18751
rect 28172 18708 28224 18717
rect 45744 18708 45796 18760
rect 46296 18751 46348 18760
rect 46296 18717 46305 18751
rect 46305 18717 46339 18751
rect 46339 18717 46348 18751
rect 46296 18708 46348 18717
rect 27344 18640 27396 18649
rect 17500 18615 17552 18624
rect 17500 18581 17509 18615
rect 17509 18581 17543 18615
rect 17543 18581 17552 18615
rect 17500 18572 17552 18581
rect 24216 18572 24268 18624
rect 26240 18572 26292 18624
rect 27528 18615 27580 18624
rect 27528 18581 27553 18615
rect 27553 18581 27580 18615
rect 27528 18572 27580 18581
rect 28264 18615 28316 18624
rect 28264 18581 28273 18615
rect 28273 18581 28307 18615
rect 28307 18581 28316 18615
rect 28264 18572 28316 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 9036 18368 9088 18420
rect 10324 18368 10376 18420
rect 12072 18368 12124 18420
rect 14832 18368 14884 18420
rect 16672 18368 16724 18420
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 9864 18232 9916 18284
rect 11704 18232 11756 18284
rect 13452 18232 13504 18284
rect 14464 18232 14516 18284
rect 14832 18232 14884 18284
rect 16396 18300 16448 18352
rect 17500 18300 17552 18352
rect 19432 18368 19484 18420
rect 20076 18411 20128 18420
rect 20076 18377 20085 18411
rect 20085 18377 20119 18411
rect 20119 18377 20128 18411
rect 20076 18368 20128 18377
rect 20536 18368 20588 18420
rect 22652 18411 22704 18420
rect 22652 18377 22661 18411
rect 22661 18377 22695 18411
rect 22695 18377 22704 18411
rect 22652 18368 22704 18377
rect 22928 18300 22980 18352
rect 24216 18343 24268 18352
rect 24216 18309 24225 18343
rect 24225 18309 24259 18343
rect 24259 18309 24268 18343
rect 24216 18300 24268 18309
rect 28264 18368 28316 18420
rect 47676 18411 47728 18420
rect 47676 18377 47685 18411
rect 47685 18377 47719 18411
rect 47719 18377 47728 18411
rect 47676 18368 47728 18377
rect 27988 18300 28040 18352
rect 13360 18207 13412 18216
rect 13360 18173 13369 18207
rect 13369 18173 13403 18207
rect 13403 18173 13412 18207
rect 13360 18164 13412 18173
rect 13636 18207 13688 18216
rect 13636 18173 13645 18207
rect 13645 18173 13679 18207
rect 13679 18173 13688 18207
rect 13636 18164 13688 18173
rect 16856 18232 16908 18284
rect 16948 18275 17000 18284
rect 16948 18241 16957 18275
rect 16957 18241 16991 18275
rect 16991 18241 17000 18275
rect 16948 18232 17000 18241
rect 18420 18232 18472 18284
rect 18512 18232 18564 18284
rect 20260 18232 20312 18284
rect 23204 18275 23256 18284
rect 23204 18241 23213 18275
rect 23213 18241 23247 18275
rect 23247 18241 23256 18275
rect 23204 18232 23256 18241
rect 46388 18275 46440 18284
rect 46388 18241 46397 18275
rect 46397 18241 46431 18275
rect 46431 18241 46440 18275
rect 46388 18232 46440 18241
rect 47032 18275 47084 18284
rect 47032 18241 47041 18275
rect 47041 18241 47075 18275
rect 47075 18241 47084 18275
rect 47032 18232 47084 18241
rect 47584 18275 47636 18284
rect 47584 18241 47593 18275
rect 47593 18241 47627 18275
rect 47627 18241 47636 18275
rect 47584 18232 47636 18241
rect 15660 18164 15712 18216
rect 19340 18164 19392 18216
rect 24584 18164 24636 18216
rect 24860 18207 24912 18216
rect 24860 18173 24869 18207
rect 24869 18173 24903 18207
rect 24903 18173 24912 18207
rect 24860 18164 24912 18173
rect 26976 18207 27028 18216
rect 26976 18173 26985 18207
rect 26985 18173 27019 18207
rect 27019 18173 27028 18207
rect 26976 18164 27028 18173
rect 16672 18139 16724 18148
rect 14280 18028 14332 18080
rect 16672 18105 16681 18139
rect 16681 18105 16715 18139
rect 16715 18105 16724 18139
rect 16672 18096 16724 18105
rect 17132 18096 17184 18148
rect 17500 18028 17552 18080
rect 20720 18071 20772 18080
rect 20720 18037 20729 18071
rect 20729 18037 20763 18071
rect 20763 18037 20772 18071
rect 20720 18028 20772 18037
rect 22744 18028 22796 18080
rect 27344 18028 27396 18080
rect 29092 18028 29144 18080
rect 46204 18071 46256 18080
rect 46204 18037 46213 18071
rect 46213 18037 46247 18071
rect 46247 18037 46256 18071
rect 46204 18028 46256 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 14004 17824 14056 17876
rect 17316 17824 17368 17876
rect 19340 17867 19392 17876
rect 19340 17833 19349 17867
rect 19349 17833 19383 17867
rect 19383 17833 19392 17867
rect 19340 17824 19392 17833
rect 19984 17824 20036 17876
rect 24400 17824 24452 17876
rect 26884 17824 26936 17876
rect 27988 17824 28040 17876
rect 12440 17663 12492 17672
rect 12440 17629 12449 17663
rect 12449 17629 12483 17663
rect 12483 17629 12492 17663
rect 12440 17620 12492 17629
rect 13360 17620 13412 17672
rect 16948 17756 17000 17808
rect 16672 17688 16724 17740
rect 16212 17620 16264 17672
rect 18420 17688 18472 17740
rect 13820 17552 13872 17604
rect 12716 17484 12768 17536
rect 12992 17484 13044 17536
rect 14280 17595 14332 17604
rect 14280 17561 14305 17595
rect 14305 17561 14332 17595
rect 14280 17552 14332 17561
rect 14740 17484 14792 17536
rect 16580 17484 16632 17536
rect 16948 17620 17000 17672
rect 16856 17552 16908 17604
rect 18512 17620 18564 17672
rect 20720 17688 20772 17740
rect 25596 17688 25648 17740
rect 25228 17663 25280 17672
rect 25228 17629 25237 17663
rect 25237 17629 25271 17663
rect 25271 17629 25280 17663
rect 25228 17620 25280 17629
rect 20260 17552 20312 17604
rect 20812 17552 20864 17604
rect 22744 17552 22796 17604
rect 22928 17595 22980 17604
rect 22928 17561 22937 17595
rect 22937 17561 22971 17595
rect 22971 17561 22980 17595
rect 22928 17552 22980 17561
rect 26240 17552 26292 17604
rect 17500 17484 17552 17536
rect 18144 17484 18196 17536
rect 46020 17688 46072 17740
rect 27068 17620 27120 17672
rect 29644 17595 29696 17604
rect 29644 17561 29653 17595
rect 29653 17561 29687 17595
rect 29687 17561 29696 17595
rect 29644 17552 29696 17561
rect 30012 17552 30064 17604
rect 30656 17595 30708 17604
rect 30656 17561 30665 17595
rect 30665 17561 30699 17595
rect 30699 17561 30708 17595
rect 30656 17552 30708 17561
rect 47676 17552 47728 17604
rect 48136 17595 48188 17604
rect 48136 17561 48145 17595
rect 48145 17561 48179 17595
rect 48179 17561 48188 17595
rect 48136 17552 48188 17561
rect 40224 17484 40276 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4988 17280 5040 17332
rect 12992 17255 13044 17264
rect 12992 17221 13001 17255
rect 13001 17221 13035 17255
rect 13035 17221 13044 17255
rect 12992 17212 13044 17221
rect 19432 17212 19484 17264
rect 25228 17280 25280 17332
rect 26976 17280 27028 17332
rect 47676 17323 47728 17332
rect 47676 17289 47685 17323
rect 47685 17289 47719 17323
rect 47719 17289 47728 17323
rect 47676 17280 47728 17289
rect 23664 17255 23716 17264
rect 23664 17221 23673 17255
rect 23673 17221 23707 17255
rect 23707 17221 23716 17255
rect 23664 17212 23716 17221
rect 24400 17212 24452 17264
rect 12716 17187 12768 17196
rect 12716 17153 12725 17187
rect 12725 17153 12759 17187
rect 12759 17153 12768 17187
rect 12716 17144 12768 17153
rect 14832 17144 14884 17196
rect 15844 17187 15896 17196
rect 15844 17153 15853 17187
rect 15853 17153 15887 17187
rect 15887 17153 15896 17187
rect 15844 17144 15896 17153
rect 17316 17187 17368 17196
rect 17316 17153 17325 17187
rect 17325 17153 17359 17187
rect 17359 17153 17368 17187
rect 17316 17144 17368 17153
rect 18144 17187 18196 17196
rect 18144 17153 18153 17187
rect 18153 17153 18187 17187
rect 18187 17153 18196 17187
rect 18144 17144 18196 17153
rect 45100 17212 45152 17264
rect 47124 17212 47176 17264
rect 28448 17187 28500 17196
rect 3332 17076 3384 17128
rect 7932 17076 7984 17128
rect 14740 17119 14792 17128
rect 14740 17085 14749 17119
rect 14749 17085 14783 17119
rect 14783 17085 14792 17119
rect 14740 17076 14792 17085
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 1400 16940 1452 16992
rect 10692 16940 10744 16992
rect 16672 17008 16724 17060
rect 28448 17153 28457 17187
rect 28457 17153 28491 17187
rect 28491 17153 28500 17187
rect 28448 17144 28500 17153
rect 29092 17187 29144 17196
rect 29092 17153 29101 17187
rect 29101 17153 29135 17187
rect 29135 17153 29144 17187
rect 29092 17144 29144 17153
rect 46848 17144 46900 17196
rect 47400 17144 47452 17196
rect 23756 17076 23808 17128
rect 30932 17119 30984 17128
rect 30932 17085 30941 17119
rect 30941 17085 30975 17119
rect 30975 17085 30984 17119
rect 30932 17076 30984 17085
rect 45192 17119 45244 17128
rect 45192 17085 45201 17119
rect 45201 17085 45235 17119
rect 45235 17085 45244 17119
rect 45192 17076 45244 17085
rect 23480 17008 23532 17060
rect 30656 17008 30708 17060
rect 15844 16940 15896 16992
rect 17316 16940 17368 16992
rect 24860 16940 24912 16992
rect 39764 16940 39816 16992
rect 45468 16940 45520 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 13820 16736 13872 16788
rect 20996 16736 21048 16788
rect 29644 16736 29696 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 2320 16600 2372 16652
rect 14740 16668 14792 16720
rect 3424 16600 3476 16652
rect 13084 16600 13136 16652
rect 15844 16643 15896 16652
rect 15844 16609 15853 16643
rect 15853 16609 15887 16643
rect 15887 16609 15896 16643
rect 15844 16600 15896 16609
rect 20996 16643 21048 16652
rect 20996 16609 21005 16643
rect 21005 16609 21039 16643
rect 21039 16609 21048 16643
rect 20996 16600 21048 16609
rect 24492 16600 24544 16652
rect 25412 16600 25464 16652
rect 39764 16600 39816 16652
rect 45928 16736 45980 16788
rect 40224 16643 40276 16652
rect 40224 16609 40233 16643
rect 40233 16609 40267 16643
rect 40267 16609 40276 16643
rect 40224 16600 40276 16609
rect 47032 16600 47084 16652
rect 10692 16575 10744 16584
rect 10692 16541 10701 16575
rect 10701 16541 10735 16575
rect 10735 16541 10744 16575
rect 10692 16532 10744 16541
rect 14280 16532 14332 16584
rect 2136 16464 2188 16516
rect 10876 16507 10928 16516
rect 10876 16473 10885 16507
rect 10885 16473 10919 16507
rect 10919 16473 10928 16507
rect 10876 16464 10928 16473
rect 14740 16464 14792 16516
rect 15844 16464 15896 16516
rect 19340 16532 19392 16584
rect 19984 16532 20036 16584
rect 23480 16532 23532 16584
rect 23664 16575 23716 16584
rect 23664 16541 23673 16575
rect 23673 16541 23707 16575
rect 23707 16541 23716 16575
rect 23664 16532 23716 16541
rect 24860 16575 24912 16584
rect 24860 16541 24869 16575
rect 24869 16541 24903 16575
rect 24903 16541 24912 16575
rect 24860 16532 24912 16541
rect 45652 16532 45704 16584
rect 46020 16532 46072 16584
rect 17500 16507 17552 16516
rect 17500 16473 17509 16507
rect 17509 16473 17543 16507
rect 17543 16473 17552 16507
rect 17500 16464 17552 16473
rect 22008 16507 22060 16516
rect 14004 16396 14056 16448
rect 15108 16396 15160 16448
rect 19340 16396 19392 16448
rect 20168 16396 20220 16448
rect 22008 16473 22017 16507
rect 22017 16473 22051 16507
rect 22051 16473 22060 16507
rect 22008 16464 22060 16473
rect 23756 16507 23808 16516
rect 23756 16473 23765 16507
rect 23765 16473 23799 16507
rect 23799 16473 23808 16507
rect 23756 16464 23808 16473
rect 30196 16507 30248 16516
rect 30196 16473 30205 16507
rect 30205 16473 30239 16507
rect 30239 16473 30248 16507
rect 30196 16464 30248 16473
rect 40408 16464 40460 16516
rect 47676 16464 47728 16516
rect 48136 16507 48188 16516
rect 48136 16473 48145 16507
rect 48145 16473 48179 16507
rect 48179 16473 48188 16507
rect 48136 16464 48188 16473
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 10876 16235 10928 16244
rect 10876 16201 10885 16235
rect 10885 16201 10919 16235
rect 10919 16201 10928 16235
rect 10876 16192 10928 16201
rect 16580 16192 16632 16244
rect 17316 16192 17368 16244
rect 19432 16192 19484 16244
rect 30196 16235 30248 16244
rect 30196 16201 30205 16235
rect 30205 16201 30239 16235
rect 30239 16201 30248 16235
rect 30196 16192 30248 16201
rect 1952 16056 2004 16108
rect 15844 16124 15896 16176
rect 16212 16124 16264 16176
rect 18052 16124 18104 16176
rect 24584 16124 24636 16176
rect 11060 16056 11112 16108
rect 16672 16056 16724 16108
rect 16856 16056 16908 16108
rect 17408 16056 17460 16108
rect 18604 16056 18656 16108
rect 19248 16056 19300 16108
rect 23756 16099 23808 16108
rect 23756 16065 23765 16099
rect 23765 16065 23799 16099
rect 23799 16065 23808 16099
rect 23756 16056 23808 16065
rect 24400 16099 24452 16108
rect 24400 16065 24409 16099
rect 24409 16065 24443 16099
rect 24443 16065 24452 16099
rect 24400 16056 24452 16065
rect 30104 16099 30156 16108
rect 30104 16065 30113 16099
rect 30113 16065 30147 16099
rect 30147 16065 30156 16099
rect 46480 16192 46532 16244
rect 47676 16235 47728 16244
rect 47676 16201 47685 16235
rect 47685 16201 47719 16235
rect 47719 16201 47728 16235
rect 47676 16192 47728 16201
rect 46664 16124 46716 16176
rect 46940 16124 46992 16176
rect 47032 16099 47084 16108
rect 30104 16056 30156 16065
rect 47032 16065 47041 16099
rect 47041 16065 47075 16099
rect 47075 16065 47084 16099
rect 47032 16056 47084 16065
rect 17224 15852 17276 15904
rect 18328 15852 18380 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 18972 15648 19024 15700
rect 2044 15580 2096 15632
rect 22008 15648 22060 15700
rect 23940 15648 23992 15700
rect 24400 15648 24452 15700
rect 9220 15512 9272 15564
rect 13360 15555 13412 15564
rect 1768 15444 1820 15496
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13360 15512 13412 15521
rect 14280 15512 14332 15564
rect 15016 15512 15068 15564
rect 16212 15512 16264 15564
rect 27068 15580 27120 15632
rect 23480 15512 23532 15564
rect 23756 15512 23808 15564
rect 9864 15419 9916 15428
rect 9864 15385 9873 15419
rect 9873 15385 9907 15419
rect 9907 15385 9916 15419
rect 9864 15376 9916 15385
rect 13636 15444 13688 15496
rect 14832 15487 14884 15496
rect 14004 15376 14056 15428
rect 14832 15453 14841 15487
rect 14841 15453 14875 15487
rect 14875 15453 14884 15487
rect 14832 15444 14884 15453
rect 16120 15419 16172 15428
rect 13820 15308 13872 15360
rect 14924 15351 14976 15360
rect 14924 15317 14933 15351
rect 14933 15317 14967 15351
rect 14967 15317 14976 15351
rect 14924 15308 14976 15317
rect 16120 15385 16129 15419
rect 16129 15385 16163 15419
rect 16163 15385 16172 15419
rect 16120 15376 16172 15385
rect 19340 15444 19392 15496
rect 19984 15444 20036 15496
rect 17776 15419 17828 15428
rect 17776 15385 17785 15419
rect 17785 15385 17819 15419
rect 17819 15385 17828 15419
rect 17776 15376 17828 15385
rect 17960 15308 18012 15360
rect 22100 15444 22152 15496
rect 23664 15444 23716 15496
rect 46388 15487 46440 15496
rect 23848 15376 23900 15428
rect 46388 15453 46397 15487
rect 46397 15453 46431 15487
rect 46431 15453 46440 15487
rect 46388 15444 46440 15453
rect 47860 15487 47912 15496
rect 47860 15453 47869 15487
rect 47869 15453 47903 15487
rect 47903 15453 47912 15487
rect 47860 15444 47912 15453
rect 24860 15376 24912 15428
rect 45192 15376 45244 15428
rect 23388 15351 23440 15360
rect 23388 15317 23397 15351
rect 23397 15317 23431 15351
rect 23431 15317 23440 15351
rect 23388 15308 23440 15317
rect 47860 15308 47912 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 9864 15104 9916 15156
rect 16120 15104 16172 15156
rect 13360 15036 13412 15088
rect 14924 15036 14976 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 11060 14968 11112 15020
rect 15936 15011 15988 15020
rect 15936 14977 15945 15011
rect 15945 14977 15979 15011
rect 15979 14977 15988 15011
rect 15936 14968 15988 14977
rect 17960 15104 18012 15156
rect 18052 15104 18104 15156
rect 23756 15147 23808 15156
rect 17224 15079 17276 15088
rect 17224 15045 17233 15079
rect 17233 15045 17267 15079
rect 17267 15045 17276 15079
rect 17224 15036 17276 15045
rect 23756 15113 23765 15147
rect 23765 15113 23799 15147
rect 23799 15113 23808 15147
rect 23756 15104 23808 15113
rect 24492 15104 24544 15156
rect 24860 15147 24912 15156
rect 24860 15113 24869 15147
rect 24869 15113 24903 15147
rect 24903 15113 24912 15147
rect 24860 15104 24912 15113
rect 18328 14968 18380 15020
rect 20352 14968 20404 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 22100 14968 22152 15020
rect 23388 15036 23440 15088
rect 23940 15036 23992 15088
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 13820 14900 13872 14952
rect 15108 14900 15160 14952
rect 20260 14900 20312 14952
rect 23756 14968 23808 15020
rect 25964 15036 26016 15088
rect 26148 15036 26200 15088
rect 20720 14764 20772 14816
rect 21180 14807 21232 14816
rect 21180 14773 21189 14807
rect 21189 14773 21223 14807
rect 21223 14773 21232 14807
rect 21180 14764 21232 14773
rect 23020 14807 23072 14816
rect 23020 14773 23029 14807
rect 23029 14773 23063 14807
rect 23063 14773 23072 14807
rect 23020 14764 23072 14773
rect 46204 15036 46256 15088
rect 47768 15079 47820 15088
rect 47768 15045 47777 15079
rect 47777 15045 47811 15079
rect 47811 15045 47820 15079
rect 47768 15036 47820 15045
rect 45192 15011 45244 15020
rect 45192 14977 45201 15011
rect 45201 14977 45235 15011
rect 45235 14977 45244 15011
rect 45192 14968 45244 14977
rect 47676 14968 47728 15020
rect 45652 14900 45704 14952
rect 46388 14764 46440 14816
rect 46848 14764 46900 14816
rect 47952 14807 48004 14816
rect 47952 14773 47961 14807
rect 47961 14773 47995 14807
rect 47995 14773 48004 14807
rect 47952 14764 48004 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 16396 14603 16448 14612
rect 16396 14569 16405 14603
rect 16405 14569 16439 14603
rect 16439 14569 16448 14603
rect 16396 14560 16448 14569
rect 17132 14560 17184 14612
rect 16856 14492 16908 14544
rect 22928 14560 22980 14612
rect 24492 14603 24544 14612
rect 24492 14569 24501 14603
rect 24501 14569 24535 14603
rect 24535 14569 24544 14603
rect 24492 14560 24544 14569
rect 45652 14603 45704 14612
rect 45652 14569 45661 14603
rect 45661 14569 45695 14603
rect 45695 14569 45704 14603
rect 45652 14560 45704 14569
rect 3884 14424 3936 14476
rect 17408 14492 17460 14544
rect 26148 14492 26200 14544
rect 46572 14492 46624 14544
rect 17224 14424 17276 14476
rect 21824 14467 21876 14476
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 14832 14356 14884 14408
rect 15016 14356 15068 14408
rect 15384 14399 15436 14408
rect 14464 14288 14516 14340
rect 15384 14365 15393 14399
rect 15393 14365 15427 14399
rect 15427 14365 15436 14399
rect 15384 14356 15436 14365
rect 16856 14331 16908 14340
rect 14280 14220 14332 14272
rect 15384 14220 15436 14272
rect 16856 14297 16865 14331
rect 16865 14297 16899 14331
rect 16899 14297 16908 14331
rect 16856 14288 16908 14297
rect 19248 14356 19300 14408
rect 20260 14399 20312 14408
rect 20260 14365 20269 14399
rect 20269 14365 20303 14399
rect 20303 14365 20312 14399
rect 20260 14356 20312 14365
rect 16948 14220 17000 14272
rect 17040 14263 17092 14272
rect 21824 14433 21833 14467
rect 21833 14433 21867 14467
rect 21867 14433 21876 14467
rect 21824 14424 21876 14433
rect 22928 14424 22980 14476
rect 23020 14399 23072 14408
rect 23020 14365 23029 14399
rect 23029 14365 23063 14399
rect 23063 14365 23072 14399
rect 23020 14356 23072 14365
rect 46664 14467 46716 14476
rect 46664 14433 46673 14467
rect 46673 14433 46707 14467
rect 46707 14433 46716 14467
rect 46664 14424 46716 14433
rect 47768 14492 47820 14544
rect 25228 14399 25280 14408
rect 17040 14229 17065 14263
rect 17065 14229 17092 14263
rect 17040 14220 17092 14229
rect 19432 14263 19484 14272
rect 19432 14229 19441 14263
rect 19441 14229 19475 14263
rect 19475 14229 19484 14263
rect 19432 14220 19484 14229
rect 22284 14288 22336 14340
rect 23756 14288 23808 14340
rect 21180 14220 21232 14272
rect 23848 14263 23900 14272
rect 23848 14229 23857 14263
rect 23857 14229 23891 14263
rect 23891 14229 23900 14263
rect 23848 14220 23900 14229
rect 24032 14288 24084 14340
rect 25228 14365 25237 14399
rect 25237 14365 25271 14399
rect 25271 14365 25280 14399
rect 25228 14356 25280 14365
rect 46296 14356 46348 14408
rect 47676 14356 47728 14408
rect 47216 14288 47268 14340
rect 48228 14288 48280 14340
rect 47860 14263 47912 14272
rect 47860 14229 47869 14263
rect 47869 14229 47903 14263
rect 47903 14229 47912 14263
rect 47860 14220 47912 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 2136 14016 2188 14068
rect 17224 14016 17276 14068
rect 14280 13948 14332 14000
rect 14464 13948 14516 14000
rect 16856 13948 16908 14000
rect 17960 13948 18012 14000
rect 13636 13880 13688 13932
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 16672 13880 16724 13932
rect 16948 13923 17000 13932
rect 16948 13889 16957 13923
rect 16957 13889 16991 13923
rect 16991 13889 17000 13923
rect 19340 14016 19392 14068
rect 23756 14059 23808 14068
rect 23756 14025 23765 14059
rect 23765 14025 23799 14059
rect 23799 14025 23808 14059
rect 23756 14016 23808 14025
rect 25228 14016 25280 14068
rect 47952 14016 48004 14068
rect 19432 13948 19484 14000
rect 46480 13948 46532 14000
rect 16948 13880 17000 13889
rect 15476 13855 15528 13864
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17040 13812 17092 13864
rect 3976 13676 4028 13728
rect 13820 13676 13872 13728
rect 16028 13719 16080 13728
rect 16028 13685 16037 13719
rect 16037 13685 16071 13719
rect 16071 13685 16080 13719
rect 16028 13676 16080 13685
rect 22928 13880 22980 13932
rect 24032 13880 24084 13932
rect 24492 13880 24544 13932
rect 46296 13880 46348 13932
rect 47216 13880 47268 13932
rect 22284 13812 22336 13864
rect 22836 13812 22888 13864
rect 46848 13855 46900 13864
rect 46848 13821 46857 13855
rect 46857 13821 46891 13855
rect 46891 13821 46900 13855
rect 46848 13812 46900 13821
rect 47860 13812 47912 13864
rect 20168 13719 20220 13728
rect 20168 13685 20177 13719
rect 20177 13685 20211 13719
rect 20211 13685 20220 13719
rect 20168 13676 20220 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19340 13472 19392 13524
rect 46664 13515 46716 13524
rect 46664 13481 46673 13515
rect 46673 13481 46707 13515
rect 46707 13481 46716 13515
rect 46664 13472 46716 13481
rect 12440 13404 12492 13456
rect 16028 13336 16080 13388
rect 19248 13404 19300 13456
rect 20168 13336 20220 13388
rect 20720 13379 20772 13388
rect 20720 13345 20729 13379
rect 20729 13345 20763 13379
rect 20763 13345 20772 13379
rect 20720 13336 20772 13345
rect 45376 13336 45428 13388
rect 47216 13336 47268 13388
rect 15476 13200 15528 13252
rect 19984 13268 20036 13320
rect 30472 13200 30524 13252
rect 45192 13200 45244 13252
rect 46112 13268 46164 13320
rect 47676 13311 47728 13320
rect 47676 13277 47685 13311
rect 47685 13277 47719 13311
rect 47719 13277 47728 13311
rect 47676 13268 47728 13277
rect 17132 13132 17184 13184
rect 18512 13175 18564 13184
rect 18512 13141 18521 13175
rect 18521 13141 18555 13175
rect 18555 13141 18564 13175
rect 18512 13132 18564 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 18512 12792 18564 12844
rect 21548 12792 21600 12844
rect 21732 12792 21784 12844
rect 23848 12792 23900 12844
rect 45192 12835 45244 12844
rect 45192 12801 45201 12835
rect 45201 12801 45235 12835
rect 45235 12801 45244 12835
rect 45192 12792 45244 12801
rect 45376 12835 45428 12844
rect 45376 12801 45385 12835
rect 45385 12801 45419 12835
rect 45419 12801 45428 12835
rect 45376 12792 45428 12801
rect 46112 12792 46164 12844
rect 46296 12835 46348 12844
rect 46296 12801 46305 12835
rect 46305 12801 46339 12835
rect 46339 12801 46348 12835
rect 46296 12792 46348 12801
rect 17040 12724 17092 12776
rect 25872 12767 25924 12776
rect 25872 12733 25881 12767
rect 25881 12733 25915 12767
rect 25915 12733 25924 12767
rect 25872 12724 25924 12733
rect 47216 12792 47268 12844
rect 25044 12656 25096 12708
rect 18880 12631 18932 12640
rect 18880 12597 18889 12631
rect 18889 12597 18923 12631
rect 18923 12597 18932 12631
rect 18880 12588 18932 12597
rect 45836 12631 45888 12640
rect 45836 12597 45845 12631
rect 45845 12597 45879 12631
rect 45879 12597 45888 12631
rect 45836 12588 45888 12597
rect 46020 12588 46072 12640
rect 46204 12588 46256 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 45744 12384 45796 12436
rect 17040 12359 17092 12368
rect 17040 12325 17049 12359
rect 17049 12325 17083 12359
rect 17083 12325 17092 12359
rect 17040 12316 17092 12325
rect 16856 12248 16908 12300
rect 45744 12291 45796 12300
rect 45744 12257 45753 12291
rect 45753 12257 45787 12291
rect 45787 12257 45796 12291
rect 45744 12248 45796 12257
rect 47676 12316 47728 12368
rect 46480 12291 46532 12300
rect 46480 12257 46489 12291
rect 46489 12257 46523 12291
rect 46523 12257 46532 12291
rect 46480 12248 46532 12257
rect 48136 12291 48188 12300
rect 48136 12257 48145 12291
rect 48145 12257 48179 12291
rect 48179 12257 48188 12291
rect 48136 12248 48188 12257
rect 15016 12180 15068 12232
rect 17960 12180 18012 12232
rect 18880 12180 18932 12232
rect 45652 12180 45704 12232
rect 45376 12112 45428 12164
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 15660 11704 15712 11756
rect 21364 11704 21416 11756
rect 45744 11747 45796 11756
rect 45744 11713 45753 11747
rect 45753 11713 45787 11747
rect 45787 11713 45796 11747
rect 45744 11704 45796 11713
rect 45836 11704 45888 11756
rect 45560 11568 45612 11620
rect 46756 11568 46808 11620
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 15200 11500 15252 11509
rect 47768 11543 47820 11552
rect 47768 11509 47777 11543
rect 47777 11509 47811 11543
rect 47811 11509 47820 11543
rect 47768 11500 47820 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3332 11296 3384 11348
rect 14832 11296 14884 11348
rect 15016 11203 15068 11212
rect 15016 11169 15025 11203
rect 15025 11169 15059 11203
rect 15059 11169 15068 11203
rect 15016 11160 15068 11169
rect 15200 11203 15252 11212
rect 15200 11169 15209 11203
rect 15209 11169 15243 11203
rect 15243 11169 15252 11203
rect 15200 11160 15252 11169
rect 21732 11296 21784 11348
rect 45560 11296 45612 11348
rect 45836 11339 45888 11348
rect 45836 11305 45845 11339
rect 45845 11305 45879 11339
rect 45879 11305 45888 11339
rect 45836 11296 45888 11305
rect 45652 11271 45704 11280
rect 45652 11237 45661 11271
rect 45661 11237 45695 11271
rect 45695 11237 45704 11271
rect 45652 11228 45704 11237
rect 45376 11203 45428 11212
rect 45376 11169 45385 11203
rect 45385 11169 45419 11203
rect 45419 11169 45428 11203
rect 45376 11160 45428 11169
rect 47768 11160 47820 11212
rect 21732 11135 21784 11144
rect 21732 11101 21741 11135
rect 21741 11101 21775 11135
rect 21775 11101 21784 11135
rect 21732 11092 21784 11101
rect 21916 11067 21968 11076
rect 21916 11033 21925 11067
rect 21925 11033 21959 11067
rect 21959 11033 21968 11067
rect 21916 11024 21968 11033
rect 46020 11024 46072 11076
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 21916 10795 21968 10804
rect 21916 10761 21925 10795
rect 21925 10761 21959 10795
rect 21959 10761 21968 10795
rect 21916 10752 21968 10761
rect 45376 10795 45428 10804
rect 45376 10761 45385 10795
rect 45385 10761 45419 10795
rect 45419 10761 45428 10795
rect 45376 10752 45428 10761
rect 46112 10727 46164 10736
rect 46112 10693 46121 10727
rect 46121 10693 46155 10727
rect 46155 10693 46164 10727
rect 46112 10684 46164 10693
rect 21640 10616 21692 10668
rect 45468 10659 45520 10668
rect 45468 10625 45477 10659
rect 45477 10625 45511 10659
rect 45511 10625 45520 10659
rect 45468 10616 45520 10625
rect 45376 10548 45428 10600
rect 46204 10548 46256 10600
rect 45560 10480 45612 10532
rect 3516 10412 3568 10464
rect 9220 10412 9272 10464
rect 46296 10412 46348 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 45652 10251 45704 10260
rect 45652 10217 45661 10251
rect 45661 10217 45695 10251
rect 45695 10217 45704 10251
rect 45652 10208 45704 10217
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 45560 10047 45612 10056
rect 45560 10013 45569 10047
rect 45569 10013 45603 10047
rect 45603 10013 45612 10047
rect 45560 10004 45612 10013
rect 45100 9936 45152 9988
rect 45468 9936 45520 9988
rect 47676 9936 47728 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 46112 9664 46164 9716
rect 47676 9639 47728 9648
rect 47676 9605 47685 9639
rect 47685 9605 47719 9639
rect 47719 9605 47728 9639
rect 47676 9596 47728 9605
rect 46848 9528 46900 9580
rect 47492 9528 47544 9580
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 16580 8984 16632 9036
rect 16672 8984 16724 9036
rect 15660 8959 15712 8968
rect 15660 8925 15669 8959
rect 15669 8925 15703 8959
rect 15703 8925 15712 8959
rect 15660 8916 15712 8925
rect 47308 8959 47360 8968
rect 47308 8925 47317 8959
rect 47317 8925 47351 8959
rect 47351 8925 47360 8959
rect 47308 8916 47360 8925
rect 47400 8916 47452 8968
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 47768 8551 47820 8560
rect 47768 8517 47777 8551
rect 47777 8517 47811 8551
rect 47811 8517 47820 8551
rect 47768 8508 47820 8517
rect 24952 8304 25004 8356
rect 2964 8236 3016 8288
rect 12440 8236 12492 8288
rect 21824 8236 21876 8288
rect 45560 8236 45612 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 30932 7964 30984 8016
rect 33876 7964 33928 8016
rect 47124 7964 47176 8016
rect 47400 7896 47452 7948
rect 47676 7939 47728 7948
rect 47676 7905 47685 7939
rect 47685 7905 47719 7939
rect 47719 7905 47728 7939
rect 47676 7896 47728 7905
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 48136 7395 48188 7404
rect 48136 7361 48145 7395
rect 48145 7361 48179 7395
rect 48179 7361 48188 7395
rect 48136 7352 48188 7361
rect 47124 7148 47176 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3516 6808 3568 6860
rect 17776 6808 17828 6860
rect 47124 6851 47176 6860
rect 47124 6817 47133 6851
rect 47133 6817 47167 6851
rect 47167 6817 47176 6851
rect 47124 6808 47176 6817
rect 48228 6808 48280 6860
rect 22376 6740 22428 6792
rect 1676 6672 1728 6724
rect 6920 6604 6972 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 6920 6375 6972 6384
rect 6920 6341 6929 6375
rect 6929 6341 6963 6375
rect 6963 6341 6972 6375
rect 6920 6332 6972 6341
rect 6920 6196 6972 6248
rect 6460 6128 6512 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 46848 5720 46900 5772
rect 21088 5652 21140 5704
rect 47216 5652 47268 5704
rect 20628 5516 20680 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 18880 5176 18932 5185
rect 20812 5176 20864 5228
rect 22376 5176 22428 5228
rect 22744 5176 22796 5228
rect 23480 5219 23532 5228
rect 23480 5185 23489 5219
rect 23489 5185 23523 5219
rect 23523 5185 23532 5219
rect 23480 5176 23532 5185
rect 46848 5176 46900 5228
rect 48320 5176 48372 5228
rect 44732 5040 44784 5092
rect 18604 4972 18656 5024
rect 21364 4972 21416 5024
rect 22468 4972 22520 5024
rect 23204 4972 23256 5024
rect 24676 4972 24728 5024
rect 47216 4972 47268 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 20812 4811 20864 4820
rect 20812 4777 20821 4811
rect 20821 4777 20855 4811
rect 20855 4777 20864 4811
rect 20812 4768 20864 4777
rect 22744 4811 22796 4820
rect 22744 4777 22753 4811
rect 22753 4777 22787 4811
rect 22787 4777 22796 4811
rect 22744 4768 22796 4777
rect 46388 4768 46440 4820
rect 47584 4768 47636 4820
rect 24492 4632 24544 4684
rect 44732 4632 44784 4684
rect 45376 4632 45428 4684
rect 48228 4632 48280 4684
rect 10324 4564 10376 4616
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 18972 4564 19024 4616
rect 20076 4607 20128 4616
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 20720 4607 20772 4616
rect 20720 4573 20729 4607
rect 20729 4573 20763 4607
rect 20763 4573 20772 4607
rect 20720 4564 20772 4573
rect 21364 4607 21416 4616
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 22008 4607 22060 4616
rect 22008 4573 22017 4607
rect 22017 4573 22051 4607
rect 22051 4573 22060 4607
rect 22008 4564 22060 4573
rect 22468 4564 22520 4616
rect 23204 4564 23256 4616
rect 43812 4564 43864 4616
rect 46388 4607 46440 4616
rect 19340 4496 19392 4548
rect 27068 4539 27120 4548
rect 27068 4505 27077 4539
rect 27077 4505 27111 4539
rect 27111 4505 27120 4539
rect 27068 4496 27120 4505
rect 27252 4496 27304 4548
rect 39672 4496 39724 4548
rect 45192 4496 45244 4548
rect 46388 4573 46397 4607
rect 46397 4573 46431 4607
rect 46431 4573 46440 4607
rect 46388 4564 46440 4573
rect 18788 4428 18840 4480
rect 19432 4428 19484 4480
rect 21824 4428 21876 4480
rect 23204 4428 23256 4480
rect 23848 4428 23900 4480
rect 43720 4428 43772 4480
rect 45744 4471 45796 4480
rect 45744 4437 45753 4471
rect 45753 4437 45787 4471
rect 45787 4437 45796 4471
rect 45744 4428 45796 4437
rect 46480 4471 46532 4480
rect 46480 4437 46489 4471
rect 46489 4437 46523 4471
rect 46523 4437 46532 4471
rect 46480 4428 46532 4437
rect 47216 4539 47268 4548
rect 47216 4505 47225 4539
rect 47225 4505 47259 4539
rect 47259 4505 47268 4539
rect 47216 4496 47268 4505
rect 47032 4428 47084 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 18512 4224 18564 4276
rect 20076 4224 20128 4276
rect 40592 4267 40644 4276
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 3424 4020 3476 4072
rect 15660 4020 15712 4072
rect 16672 3952 16724 4004
rect 1676 3884 1728 3936
rect 2780 3884 2832 3936
rect 8116 3884 8168 3936
rect 9128 3884 9180 3936
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 17684 4088 17736 4140
rect 18512 4088 18564 4140
rect 18972 4088 19024 4140
rect 19432 4131 19484 4140
rect 19432 4097 19441 4131
rect 19441 4097 19475 4131
rect 19475 4097 19484 4131
rect 19432 4088 19484 4097
rect 21640 4088 21692 4140
rect 21824 4131 21876 4140
rect 21824 4097 21833 4131
rect 21833 4097 21867 4131
rect 21867 4097 21876 4131
rect 21824 4088 21876 4097
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 40592 4233 40601 4267
rect 40601 4233 40635 4267
rect 40635 4233 40644 4267
rect 40592 4224 40644 4233
rect 22192 3952 22244 4004
rect 22836 3952 22888 4004
rect 28448 4088 28500 4140
rect 24952 4020 25004 4072
rect 35900 4088 35952 4140
rect 38476 4088 38528 4140
rect 39856 4131 39908 4140
rect 39856 4097 39865 4131
rect 39865 4097 39899 4131
rect 39899 4097 39908 4131
rect 39856 4088 39908 4097
rect 40500 4131 40552 4140
rect 40500 4097 40509 4131
rect 40509 4097 40543 4131
rect 40543 4097 40552 4131
rect 40500 4088 40552 4097
rect 41052 4156 41104 4208
rect 45284 4224 45336 4276
rect 43720 4199 43772 4208
rect 43720 4165 43729 4199
rect 43729 4165 43763 4199
rect 43763 4165 43772 4199
rect 43720 4156 43772 4165
rect 46388 4156 46440 4208
rect 47768 4199 47820 4208
rect 47768 4165 47777 4199
rect 47777 4165 47811 4199
rect 47811 4165 47820 4199
rect 47768 4156 47820 4165
rect 33784 4020 33836 4072
rect 24860 3952 24912 4004
rect 41696 4020 41748 4072
rect 44916 4088 44968 4140
rect 45008 4020 45060 4072
rect 20168 3884 20220 3936
rect 21364 3884 21416 3936
rect 22744 3884 22796 3936
rect 23940 3927 23992 3936
rect 23940 3893 23949 3927
rect 23949 3893 23983 3927
rect 23983 3893 23992 3927
rect 23940 3884 23992 3893
rect 24768 3927 24820 3936
rect 24768 3893 24777 3927
rect 24777 3893 24811 3927
rect 24811 3893 24820 3927
rect 24768 3884 24820 3893
rect 25504 3927 25556 3936
rect 25504 3893 25513 3927
rect 25513 3893 25547 3927
rect 25547 3893 25556 3927
rect 25504 3884 25556 3893
rect 39580 3884 39632 3936
rect 41052 3952 41104 4004
rect 41512 3927 41564 3936
rect 41512 3893 41521 3927
rect 41521 3893 41555 3927
rect 41555 3893 41564 3927
rect 41512 3884 41564 3893
rect 42892 3884 42944 3936
rect 46296 3884 46348 3936
rect 46664 3927 46716 3936
rect 46664 3893 46673 3927
rect 46673 3893 46707 3927
rect 46707 3893 46716 3927
rect 46664 3884 46716 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 17684 3723 17736 3732
rect 6644 3612 6696 3664
rect 17684 3689 17693 3723
rect 17693 3689 17727 3723
rect 17727 3689 17736 3723
rect 17684 3680 17736 3689
rect 20720 3680 20772 3732
rect 1308 3476 1360 3528
rect 2136 3519 2188 3528
rect 2136 3485 2145 3519
rect 2145 3485 2179 3519
rect 2179 3485 2188 3519
rect 2136 3476 2188 3485
rect 7012 3544 7064 3596
rect 10324 3587 10376 3596
rect 7472 3519 7524 3528
rect 1768 3408 1820 3460
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 7932 3476 7984 3528
rect 8392 3408 8444 3460
rect 10324 3553 10333 3587
rect 10333 3553 10367 3587
rect 10367 3553 10376 3587
rect 10324 3544 10376 3553
rect 10508 3587 10560 3596
rect 10508 3553 10517 3587
rect 10517 3553 10551 3587
rect 10551 3553 10560 3587
rect 10508 3544 10560 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 17500 3544 17552 3596
rect 17960 3476 18012 3528
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 15476 3451 15528 3460
rect 15476 3417 15485 3451
rect 15485 3417 15519 3451
rect 15519 3417 15528 3451
rect 15476 3408 15528 3417
rect 17132 3451 17184 3460
rect 17132 3417 17141 3451
rect 17141 3417 17175 3451
rect 17175 3417 17184 3451
rect 17132 3408 17184 3417
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 1952 3340 2004 3392
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 13728 3340 13780 3392
rect 18328 3383 18380 3392
rect 18328 3349 18337 3383
rect 18337 3349 18371 3383
rect 18371 3349 18380 3383
rect 18328 3340 18380 3349
rect 20076 3612 20128 3664
rect 20168 3587 20220 3596
rect 20168 3553 20177 3587
rect 20177 3553 20211 3587
rect 20211 3553 20220 3587
rect 20168 3544 20220 3553
rect 20536 3612 20588 3664
rect 23020 3680 23072 3732
rect 23112 3680 23164 3732
rect 25872 3680 25924 3732
rect 39120 3680 39172 3732
rect 40500 3680 40552 3732
rect 22376 3612 22428 3664
rect 23388 3612 23440 3664
rect 20996 3544 21048 3596
rect 23940 3544 23992 3596
rect 25412 3587 25464 3596
rect 25412 3553 25421 3587
rect 25421 3553 25455 3587
rect 25455 3553 25464 3587
rect 25412 3544 25464 3553
rect 28908 3612 28960 3664
rect 45836 3680 45888 3732
rect 29552 3587 29604 3596
rect 19340 3519 19392 3528
rect 19340 3485 19349 3519
rect 19349 3485 19383 3519
rect 19383 3485 19392 3519
rect 19340 3476 19392 3485
rect 19984 3519 20036 3528
rect 19984 3485 19993 3519
rect 19993 3485 20027 3519
rect 20027 3485 20036 3519
rect 19984 3476 20036 3485
rect 22560 3476 22612 3528
rect 23204 3519 23256 3528
rect 23204 3485 23213 3519
rect 23213 3485 23247 3519
rect 23247 3485 23256 3519
rect 23204 3476 23256 3485
rect 20812 3340 20864 3392
rect 22652 3408 22704 3460
rect 24860 3476 24912 3528
rect 24492 3408 24544 3460
rect 25596 3451 25648 3460
rect 25596 3417 25605 3451
rect 25605 3417 25639 3451
rect 25639 3417 25648 3451
rect 25596 3408 25648 3417
rect 27252 3451 27304 3460
rect 27252 3417 27261 3451
rect 27261 3417 27295 3451
rect 27295 3417 27304 3451
rect 27252 3408 27304 3417
rect 24584 3340 24636 3392
rect 29552 3553 29561 3587
rect 29561 3553 29595 3587
rect 29595 3553 29604 3587
rect 29552 3544 29604 3553
rect 39948 3544 40000 3596
rect 40040 3587 40092 3596
rect 40040 3553 40049 3587
rect 40049 3553 40083 3587
rect 40083 3553 40092 3587
rect 40040 3544 40092 3553
rect 40684 3544 40736 3596
rect 41512 3587 41564 3596
rect 41512 3553 41521 3587
rect 41521 3553 41555 3587
rect 41555 3553 41564 3587
rect 41512 3544 41564 3553
rect 33784 3476 33836 3528
rect 35900 3519 35952 3528
rect 29736 3451 29788 3460
rect 29736 3417 29745 3451
rect 29745 3417 29779 3451
rect 29779 3417 29788 3451
rect 29736 3408 29788 3417
rect 32956 3408 33008 3460
rect 35900 3485 35909 3519
rect 35909 3485 35943 3519
rect 35943 3485 35952 3519
rect 35900 3476 35952 3485
rect 37740 3519 37792 3528
rect 37740 3485 37749 3519
rect 37749 3485 37783 3519
rect 37783 3485 37792 3519
rect 37740 3476 37792 3485
rect 39212 3476 39264 3528
rect 36176 3408 36228 3460
rect 39672 3408 39724 3460
rect 39764 3408 39816 3460
rect 41696 3451 41748 3460
rect 41696 3417 41705 3451
rect 41705 3417 41739 3451
rect 41739 3417 41748 3451
rect 41696 3408 41748 3417
rect 42708 3408 42760 3460
rect 45192 3519 45244 3528
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 47492 3612 47544 3664
rect 46296 3587 46348 3596
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 47676 3408 47728 3460
rect 48964 3408 49016 3460
rect 32220 3340 32272 3392
rect 33140 3383 33192 3392
rect 33140 3349 33149 3383
rect 33149 3349 33183 3383
rect 33183 3349 33192 3383
rect 33140 3340 33192 3349
rect 33876 3340 33928 3392
rect 42524 3340 42576 3392
rect 45376 3340 45428 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 1584 3136 1636 3188
rect 18236 3179 18288 3188
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 8116 3111 8168 3120
rect 8116 3077 8125 3111
rect 8125 3077 8159 3111
rect 8159 3077 8168 3111
rect 8116 3068 8168 3077
rect 13728 3111 13780 3120
rect 13728 3077 13737 3111
rect 13737 3077 13771 3111
rect 13771 3077 13780 3111
rect 13728 3068 13780 3077
rect 18236 3145 18245 3179
rect 18245 3145 18279 3179
rect 18279 3145 18288 3179
rect 18236 3136 18288 3145
rect 18880 3179 18932 3188
rect 18880 3145 18889 3179
rect 18889 3145 18923 3179
rect 18923 3145 18932 3179
rect 18880 3136 18932 3145
rect 19340 3136 19392 3188
rect 20536 3136 20588 3188
rect 22008 3136 22060 3188
rect 22192 3136 22244 3188
rect 22100 3068 22152 3120
rect 22744 3111 22796 3120
rect 22744 3077 22753 3111
rect 22753 3077 22787 3111
rect 22787 3077 22796 3111
rect 22744 3068 22796 3077
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 7932 3043 7984 3052
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 13544 3043 13596 3052
rect 664 2932 716 2984
rect 7748 2932 7800 2984
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 15200 2932 15252 2984
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 19984 3000 20036 3052
rect 21364 3000 21416 3052
rect 21916 3043 21968 3052
rect 21916 3009 21925 3043
rect 21925 3009 21959 3043
rect 21959 3009 21968 3043
rect 21916 3000 21968 3009
rect 22560 3043 22612 3052
rect 22560 3009 22569 3043
rect 22569 3009 22603 3043
rect 22603 3009 22612 3043
rect 22560 3000 22612 3009
rect 20628 2932 20680 2984
rect 20812 2932 20864 2984
rect 22100 2907 22152 2916
rect 10324 2839 10376 2848
rect 10324 2805 10333 2839
rect 10333 2805 10367 2839
rect 10367 2805 10376 2839
rect 10324 2796 10376 2805
rect 18696 2796 18748 2848
rect 20720 2796 20772 2848
rect 22100 2873 22109 2907
rect 22109 2873 22143 2907
rect 22143 2873 22152 2907
rect 22100 2864 22152 2873
rect 22468 2932 22520 2984
rect 23112 2932 23164 2984
rect 24676 3068 24728 3120
rect 35808 3136 35860 3188
rect 36176 3179 36228 3188
rect 36176 3145 36185 3179
rect 36185 3145 36219 3179
rect 36219 3145 36228 3179
rect 36176 3136 36228 3145
rect 39856 3136 39908 3188
rect 40132 3136 40184 3188
rect 25964 3111 26016 3120
rect 25964 3077 25973 3111
rect 25973 3077 26007 3111
rect 26007 3077 26016 3111
rect 25964 3068 26016 3077
rect 27620 3111 27672 3120
rect 27620 3077 27629 3111
rect 27629 3077 27663 3111
rect 27663 3077 27672 3111
rect 27620 3068 27672 3077
rect 33140 3111 33192 3120
rect 33140 3077 33149 3111
rect 33149 3077 33183 3111
rect 33183 3077 33192 3111
rect 33140 3068 33192 3077
rect 27068 3000 27120 3052
rect 32956 3043 33008 3052
rect 32956 3009 32965 3043
rect 32965 3009 32999 3043
rect 32999 3009 33008 3043
rect 32956 3000 33008 3009
rect 36084 3000 36136 3052
rect 38476 3043 38528 3052
rect 38476 3009 38485 3043
rect 38485 3009 38519 3043
rect 38519 3009 38528 3043
rect 38476 3000 38528 3009
rect 40592 3068 40644 3120
rect 42892 3111 42944 3120
rect 42892 3077 42901 3111
rect 42901 3077 42935 3111
rect 42935 3077 42944 3111
rect 42892 3068 42944 3077
rect 43168 3068 43220 3120
rect 45376 3111 45428 3120
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 42708 3043 42760 3052
rect 33508 2975 33560 2984
rect 23388 2864 23440 2916
rect 26056 2864 26108 2916
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 39764 2975 39816 2984
rect 39764 2941 39773 2975
rect 39773 2941 39807 2975
rect 39807 2941 39816 2975
rect 39764 2932 39816 2941
rect 39856 2932 39908 2984
rect 40684 2932 40736 2984
rect 42708 3009 42717 3043
rect 42717 3009 42751 3043
rect 42751 3009 42760 3043
rect 42708 3000 42760 3009
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 47768 3043 47820 3052
rect 47768 3009 47777 3043
rect 47777 3009 47811 3043
rect 47811 3009 47820 3043
rect 47768 3000 47820 3009
rect 46940 2932 46992 2984
rect 47676 2932 47728 2984
rect 27252 2796 27304 2848
rect 39672 2796 39724 2848
rect 40132 2796 40184 2848
rect 45008 2796 45060 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 15476 2592 15528 2644
rect 17960 2635 18012 2644
rect 17960 2601 17969 2635
rect 17969 2601 18003 2635
rect 18003 2601 18012 2635
rect 17960 2592 18012 2601
rect 18512 2592 18564 2644
rect 20904 2635 20956 2644
rect 20904 2601 20913 2635
rect 20913 2601 20947 2635
rect 20947 2601 20956 2635
rect 20904 2592 20956 2601
rect 21180 2592 21232 2644
rect 24952 2592 25004 2644
rect 26792 2592 26844 2644
rect 29736 2635 29788 2644
rect 29736 2601 29745 2635
rect 29745 2601 29779 2635
rect 29779 2601 29788 2635
rect 29736 2592 29788 2601
rect 39212 2635 39264 2644
rect 39212 2601 39221 2635
rect 39221 2601 39255 2635
rect 39255 2601 39264 2635
rect 39212 2592 39264 2601
rect 40408 2635 40460 2644
rect 40408 2601 40417 2635
rect 40417 2601 40451 2635
rect 40451 2601 40460 2635
rect 40408 2592 40460 2601
rect 2780 2524 2832 2576
rect 1676 2456 1728 2508
rect 2872 2499 2924 2508
rect 2872 2465 2881 2499
rect 2881 2465 2915 2499
rect 2915 2465 2924 2499
rect 2872 2456 2924 2465
rect 15200 2524 15252 2576
rect 17592 2524 17644 2576
rect 21088 2524 21140 2576
rect 6736 2499 6788 2508
rect 6736 2465 6745 2499
rect 6745 2465 6779 2499
rect 6779 2465 6788 2499
rect 6736 2456 6788 2465
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 9128 2499 9180 2508
rect 9128 2465 9137 2499
rect 9137 2465 9171 2499
rect 9171 2465 9180 2499
rect 9128 2456 9180 2465
rect 10324 2456 10376 2508
rect 2596 2320 2648 2372
rect 5172 2388 5224 2440
rect 7472 2320 7524 2372
rect 9036 2320 9088 2372
rect 20720 2456 20772 2508
rect 25504 2524 25556 2576
rect 25596 2524 25648 2576
rect 45284 2524 45336 2576
rect 15476 2388 15528 2440
rect 18328 2388 18380 2440
rect 18604 2388 18656 2440
rect 20996 2388 21048 2440
rect 22100 2431 22152 2440
rect 22100 2397 22109 2431
rect 22109 2397 22143 2431
rect 22143 2397 22152 2431
rect 22100 2388 22152 2397
rect 24768 2499 24820 2508
rect 24768 2465 24777 2499
rect 24777 2465 24811 2499
rect 24811 2465 24820 2499
rect 24768 2456 24820 2465
rect 25136 2499 25188 2508
rect 25136 2465 25145 2499
rect 25145 2465 25179 2499
rect 25179 2465 25188 2499
rect 25136 2456 25188 2465
rect 35808 2499 35860 2508
rect 35808 2465 35817 2499
rect 35817 2465 35851 2499
rect 35851 2465 35860 2499
rect 35808 2456 35860 2465
rect 41696 2456 41748 2508
rect 45100 2456 45152 2508
rect 45744 2456 45796 2508
rect 45836 2499 45888 2508
rect 45836 2465 45845 2499
rect 45845 2465 45879 2499
rect 45879 2465 45888 2499
rect 45836 2456 45888 2465
rect 26424 2388 26476 2440
rect 16120 2320 16172 2372
rect 20628 2320 20680 2372
rect 24032 2320 24084 2372
rect 29644 2388 29696 2440
rect 35440 2388 35492 2440
rect 38016 2388 38068 2440
rect 39580 2388 39632 2440
rect 41236 2388 41288 2440
rect 28356 2320 28408 2372
rect 29828 2320 29880 2372
rect 16856 2252 16908 2304
rect 29460 2252 29512 2304
rect 39304 2320 39356 2372
rect 40592 2320 40644 2372
rect 45468 2320 45520 2372
rect 47952 2320 48004 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4844 49314
rect 4498 49200 4610 49286
rect 32 21418 60 49200
rect 1398 47696 1454 47705
rect 1398 47631 1454 47640
rect 1412 46578 1440 47631
rect 1964 47054 1992 49200
rect 2608 47054 2636 49200
rect 3252 47054 3280 49200
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2596 47048 2648 47054
rect 2596 46990 2648 46996
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3422 47016 3478 47025
rect 3422 46951 3478 46960
rect 2136 46912 2188 46918
rect 2136 46854 2188 46860
rect 2872 46912 2924 46918
rect 2872 46854 2924 46860
rect 1400 46572 1452 46578
rect 1400 46514 1452 46520
rect 1676 46368 1728 46374
rect 1676 46310 1728 46316
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1584 41540 1636 41546
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1400 40520 1452 40526
rect 1400 40462 1452 40468
rect 1412 40225 1440 40462
rect 1398 40216 1454 40225
rect 1398 40151 1454 40160
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1492 35488 1544 35494
rect 1596 35465 1624 35634
rect 1492 35430 1544 35436
rect 1582 35456 1638 35465
rect 1308 33992 1360 33998
rect 1308 33934 1360 33940
rect 1320 32745 1348 33934
rect 1400 33448 1452 33454
rect 1398 33416 1400 33425
rect 1452 33416 1454 33425
rect 1398 33351 1454 33360
rect 1504 33046 1532 35430
rect 1582 35391 1638 35400
rect 1584 33856 1636 33862
rect 1584 33798 1636 33804
rect 1492 33040 1544 33046
rect 1492 32982 1544 32988
rect 1596 32978 1624 33798
rect 1584 32972 1636 32978
rect 1584 32914 1636 32920
rect 1306 32736 1362 32745
rect 1306 32671 1362 32680
rect 1400 32224 1452 32230
rect 1400 32166 1452 32172
rect 1412 31890 1440 32166
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1596 31482 1624 31690
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 1688 28218 1716 46310
rect 1860 43308 1912 43314
rect 1860 43250 1912 43256
rect 1872 42945 1900 43250
rect 1952 43104 2004 43110
rect 1952 43046 2004 43052
rect 1858 42936 1914 42945
rect 1858 42871 1914 42880
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1780 36786 1808 37198
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1964 35894 1992 43046
rect 2148 40458 2176 46854
rect 2884 46646 2912 46854
rect 2872 46640 2924 46646
rect 2872 46582 2924 46588
rect 2320 46368 2372 46374
rect 2320 46310 2372 46316
rect 2778 46336 2834 46345
rect 2332 46034 2360 46310
rect 2778 46271 2834 46280
rect 2792 46034 2820 46271
rect 2320 46028 2372 46034
rect 2320 45970 2372 45976
rect 2780 46028 2832 46034
rect 2780 45970 2832 45976
rect 2228 45892 2280 45898
rect 2228 45834 2280 45840
rect 2240 45626 2268 45834
rect 2228 45620 2280 45626
rect 2228 45562 2280 45568
rect 2412 45484 2464 45490
rect 2412 45426 2464 45432
rect 2136 40452 2188 40458
rect 2136 40394 2188 40400
rect 2228 36712 2280 36718
rect 2228 36654 2280 36660
rect 2240 36378 2268 36654
rect 2228 36372 2280 36378
rect 2228 36314 2280 36320
rect 2228 36168 2280 36174
rect 2228 36110 2280 36116
rect 1964 35866 2084 35894
rect 1858 32056 1914 32065
rect 1858 31991 1914 32000
rect 1872 31890 1900 31991
rect 1860 31884 1912 31890
rect 1860 31826 1912 31832
rect 1676 28212 1728 28218
rect 1676 28154 1728 28160
rect 1400 25288 1452 25294
rect 1398 25256 1400 25265
rect 1452 25256 1454 25265
rect 1398 25191 1454 25200
rect 1676 25220 1728 25226
rect 1676 25162 1728 25168
rect 20 21412 72 21418
rect 20 21354 72 21360
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1688 6730 1716 25162
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 23225 1900 23666
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1872 17785 1900 18226
rect 1858 17776 1914 17785
rect 1858 17711 1914 17720
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1872 16425 1900 16594
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1964 6914 1992 16050
rect 2056 15638 2084 35866
rect 2136 31340 2188 31346
rect 2136 31282 2188 31288
rect 2148 23186 2176 31282
rect 2136 23180 2188 23186
rect 2136 23122 2188 23128
rect 2240 20074 2268 36110
rect 2320 32360 2372 32366
rect 2320 32302 2372 32308
rect 2148 20046 2268 20074
rect 2148 18766 2176 20046
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2332 16658 2360 32302
rect 2424 31346 2452 45426
rect 2962 44976 3018 44985
rect 2962 44911 3018 44920
rect 2976 44266 3004 44911
rect 2964 44260 3016 44266
rect 2964 44202 3016 44208
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36718 2820 36751
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 2504 33448 2556 33454
rect 2504 33390 2556 33396
rect 2516 32502 2544 33390
rect 2504 32496 2556 32502
rect 2504 32438 2556 32444
rect 2412 31340 2464 31346
rect 2412 31282 2464 31288
rect 3330 28656 3386 28665
rect 3330 28591 3386 28600
rect 3344 27946 3372 28591
rect 3332 27940 3384 27946
rect 3332 27882 3384 27888
rect 3436 22386 3464 46951
rect 3896 46442 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4816 47054 4844 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49200 7186 50000
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49314 13626 50000
rect 13514 49286 13768 49314
rect 13514 49200 13626 49286
rect 5828 47054 5856 49200
rect 7116 47054 7144 49200
rect 4804 47048 4856 47054
rect 4804 46990 4856 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7104 47048 7156 47054
rect 7104 46990 7156 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 5080 46980 5132 46986
rect 5080 46922 5132 46928
rect 7840 46980 7892 46986
rect 7840 46922 7892 46928
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 3884 46436 3936 46442
rect 3884 46378 3936 46384
rect 3988 46170 4016 46446
rect 3976 46164 4028 46170
rect 3976 46106 4028 46112
rect 3514 43616 3570 43625
rect 3514 43551 3570 43560
rect 3528 22506 3556 43551
rect 3698 39536 3754 39545
rect 3698 39471 3754 39480
rect 3606 31376 3662 31385
rect 3606 31311 3662 31320
rect 3516 22500 3568 22506
rect 3516 22442 3568 22448
rect 3436 22358 3556 22386
rect 3528 19446 3556 22358
rect 3620 21010 3648 31311
rect 3712 22778 3740 39471
rect 3976 32836 4028 32842
rect 3976 32778 4028 32784
rect 3988 32366 4016 32778
rect 3976 32360 4028 32366
rect 3976 32302 4028 32308
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 3988 22094 4016 32302
rect 3896 22066 4016 22094
rect 3608 21004 3660 21010
rect 3608 20946 3660 20952
rect 3516 19440 3568 19446
rect 3516 19382 3568 19388
rect 3332 17128 3384 17134
rect 3330 17096 3332 17105
rect 3384 17096 3386 17105
rect 3330 17031 3386 17040
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 2148 16250 2176 16458
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2044 15632 2096 15638
rect 2044 15574 2096 15580
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2148 14074 2176 14350
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 1964 6886 2084 6914
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 2056 4146 2084 6886
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1320 800 1348 3470
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1596 3194 1624 3334
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1688 2514 1716 3878
rect 2148 3534 2176 14010
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7585 3004 8230
rect 2962 7576 3018 7585
rect 2962 7511 3018 7520
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 1768 3460 1820 3466
rect 1768 3402 1820 3408
rect 1780 3058 1808 3402
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1964 3126 1992 3334
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2792 2582 2820 3878
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2608 800 2636 2314
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 2884 785 2912 2450
rect 3344 898 3372 11290
rect 3436 4162 3464 16594
rect 3896 14482 3924 22066
rect 3976 19916 4028 19922
rect 3976 19858 4028 19864
rect 3988 19825 4016 19858
rect 3974 19816 4030 19825
rect 3974 19751 4030 19760
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3988 18465 4016 18906
rect 3974 18456 4030 18465
rect 3974 18391 4030 18400
rect 3884 14476 3936 14482
rect 3884 14418 3936 14424
rect 3976 13728 4028 13734
rect 3974 13696 3976 13705
rect 4028 13696 4030 13705
rect 3974 13631 4030 13640
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 10305 3556 10406
rect 3514 10296 3570 10305
rect 3514 10231 3570 10240
rect 4080 6914 4108 46922
rect 4988 46504 5040 46510
rect 4988 46446 5040 46452
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 5000 46170 5028 46446
rect 4988 46164 5040 46170
rect 4988 46106 5040 46112
rect 4896 45960 4948 45966
rect 4896 45902 4948 45908
rect 4908 45354 4936 45902
rect 4896 45348 4948 45354
rect 4896 45290 4948 45296
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 5092 26234 5120 46922
rect 6920 46912 6972 46918
rect 6920 46854 6972 46860
rect 5000 26206 5120 26234
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 5000 17338 5028 26206
rect 6932 22094 6960 46854
rect 7852 29034 7880 46922
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9496 46980 9548 46986
rect 9496 46922 9548 46928
rect 8312 45526 8432 45554
rect 8312 30122 8340 45526
rect 9508 36922 9536 46922
rect 10600 46368 10652 46374
rect 10600 46310 10652 46316
rect 10612 46034 10640 46310
rect 10980 46034 11008 49200
rect 11624 46578 11652 49200
rect 12268 47122 12296 49200
rect 12256 47116 12308 47122
rect 12256 47058 12308 47064
rect 12624 47048 12676 47054
rect 12624 46990 12676 46996
rect 11612 46572 11664 46578
rect 11612 46514 11664 46520
rect 10600 46028 10652 46034
rect 10600 45970 10652 45976
rect 10968 46028 11020 46034
rect 10968 45970 11020 45976
rect 10784 45892 10836 45898
rect 10784 45834 10836 45840
rect 10796 45626 10824 45834
rect 10784 45620 10836 45626
rect 10784 45562 10836 45568
rect 10968 40384 11020 40390
rect 10968 40326 11020 40332
rect 9496 36916 9548 36922
rect 9496 36858 9548 36864
rect 10980 36310 11008 40326
rect 12636 37126 12664 46990
rect 12912 45966 12940 49200
rect 13740 47138 13768 49286
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49314 16202 50000
rect 16090 49286 16528 49314
rect 16090 49200 16202 49286
rect 14200 47274 14228 49200
rect 14200 47246 14320 47274
rect 13740 47122 13860 47138
rect 13740 47116 13872 47122
rect 13740 47110 13820 47116
rect 13820 47058 13872 47064
rect 14292 46510 14320 47246
rect 14464 47048 14516 47054
rect 14464 46990 14516 46996
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 14200 46170 14228 46446
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 12900 45960 12952 45966
rect 12900 45902 12952 45908
rect 14096 45960 14148 45966
rect 14096 45902 14148 45908
rect 14108 41138 14136 45902
rect 14476 41414 14504 46990
rect 15488 45554 15516 49200
rect 16500 47054 16528 49286
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49314 25218 50000
rect 25106 49286 25452 49314
rect 25106 49200 25218 49286
rect 17420 47410 17448 49200
rect 16776 47382 17448 47410
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 15488 45526 15976 45554
rect 14476 41386 14596 41414
rect 14096 41132 14148 41138
rect 14096 41074 14148 41080
rect 14188 37256 14240 37262
rect 14188 37198 14240 37204
rect 12624 37120 12676 37126
rect 12624 37062 12676 37068
rect 14200 36718 14228 37198
rect 14188 36712 14240 36718
rect 14188 36654 14240 36660
rect 10968 36304 11020 36310
rect 10968 36246 11020 36252
rect 14200 35630 14228 36654
rect 14188 35624 14240 35630
rect 14188 35566 14240 35572
rect 14200 35086 14228 35566
rect 14188 35080 14240 35086
rect 14188 35022 14240 35028
rect 14200 33998 14228 35022
rect 14464 35012 14516 35018
rect 14464 34954 14516 34960
rect 14476 34746 14504 34954
rect 14464 34740 14516 34746
rect 14464 34682 14516 34688
rect 14188 33992 14240 33998
rect 14188 33934 14240 33940
rect 14200 31890 14228 33934
rect 14464 33924 14516 33930
rect 14464 33866 14516 33872
rect 14476 33658 14504 33866
rect 14464 33652 14516 33658
rect 14464 33594 14516 33600
rect 14188 31884 14240 31890
rect 14188 31826 14240 31832
rect 14568 30802 14596 41386
rect 15292 37868 15344 37874
rect 15292 37810 15344 37816
rect 15200 36848 15252 36854
rect 15200 36790 15252 36796
rect 15212 36378 15240 36790
rect 15200 36372 15252 36378
rect 15200 36314 15252 36320
rect 15304 36174 15332 37810
rect 15844 37732 15896 37738
rect 15844 37674 15896 37680
rect 15856 37330 15884 37674
rect 15844 37324 15896 37330
rect 15844 37266 15896 37272
rect 15568 36372 15620 36378
rect 15568 36314 15620 36320
rect 15580 36242 15608 36314
rect 15568 36236 15620 36242
rect 15568 36178 15620 36184
rect 15292 36168 15344 36174
rect 15292 36110 15344 36116
rect 15304 36038 15332 36110
rect 15292 36032 15344 36038
rect 15292 35974 15344 35980
rect 15304 32434 15332 35974
rect 15476 35488 15528 35494
rect 15476 35430 15528 35436
rect 15488 35018 15516 35430
rect 15476 35012 15528 35018
rect 15476 34954 15528 34960
rect 15476 34604 15528 34610
rect 15580 34592 15608 36178
rect 15844 34944 15896 34950
rect 15844 34886 15896 34892
rect 15856 34610 15884 34886
rect 15528 34564 15608 34592
rect 15844 34604 15896 34610
rect 15476 34546 15528 34552
rect 15844 34546 15896 34552
rect 15752 34536 15804 34542
rect 15580 34496 15752 34524
rect 15292 32428 15344 32434
rect 15292 32370 15344 32376
rect 15304 31754 15332 32370
rect 15304 31726 15516 31754
rect 15488 31482 15516 31726
rect 15476 31476 15528 31482
rect 15476 31418 15528 31424
rect 14556 30796 14608 30802
rect 14556 30738 14608 30744
rect 15488 30734 15516 31418
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 12992 30184 13044 30190
rect 12992 30126 13044 30132
rect 13452 30184 13504 30190
rect 13452 30126 13504 30132
rect 8300 30116 8352 30122
rect 8300 30058 8352 30064
rect 11704 29096 11756 29102
rect 11704 29038 11756 29044
rect 7840 29028 7892 29034
rect 7840 28970 7892 28976
rect 11612 28620 11664 28626
rect 11612 28562 11664 28568
rect 10876 28552 10928 28558
rect 10876 28494 10928 28500
rect 10888 28218 10916 28494
rect 11624 28218 11652 28562
rect 10876 28212 10928 28218
rect 10876 28154 10928 28160
rect 11612 28212 11664 28218
rect 11612 28154 11664 28160
rect 11716 28082 11744 29038
rect 11980 28756 12032 28762
rect 11980 28698 12032 28704
rect 10508 28076 10560 28082
rect 10508 28018 10560 28024
rect 11520 28076 11572 28082
rect 11520 28018 11572 28024
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 10520 26994 10548 28018
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 10784 27328 10836 27334
rect 10784 27270 10836 27276
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 10520 26874 10548 26930
rect 10428 26846 10548 26874
rect 10428 25906 10456 26846
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10520 26450 10548 26726
rect 10796 26450 10824 27270
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10784 26444 10836 26450
rect 10784 26386 10836 26392
rect 11164 26042 11192 27406
rect 11532 27130 11560 28018
rect 11520 27124 11572 27130
rect 11520 27066 11572 27072
rect 11716 27062 11744 28018
rect 11428 27056 11480 27062
rect 11428 26998 11480 27004
rect 11704 27056 11756 27062
rect 11704 26998 11756 27004
rect 11440 26246 11468 26998
rect 11992 26994 12020 28698
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 12544 28218 12572 28426
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12360 27470 12388 28018
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 12440 27396 12492 27402
rect 12440 27338 12492 27344
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 11980 26988 12032 26994
rect 11980 26930 12032 26936
rect 11888 26852 11940 26858
rect 11888 26794 11940 26800
rect 11428 26240 11480 26246
rect 11428 26182 11480 26188
rect 11152 26036 11204 26042
rect 11152 25978 11204 25984
rect 11440 25974 11468 26182
rect 11428 25968 11480 25974
rect 11428 25910 11480 25916
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 10968 25900 11020 25906
rect 10968 25842 11020 25848
rect 9404 25696 9456 25702
rect 9404 25638 9456 25644
rect 9416 25362 9444 25638
rect 10428 25378 10456 25842
rect 9404 25356 9456 25362
rect 9404 25298 9456 25304
rect 10336 25350 10456 25378
rect 9680 25220 9732 25226
rect 9680 25162 9732 25168
rect 9692 24682 9720 25162
rect 9956 24744 10008 24750
rect 9956 24686 10008 24692
rect 9680 24676 9732 24682
rect 9680 24618 9732 24624
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7932 23656 7984 23662
rect 7932 23598 7984 23604
rect 7668 23322 7696 23598
rect 7656 23316 7708 23322
rect 7656 23258 7708 23264
rect 7656 23112 7708 23118
rect 7656 23054 7708 23060
rect 7668 22658 7696 23054
rect 7484 22642 7696 22658
rect 7472 22636 7696 22642
rect 7524 22630 7696 22636
rect 7472 22578 7524 22584
rect 7668 22094 7696 22630
rect 6932 22066 7052 22094
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3514 6896 3570 6905
rect 3514 6831 3516 6840
rect 3568 6831 3570 6840
rect 3988 6886 4108 6914
rect 3516 6802 3568 6808
rect 3436 4134 3556 4162
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3436 3505 3464 4014
rect 3422 3496 3478 3505
rect 3422 3431 3478 3440
rect 3528 1465 3556 4134
rect 3988 3641 4016 6886
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3974 3632 4030 3641
rect 3974 3567 4030 3576
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 3514 1456 3570 1465
rect 3514 1391 3570 1400
rect 3344 870 3556 898
rect 2870 776 2926 785
rect 2870 711 2926 720
rect 3210 0 3322 800
rect 3528 762 3556 870
rect 3712 870 3924 898
rect 3712 762 3740 870
rect 3896 800 3924 870
rect 5184 800 5212 2382
rect 6472 800 6500 6122
rect 6656 3670 6684 18634
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6390 6960 6598
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5914 6960 6190
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 7024 3602 7052 22066
rect 7576 22066 7696 22094
rect 7576 22030 7604 22066
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7472 21888 7524 21894
rect 7472 21830 7524 21836
rect 7484 21622 7512 21830
rect 7576 21622 7604 21966
rect 7472 21616 7524 21622
rect 7472 21558 7524 21564
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7944 17134 7972 23598
rect 9968 23118 9996 24686
rect 10336 23730 10364 25350
rect 10416 25220 10468 25226
rect 10416 25162 10468 25168
rect 10428 24410 10456 25162
rect 10980 24750 11008 25842
rect 11440 25226 11468 25910
rect 11900 25906 11928 26794
rect 11888 25900 11940 25906
rect 11888 25842 11940 25848
rect 11428 25220 11480 25226
rect 11428 25162 11480 25168
rect 11440 24818 11468 25162
rect 11428 24812 11480 24818
rect 11428 24754 11480 24760
rect 10968 24744 11020 24750
rect 10968 24686 11020 24692
rect 10980 24614 11008 24686
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 10324 23724 10376 23730
rect 10244 23684 10324 23712
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8956 22098 8984 22918
rect 9312 22568 9364 22574
rect 9312 22510 9364 22516
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9232 21690 9260 21898
rect 9324 21894 9352 22510
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9128 21684 9180 21690
rect 9128 21626 9180 21632
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9140 19786 9168 21626
rect 9324 21486 9352 21830
rect 9312 21480 9364 21486
rect 9312 21422 9364 21428
rect 9324 20874 9352 21422
rect 9692 21418 9720 23054
rect 10244 22982 10272 23684
rect 10324 23666 10376 23672
rect 10324 23520 10376 23526
rect 10324 23462 10376 23468
rect 10336 23118 10364 23462
rect 10324 23112 10376 23118
rect 10324 23054 10376 23060
rect 10232 22976 10284 22982
rect 10232 22918 10284 22924
rect 10244 22778 10272 22918
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 10428 22438 10456 24142
rect 11900 23798 11928 25842
rect 11992 25838 12020 26930
rect 12084 26314 12112 27270
rect 12452 27130 12480 27338
rect 13004 27282 13032 30126
rect 13464 29306 13492 30126
rect 13820 29640 13872 29646
rect 13820 29582 13872 29588
rect 13452 29300 13504 29306
rect 13452 29242 13504 29248
rect 13832 29170 13860 29582
rect 14280 29504 14332 29510
rect 14280 29446 14332 29452
rect 14924 29504 14976 29510
rect 14924 29446 14976 29452
rect 14292 29238 14320 29446
rect 14280 29232 14332 29238
rect 14280 29174 14332 29180
rect 13820 29164 13872 29170
rect 13820 29106 13872 29112
rect 13268 28620 13320 28626
rect 13268 28562 13320 28568
rect 13004 27254 13216 27282
rect 12440 27124 12492 27130
rect 12440 27066 12492 27072
rect 12256 26852 12308 26858
rect 12256 26794 12308 26800
rect 12268 26586 12296 26794
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 12268 26314 12296 26522
rect 13004 26314 13032 27254
rect 13188 27130 13216 27254
rect 13084 27124 13136 27130
rect 13084 27066 13136 27072
rect 13176 27124 13228 27130
rect 13176 27066 13228 27072
rect 12072 26308 12124 26314
rect 12072 26250 12124 26256
rect 12256 26308 12308 26314
rect 12256 26250 12308 26256
rect 12992 26308 13044 26314
rect 12992 26250 13044 26256
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 11980 25832 12032 25838
rect 11980 25774 12032 25780
rect 12820 24274 12848 25842
rect 13004 25770 13032 26250
rect 13096 25906 13124 27066
rect 13176 26920 13228 26926
rect 13176 26862 13228 26868
rect 13188 26042 13216 26862
rect 13280 26382 13308 28562
rect 13832 27538 13860 29106
rect 14936 28626 14964 29446
rect 14924 28620 14976 28626
rect 14924 28562 14976 28568
rect 14096 28008 14148 28014
rect 14464 28008 14516 28014
rect 14096 27950 14148 27956
rect 13820 27532 13872 27538
rect 13820 27474 13872 27480
rect 13912 27464 13964 27470
rect 13912 27406 13964 27412
rect 13452 27056 13504 27062
rect 13452 26998 13504 27004
rect 13464 26450 13492 26998
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 13452 26444 13504 26450
rect 13452 26386 13504 26392
rect 13268 26376 13320 26382
rect 13268 26318 13320 26324
rect 13452 26308 13504 26314
rect 13452 26250 13504 26256
rect 13176 26036 13228 26042
rect 13176 25978 13228 25984
rect 13464 25974 13492 26250
rect 13832 26042 13860 26726
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13452 25968 13504 25974
rect 13452 25910 13504 25916
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 12992 25764 13044 25770
rect 12992 25706 13044 25712
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13096 24342 13124 24686
rect 13372 24410 13400 24686
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 12992 24336 13044 24342
rect 12992 24278 13044 24284
rect 13084 24336 13136 24342
rect 13084 24278 13136 24284
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 13004 24206 13032 24278
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 11888 23792 11940 23798
rect 11888 23734 11940 23740
rect 12820 23730 12848 24074
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 13004 23798 13032 24006
rect 12992 23792 13044 23798
rect 12992 23734 13044 23740
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 11888 23656 11940 23662
rect 11888 23598 11940 23604
rect 11520 22976 11572 22982
rect 11520 22918 11572 22924
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 10416 22432 10468 22438
rect 10416 22374 10468 22380
rect 9968 21962 9996 22374
rect 11440 22098 11468 22578
rect 11532 22574 11560 22918
rect 11520 22568 11572 22574
rect 11520 22510 11572 22516
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 11428 22092 11480 22098
rect 11428 22034 11480 22040
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9680 21412 9732 21418
rect 9680 21354 9732 21360
rect 9784 21350 9812 21626
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10232 21480 10284 21486
rect 10232 21422 10284 21428
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9312 20868 9364 20874
rect 9312 20810 9364 20816
rect 10244 20806 10272 21422
rect 10980 21350 11008 21490
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 9692 20398 9720 20742
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 9692 19378 9720 20334
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9968 19990 9996 20198
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 10244 19854 10272 20742
rect 10336 20466 10364 21286
rect 10980 21146 11008 21286
rect 10600 21140 10652 21146
rect 10600 21082 10652 21088
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10968 21140 11020 21146
rect 10968 21082 11020 21088
rect 10612 20874 10640 21082
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10612 20602 10640 20810
rect 10600 20596 10652 20602
rect 10600 20538 10652 20544
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10336 19922 10364 20402
rect 10796 20398 10824 21082
rect 11072 21078 11100 21422
rect 11164 21078 11192 21966
rect 11532 21962 11560 22510
rect 11716 22234 11744 22510
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 11796 22228 11848 22234
rect 11796 22170 11848 22176
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11532 21622 11560 21898
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11520 21616 11572 21622
rect 11520 21558 11572 21564
rect 11060 21072 11112 21078
rect 11060 21014 11112 21020
rect 11152 21072 11204 21078
rect 11152 21014 11204 21020
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9324 18834 9352 19110
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 9048 18426 9076 18702
rect 9416 18698 9444 18770
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9692 18630 9720 19314
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9232 10470 9260 15506
rect 9692 15502 9720 18566
rect 9876 18290 9904 19314
rect 10336 19310 10364 19858
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10612 19378 10640 19790
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10796 19378 10824 19654
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10336 18426 10364 18634
rect 11164 18578 11192 21014
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11624 20058 11652 20334
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11348 18834 11376 19110
rect 11624 18834 11652 19450
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11072 18550 11192 18578
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10704 16590 10732 16934
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10876 16516 10928 16522
rect 10876 16458 10928 16464
rect 10888 16250 10916 16458
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 11072 16114 11100 18550
rect 11716 18290 11744 21830
rect 11808 21486 11836 22170
rect 11900 22030 11928 23598
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 11992 22438 12020 23054
rect 12268 22982 12296 23462
rect 12256 22976 12308 22982
rect 12256 22918 12308 22924
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13464 22710 13492 22918
rect 13452 22704 13504 22710
rect 13452 22646 13504 22652
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11900 21554 11928 21966
rect 11992 21894 12020 22374
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 12268 21350 12296 22034
rect 13648 21894 13676 25298
rect 13924 25294 13952 27406
rect 14004 25900 14056 25906
rect 14004 25842 14056 25848
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13728 25220 13780 25226
rect 13728 25162 13780 25168
rect 13740 24138 13768 25162
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13740 23866 13768 24074
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 11992 19378 12020 21286
rect 12360 20482 12388 21490
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 12360 20454 12480 20482
rect 12452 20398 12480 20454
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12360 20058 12388 20334
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12072 19780 12124 19786
rect 12072 19722 12124 19728
rect 12084 19514 12112 19722
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12084 19378 12112 19450
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 12084 18426 12112 18634
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 12452 17678 12480 19314
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 12912 18834 12940 19110
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 13004 18630 13032 19110
rect 13096 18630 13124 20538
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13464 19242 13492 19654
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13464 18630 13492 19178
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12728 17202 12756 17478
rect 13004 17270 13032 17478
rect 12992 17264 13044 17270
rect 12992 17206 13044 17212
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 13096 16658 13124 18566
rect 13464 18290 13492 18566
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13648 18222 13676 18634
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13372 17678 13400 18158
rect 13832 17762 13860 23598
rect 13924 23118 13952 25230
rect 14016 25226 14044 25842
rect 14108 25770 14136 27950
rect 14200 27946 14412 27962
rect 15580 27962 15608 34496
rect 15752 34478 15804 34484
rect 15660 32224 15712 32230
rect 15660 32166 15712 32172
rect 15672 31822 15700 32166
rect 15660 31816 15712 31822
rect 15660 31758 15712 31764
rect 15660 31408 15712 31414
rect 15660 31350 15712 31356
rect 15672 30938 15700 31350
rect 15660 30932 15712 30938
rect 15660 30874 15712 30880
rect 15948 29238 15976 45526
rect 16776 41414 16804 47382
rect 18708 47054 18736 49200
rect 19996 48226 20024 49200
rect 19996 48198 20116 48226
rect 19984 47184 20036 47190
rect 19984 47126 20036 47132
rect 18696 47048 18748 47054
rect 18696 46990 18748 46996
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19616 46504 19668 46510
rect 19616 46446 19668 46452
rect 17224 46368 17276 46374
rect 17224 46310 17276 46316
rect 16684 41386 16804 41414
rect 16580 37664 16632 37670
rect 16580 37606 16632 37612
rect 16592 37194 16620 37606
rect 16580 37188 16632 37194
rect 16580 37130 16632 37136
rect 16488 36712 16540 36718
rect 16488 36654 16540 36660
rect 16028 36644 16080 36650
rect 16028 36586 16080 36592
rect 16040 36242 16068 36586
rect 16500 36378 16528 36654
rect 16684 36530 16712 41386
rect 16856 38208 16908 38214
rect 16856 38150 16908 38156
rect 16868 37874 16896 38150
rect 17236 37942 17264 46310
rect 19628 46170 19656 46446
rect 19616 46164 19668 46170
rect 19616 46106 19668 46112
rect 18972 45960 19024 45966
rect 18972 45902 19024 45908
rect 18984 41414 19012 45902
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19996 45554 20024 47126
rect 20088 47122 20116 48198
rect 20076 47116 20128 47122
rect 20076 47058 20128 47064
rect 20536 47116 20588 47122
rect 20536 47058 20588 47064
rect 20352 47048 20404 47054
rect 20352 46990 20404 46996
rect 20168 46980 20220 46986
rect 20168 46922 20220 46928
rect 20076 46436 20128 46442
rect 20076 46378 20128 46384
rect 20088 46170 20116 46378
rect 20076 46164 20128 46170
rect 20076 46106 20128 46112
rect 19996 45526 20116 45554
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 18984 41386 19196 41414
rect 18328 38412 18380 38418
rect 18328 38354 18380 38360
rect 17500 38208 17552 38214
rect 17500 38150 17552 38156
rect 17592 38208 17644 38214
rect 17592 38150 17644 38156
rect 17224 37936 17276 37942
rect 17224 37878 17276 37884
rect 16856 37868 16908 37874
rect 16856 37810 16908 37816
rect 17512 37466 17540 38150
rect 17604 38010 17632 38150
rect 17592 38004 17644 38010
rect 17592 37946 17644 37952
rect 18052 37800 18104 37806
rect 18052 37742 18104 37748
rect 18064 37466 18092 37742
rect 17500 37460 17552 37466
rect 17500 37402 17552 37408
rect 18052 37460 18104 37466
rect 18052 37402 18104 37408
rect 17512 37262 17540 37402
rect 18052 37324 18104 37330
rect 18052 37266 18104 37272
rect 17500 37256 17552 37262
rect 17500 37198 17552 37204
rect 17512 36786 17540 37198
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 18064 36718 18092 37266
rect 18052 36712 18104 36718
rect 18052 36654 18104 36660
rect 16592 36502 16712 36530
rect 17408 36576 17460 36582
rect 17408 36518 17460 36524
rect 16488 36372 16540 36378
rect 16488 36314 16540 36320
rect 16028 36236 16080 36242
rect 16028 36178 16080 36184
rect 16488 36236 16540 36242
rect 16488 36178 16540 36184
rect 16212 36168 16264 36174
rect 16212 36110 16264 36116
rect 16224 34626 16252 36110
rect 16500 36038 16528 36178
rect 16488 36032 16540 36038
rect 16488 35974 16540 35980
rect 16396 35692 16448 35698
rect 16396 35634 16448 35640
rect 16132 34610 16252 34626
rect 16120 34604 16252 34610
rect 16172 34598 16252 34604
rect 16120 34546 16172 34552
rect 16224 34066 16252 34598
rect 16212 34060 16264 34066
rect 16212 34002 16264 34008
rect 16408 33998 16436 35634
rect 16396 33992 16448 33998
rect 16396 33934 16448 33940
rect 16396 33856 16448 33862
rect 16396 33798 16448 33804
rect 16408 33658 16436 33798
rect 16396 33652 16448 33658
rect 16396 33594 16448 33600
rect 16408 32910 16436 33594
rect 16396 32904 16448 32910
rect 16396 32846 16448 32852
rect 16028 31136 16080 31142
rect 16028 31078 16080 31084
rect 15936 29232 15988 29238
rect 15936 29174 15988 29180
rect 16040 28626 16068 31078
rect 16028 28620 16080 28626
rect 16028 28562 16080 28568
rect 16040 28082 16068 28562
rect 16592 28490 16620 36502
rect 17420 36242 17448 36518
rect 17408 36236 17460 36242
rect 17408 36178 17460 36184
rect 18340 36174 18368 38354
rect 18696 37868 18748 37874
rect 18696 37810 18748 37816
rect 18604 36712 18656 36718
rect 18604 36654 18656 36660
rect 18616 36582 18644 36654
rect 18420 36576 18472 36582
rect 18420 36518 18472 36524
rect 18604 36576 18656 36582
rect 18604 36518 18656 36524
rect 17040 36168 17092 36174
rect 17040 36110 17092 36116
rect 18328 36168 18380 36174
rect 18328 36110 18380 36116
rect 17052 33998 17080 36110
rect 18328 35148 18380 35154
rect 18328 35090 18380 35096
rect 17684 34944 17736 34950
rect 17684 34886 17736 34892
rect 17696 34610 17724 34886
rect 17960 34672 18012 34678
rect 17960 34614 18012 34620
rect 17408 34604 17460 34610
rect 17408 34546 17460 34552
rect 17684 34604 17736 34610
rect 17684 34546 17736 34552
rect 17420 34202 17448 34546
rect 17868 34400 17920 34406
rect 17868 34342 17920 34348
rect 17408 34196 17460 34202
rect 17408 34138 17460 34144
rect 17040 33992 17092 33998
rect 17224 33992 17276 33998
rect 17040 33934 17092 33940
rect 17144 33952 17224 33980
rect 16948 33584 17000 33590
rect 16948 33526 17000 33532
rect 16960 33114 16988 33526
rect 16948 33108 17000 33114
rect 16948 33050 17000 33056
rect 16672 32904 16724 32910
rect 16672 32846 16724 32852
rect 16684 30666 16712 32846
rect 16948 32836 17000 32842
rect 16948 32778 17000 32784
rect 16764 31884 16816 31890
rect 16764 31826 16816 31832
rect 16776 31346 16804 31826
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 16672 30660 16724 30666
rect 16672 30602 16724 30608
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16684 28626 16712 29446
rect 16672 28620 16724 28626
rect 16672 28562 16724 28568
rect 16580 28484 16632 28490
rect 16580 28426 16632 28432
rect 16028 28076 16080 28082
rect 16028 28018 16080 28024
rect 14464 27950 14516 27956
rect 14188 27940 14424 27946
rect 14240 27934 14372 27940
rect 14188 27882 14240 27888
rect 14372 27882 14424 27888
rect 14476 27674 14504 27950
rect 15304 27934 15608 27962
rect 14464 27668 14516 27674
rect 14464 27610 14516 27616
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14188 27328 14240 27334
rect 14188 27270 14240 27276
rect 14200 27062 14228 27270
rect 14188 27056 14240 27062
rect 14188 26998 14240 27004
rect 14096 25764 14148 25770
rect 14096 25706 14148 25712
rect 14004 25220 14056 25226
rect 14004 25162 14056 25168
rect 14016 24206 14044 25162
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14108 24886 14136 25094
rect 14096 24880 14148 24886
rect 14096 24822 14148 24828
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 14016 23118 14044 24142
rect 14752 24070 14780 27406
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 15304 23594 15332 27934
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15660 25968 15712 25974
rect 15660 25910 15712 25916
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15580 25362 15608 25842
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15672 25294 15700 25910
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15488 24274 15516 24550
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15488 23798 15516 24210
rect 15476 23792 15528 23798
rect 15476 23734 15528 23740
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 15488 23254 15516 23734
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 14016 22234 14044 23054
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14384 22642 14412 22918
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14004 22228 14056 22234
rect 14004 22170 14056 22176
rect 14924 21956 14976 21962
rect 14924 21898 14976 21904
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14108 20346 14136 20878
rect 14752 20874 14780 21490
rect 14936 21146 14964 21898
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 14740 20868 14792 20874
rect 14740 20810 14792 20816
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 14200 20534 14228 20742
rect 14188 20528 14240 20534
rect 14188 20470 14240 20476
rect 13912 20324 13964 20330
rect 14108 20318 14228 20346
rect 13912 20266 13964 20272
rect 13924 19990 13952 20266
rect 14200 20262 14228 20318
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14108 19990 14136 20198
rect 13912 19984 13964 19990
rect 13912 19926 13964 19932
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 14016 19310 14044 19858
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13924 19122 13952 19178
rect 13924 19094 14044 19122
rect 14016 17882 14044 19094
rect 14292 18086 14320 19314
rect 14476 18290 14504 20198
rect 14936 20058 14964 21082
rect 15672 20874 15700 25230
rect 15764 24682 15792 26318
rect 15856 25158 15884 26930
rect 16120 26784 16172 26790
rect 16120 26726 16172 26732
rect 16132 26518 16160 26726
rect 16120 26512 16172 26518
rect 16120 26454 16172 26460
rect 16212 26308 16264 26314
rect 16212 26250 16264 26256
rect 15936 26240 15988 26246
rect 15936 26182 15988 26188
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15752 24676 15804 24682
rect 15752 24618 15804 24624
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 15764 23254 15792 24142
rect 15752 23248 15804 23254
rect 15752 23190 15804 23196
rect 15856 23118 15884 25094
rect 15948 23866 15976 26182
rect 16224 25770 16252 26250
rect 16396 26240 16448 26246
rect 16396 26182 16448 26188
rect 16408 26042 16436 26182
rect 16396 26036 16448 26042
rect 16396 25978 16448 25984
rect 16212 25764 16264 25770
rect 16212 25706 16264 25712
rect 16408 24206 16436 25978
rect 16580 25832 16632 25838
rect 16580 25774 16632 25780
rect 16592 25498 16620 25774
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 16580 25220 16632 25226
rect 16580 25162 16632 25168
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 16500 24206 16528 24618
rect 16592 24274 16620 25162
rect 16580 24268 16632 24274
rect 16580 24210 16632 24216
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15844 22976 15896 22982
rect 15948 22964 15976 23802
rect 16040 23322 16068 24142
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16316 23798 16344 24006
rect 16408 23866 16436 24142
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 16684 23730 16712 24006
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 15896 22936 15976 22964
rect 16028 22976 16080 22982
rect 15844 22918 15896 22924
rect 16028 22918 16080 22924
rect 15936 22568 15988 22574
rect 15936 22510 15988 22516
rect 15948 22098 15976 22510
rect 16040 22166 16068 22918
rect 16132 22778 16160 23598
rect 16672 23588 16724 23594
rect 16672 23530 16724 23536
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16592 23186 16620 23258
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16684 23118 16712 23530
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16580 23044 16632 23050
rect 16580 22986 16632 22992
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 16028 22160 16080 22166
rect 16028 22102 16080 22108
rect 15936 22092 15988 22098
rect 15936 22034 15988 22040
rect 16132 22030 16160 22714
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16592 21486 16620 22986
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 16684 21554 16712 22034
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 14740 19780 14792 19786
rect 14740 19722 14792 19728
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14568 19242 14596 19654
rect 14752 19446 14780 19722
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14556 19236 14608 19242
rect 14556 19178 14608 19184
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 13832 17734 13952 17762
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13832 16794 13860 17546
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 9876 15162 9904 15370
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 11072 15026 11100 16050
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13372 15094 13400 15506
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13360 15088 13412 15094
rect 13360 15030 13412 15036
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 13648 13938 13676 15438
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13832 14958 13860 15302
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13924 13818 13952 17734
rect 14016 16454 14044 17818
rect 14292 17610 14320 18022
rect 14280 17604 14332 17610
rect 14280 17546 14332 17552
rect 14292 16590 14320 17546
rect 14752 17542 14780 19382
rect 14832 18692 14884 18698
rect 14832 18634 14884 18640
rect 14844 18426 14872 18634
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14752 17134 14780 17478
rect 14844 17202 14872 18226
rect 15672 18222 15700 20810
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15856 17202 15884 20402
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15948 19922 15976 20198
rect 15936 19916 15988 19922
rect 15936 19858 15988 19864
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14752 16726 14780 17070
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 14016 15434 14044 16390
rect 14292 15570 14320 16526
rect 14752 16522 14780 16662
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14844 15502 14872 17138
rect 15856 17082 15884 17138
rect 15856 17054 15976 17082
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15856 16658 15884 16934
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14004 15428 14056 15434
rect 14004 15370 14056 15376
rect 14844 14414 14872 15438
rect 14924 15360 14976 15366
rect 14924 15302 14976 15308
rect 14936 15094 14964 15302
rect 14924 15088 14976 15094
rect 14924 15030 14976 15036
rect 15028 14414 15056 15506
rect 15120 14958 15148 16390
rect 15856 16182 15884 16458
rect 15844 16176 15896 16182
rect 15844 16118 15896 16124
rect 15948 15026 15976 17054
rect 16224 16182 16252 17614
rect 16212 16176 16264 16182
rect 16212 16118 16264 16124
rect 16224 15570 16252 16118
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 16132 15162 16160 15370
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 14006 14320 14214
rect 14476 14006 14504 14282
rect 15396 14278 15424 14350
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 15396 13852 15424 14214
rect 15948 13938 15976 14962
rect 16408 14618 16436 18294
rect 16592 17542 16620 18634
rect 16684 18426 16712 18702
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16672 18148 16724 18154
rect 16672 18090 16724 18096
rect 16684 17746 16712 18090
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16684 17066 16712 17682
rect 16672 17060 16724 17066
rect 16672 17002 16724 17008
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15476 13864 15528 13870
rect 15396 13824 15476 13852
rect 13832 13790 13952 13818
rect 15476 13806 15528 13812
rect 13832 13734 13860 13790
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 12452 8294 12480 13398
rect 15488 13258 15516 13806
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 13394 16068 13670
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 2514 6776 3334
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7116 800 7144 2450
rect 7484 2378 7512 3470
rect 7944 3058 7972 3470
rect 8128 3126 8156 3878
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 7760 800 7788 2926
rect 8404 800 8432 3402
rect 9140 2514 9168 3878
rect 10336 3602 10364 4558
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 3602 10548 3878
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10336 2514 10364 2790
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 9048 800 9076 2314
rect 10980 800 11008 3538
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13556 3058 13584 3470
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 3126 13768 3334
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14200 800 14228 2926
rect 14844 800 14872 11290
rect 15028 11218 15056 12174
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 11218 15240 11494
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15672 8974 15700 11698
rect 16592 9042 16620 16186
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16684 13938 16712 16050
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15672 4078 15700 8910
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 16684 4010 16712 8978
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15212 2582 15240 2926
rect 15488 2650 15516 3402
rect 16776 2774 16804 31078
rect 16960 30734 16988 32778
rect 17052 32502 17080 33934
rect 17040 32496 17092 32502
rect 17040 32438 17092 32444
rect 17144 32434 17172 33952
rect 17224 33934 17276 33940
rect 17420 33590 17448 34138
rect 17880 33946 17908 34342
rect 17972 34066 18000 34614
rect 18052 34468 18104 34474
rect 18052 34410 18104 34416
rect 17960 34060 18012 34066
rect 17960 34002 18012 34008
rect 18064 33998 18092 34410
rect 18144 34400 18196 34406
rect 18144 34342 18196 34348
rect 18052 33992 18104 33998
rect 17880 33918 18000 33946
rect 18052 33934 18104 33940
rect 17408 33584 17460 33590
rect 17408 33526 17460 33532
rect 17776 33516 17828 33522
rect 17776 33458 17828 33464
rect 17788 32910 17816 33458
rect 17684 32904 17736 32910
rect 17684 32846 17736 32852
rect 17776 32904 17828 32910
rect 17776 32846 17828 32852
rect 17132 32428 17184 32434
rect 17132 32370 17184 32376
rect 17144 32026 17172 32370
rect 17224 32224 17276 32230
rect 17224 32166 17276 32172
rect 17132 32020 17184 32026
rect 17132 31962 17184 31968
rect 17236 31890 17264 32166
rect 17224 31884 17276 31890
rect 17224 31826 17276 31832
rect 17408 31680 17460 31686
rect 17408 31622 17460 31628
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 17144 30938 17172 31282
rect 17132 30932 17184 30938
rect 17132 30874 17184 30880
rect 16856 30728 16908 30734
rect 16856 30670 16908 30676
rect 16948 30728 17000 30734
rect 16948 30670 17000 30676
rect 16868 29170 16896 30670
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 17328 29646 17356 30534
rect 17316 29640 17368 29646
rect 17316 29582 17368 29588
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 17420 28642 17448 31622
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17604 29306 17632 29582
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17328 28614 17448 28642
rect 17040 26240 17092 26246
rect 17040 26182 17092 26188
rect 17052 25974 17080 26182
rect 17040 25968 17092 25974
rect 17040 25910 17092 25916
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16868 22778 16896 22918
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17132 19780 17184 19786
rect 17132 19722 17184 19728
rect 16856 19236 16908 19242
rect 16856 19178 16908 19184
rect 16868 18290 16896 19178
rect 17144 18834 17172 19722
rect 17236 19446 17264 20198
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16960 17814 16988 18226
rect 17144 18154 17172 18770
rect 17236 18698 17264 19246
rect 17328 19242 17356 28614
rect 17408 28484 17460 28490
rect 17408 28426 17460 28432
rect 17420 27606 17448 28426
rect 17408 27600 17460 27606
rect 17408 27542 17460 27548
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 17604 22234 17632 22510
rect 17592 22228 17644 22234
rect 17592 22170 17644 22176
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17512 21690 17540 21966
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17420 19258 17448 21422
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17512 19378 17540 20198
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 17316 19236 17368 19242
rect 17420 19230 17540 19258
rect 17316 19178 17368 19184
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 17132 18148 17184 18154
rect 17132 18090 17184 18096
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 16960 17678 16988 17750
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16868 16114 16896 17546
rect 17328 17202 17356 17818
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17328 16998 17356 17138
rect 17420 17134 17448 18702
rect 17512 18630 17540 19230
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17512 18358 17540 18566
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17512 18086 17540 18294
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17512 17542 17540 18022
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17328 16250 17356 16934
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17420 16114 17448 17070
rect 17500 16516 17552 16522
rect 17500 16458 17552 16464
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17236 15094 17264 15846
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 16856 14544 16908 14550
rect 17144 14498 17172 14554
rect 16856 14486 16908 14492
rect 16868 14346 16896 14486
rect 16960 14470 17172 14498
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17224 14476 17276 14482
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16868 14006 16896 14282
rect 16960 14278 16988 14470
rect 17224 14418 17276 14424
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16960 13938 16988 14214
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 17052 13870 17080 14214
rect 17236 14074 17264 14418
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 16868 12306 16896 13806
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17144 12850 17172 13126
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17052 12374 17080 12718
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 17130 3496 17186 3505
rect 17130 3431 17132 3440
rect 17184 3431 17186 3440
rect 17132 3402 17184 3408
rect 16776 2746 16896 2774
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15488 800 15516 2382
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16132 800 16160 2314
rect 16868 2310 16896 2746
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 17420 800 17448 14486
rect 17512 3602 17540 16458
rect 17696 12434 17724 32846
rect 17868 32428 17920 32434
rect 17868 32370 17920 32376
rect 17880 31686 17908 32370
rect 17972 32298 18000 33918
rect 18156 33658 18184 34342
rect 18236 34196 18288 34202
rect 18236 34138 18288 34144
rect 18144 33652 18196 33658
rect 18144 33594 18196 33600
rect 18156 32910 18184 33594
rect 18144 32904 18196 32910
rect 18144 32846 18196 32852
rect 18052 32836 18104 32842
rect 18052 32778 18104 32784
rect 18064 32298 18092 32778
rect 18248 32434 18276 34138
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 17960 32292 18012 32298
rect 17960 32234 18012 32240
rect 18052 32292 18104 32298
rect 18052 32234 18104 32240
rect 17972 31890 18000 32234
rect 17960 31884 18012 31890
rect 17960 31826 18012 31832
rect 18248 31754 18276 32370
rect 18340 32026 18368 35090
rect 18432 34066 18460 36518
rect 18512 35012 18564 35018
rect 18512 34954 18564 34960
rect 18524 34746 18552 34954
rect 18512 34740 18564 34746
rect 18512 34682 18564 34688
rect 18524 34542 18552 34682
rect 18708 34610 18736 37810
rect 19064 36168 19116 36174
rect 19064 36110 19116 36116
rect 18880 35284 18932 35290
rect 18880 35226 18932 35232
rect 18696 34604 18748 34610
rect 18696 34546 18748 34552
rect 18512 34536 18564 34542
rect 18512 34478 18564 34484
rect 18420 34060 18472 34066
rect 18420 34002 18472 34008
rect 18696 33584 18748 33590
rect 18696 33526 18748 33532
rect 18708 33114 18736 33526
rect 18892 33454 18920 35226
rect 19076 34474 19104 36110
rect 19064 34468 19116 34474
rect 19064 34410 19116 34416
rect 18972 34060 19024 34066
rect 18972 34002 19024 34008
rect 18880 33448 18932 33454
rect 18880 33390 18932 33396
rect 18696 33108 18748 33114
rect 18696 33050 18748 33056
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 18328 32020 18380 32026
rect 18328 31962 18380 31968
rect 18524 31822 18552 32166
rect 18512 31816 18564 31822
rect 18512 31758 18564 31764
rect 17972 31726 18276 31754
rect 18328 31748 18380 31754
rect 17868 31680 17920 31686
rect 17868 31622 17920 31628
rect 17972 31210 18000 31726
rect 18328 31690 18380 31696
rect 18236 31680 18288 31686
rect 18236 31622 18288 31628
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 17960 31204 18012 31210
rect 17960 31146 18012 31152
rect 17972 30734 18000 31146
rect 18064 31142 18092 31214
rect 18052 31136 18104 31142
rect 18052 31078 18104 31084
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 17960 29164 18012 29170
rect 17960 29106 18012 29112
rect 17972 28762 18000 29106
rect 18064 29050 18092 31078
rect 18248 30734 18276 31622
rect 18340 31278 18368 31690
rect 18524 31346 18552 31758
rect 18892 31414 18920 33390
rect 18880 31408 18932 31414
rect 18880 31350 18932 31356
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18328 31272 18380 31278
rect 18328 31214 18380 31220
rect 18236 30728 18288 30734
rect 18236 30670 18288 30676
rect 18248 30190 18276 30670
rect 18236 30184 18288 30190
rect 18236 30126 18288 30132
rect 18236 29640 18288 29646
rect 18236 29582 18288 29588
rect 18248 29170 18276 29582
rect 18892 29510 18920 31350
rect 18984 30122 19012 34002
rect 19076 33998 19104 34410
rect 19064 33992 19116 33998
rect 19064 33934 19116 33940
rect 19168 31754 19196 41386
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19524 38752 19576 38758
rect 19524 38694 19576 38700
rect 19536 38282 19564 38694
rect 19524 38276 19576 38282
rect 19524 38218 19576 38224
rect 19248 38208 19300 38214
rect 19248 38150 19300 38156
rect 19260 37874 19288 38150
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19248 37868 19300 37874
rect 19248 37810 19300 37816
rect 19340 37732 19392 37738
rect 19340 37674 19392 37680
rect 19352 35170 19380 37674
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19984 36100 20036 36106
rect 19984 36042 20036 36048
rect 19432 36032 19484 36038
rect 19432 35974 19484 35980
rect 19444 35766 19472 35974
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19996 35766 20024 36042
rect 19432 35760 19484 35766
rect 19432 35702 19484 35708
rect 19984 35760 20036 35766
rect 19984 35702 20036 35708
rect 19352 35142 19472 35170
rect 19340 35012 19392 35018
rect 19340 34954 19392 34960
rect 19352 34610 19380 34954
rect 19340 34604 19392 34610
rect 19340 34546 19392 34552
rect 19340 33856 19392 33862
rect 19340 33798 19392 33804
rect 19352 33590 19380 33798
rect 19444 33658 19472 35142
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 19340 33584 19392 33590
rect 19340 33526 19392 33532
rect 19708 33516 19760 33522
rect 19708 33458 19760 33464
rect 19984 33516 20036 33522
rect 19984 33458 20036 33464
rect 19248 33108 19300 33114
rect 19248 33050 19300 33056
rect 19260 31754 19288 33050
rect 19720 32842 19748 33458
rect 19708 32836 19760 32842
rect 19708 32778 19760 32784
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19076 31726 19196 31754
rect 19248 31748 19300 31754
rect 18972 30116 19024 30122
rect 18972 30058 19024 30064
rect 18604 29504 18656 29510
rect 18604 29446 18656 29452
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 18616 29170 18644 29446
rect 18236 29164 18288 29170
rect 18236 29106 18288 29112
rect 18604 29164 18656 29170
rect 18604 29106 18656 29112
rect 19076 29050 19104 31726
rect 19248 31690 19300 31696
rect 19352 31278 19380 32710
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19996 32502 20024 33458
rect 19984 32496 20036 32502
rect 19984 32438 20036 32444
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19340 31272 19392 31278
rect 19340 31214 19392 31220
rect 19444 30054 19472 31758
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19996 30326 20024 32438
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 19432 30048 19484 30054
rect 19432 29990 19484 29996
rect 18064 29022 18276 29050
rect 18052 28960 18104 28966
rect 18052 28902 18104 28908
rect 17960 28756 18012 28762
rect 17960 28698 18012 28704
rect 18064 28150 18092 28902
rect 18052 28144 18104 28150
rect 18052 28086 18104 28092
rect 18248 26790 18276 29022
rect 18984 29022 19104 29050
rect 19156 29096 19208 29102
rect 19156 29038 19208 29044
rect 18512 28144 18564 28150
rect 18512 28086 18564 28092
rect 18524 27606 18552 28086
rect 18512 27600 18564 27606
rect 18512 27542 18564 27548
rect 18236 26784 18288 26790
rect 18236 26726 18288 26732
rect 17960 25968 18012 25974
rect 17960 25910 18012 25916
rect 17972 24818 18000 25910
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 17972 24206 18000 24618
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 17972 23866 18000 24142
rect 18052 24064 18104 24070
rect 18052 24006 18104 24012
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 18064 23730 18092 24006
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 18248 19854 18276 26726
rect 18880 26240 18932 26246
rect 18880 26182 18932 26188
rect 18892 25906 18920 26182
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 18892 25430 18920 25842
rect 18880 25424 18932 25430
rect 18880 25366 18932 25372
rect 18892 24818 18920 25366
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 18984 23050 19012 29022
rect 19064 28960 19116 28966
rect 19064 28902 19116 28908
rect 19076 28762 19104 28902
rect 19064 28756 19116 28762
rect 19064 28698 19116 28704
rect 19076 28150 19104 28698
rect 19064 28144 19116 28150
rect 19064 28086 19116 28092
rect 19168 28014 19196 29038
rect 19340 29028 19392 29034
rect 19340 28970 19392 28976
rect 19352 28762 19380 28970
rect 19340 28756 19392 28762
rect 19340 28698 19392 28704
rect 19444 28626 19472 29990
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19800 29232 19852 29238
rect 19800 29174 19852 29180
rect 19812 28762 19840 29174
rect 19800 28756 19852 28762
rect 19800 28698 19852 28704
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19444 28218 19472 28562
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19248 28212 19300 28218
rect 19248 28154 19300 28160
rect 19432 28212 19484 28218
rect 19432 28154 19484 28160
rect 19156 28008 19208 28014
rect 19156 27950 19208 27956
rect 19064 27464 19116 27470
rect 19064 27406 19116 27412
rect 19076 25770 19104 27406
rect 19064 25764 19116 25770
rect 19064 25706 19116 25712
rect 19260 25362 19288 28154
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19996 25770 20024 25842
rect 19984 25764 20036 25770
rect 19984 25706 20036 25712
rect 19524 25696 19576 25702
rect 19524 25638 19576 25644
rect 19536 25362 19564 25638
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19168 24154 19196 24550
rect 19260 24274 19288 25298
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19996 24818 20024 25706
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19248 24268 19300 24274
rect 19248 24210 19300 24216
rect 19168 24126 19288 24154
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18972 23044 19024 23050
rect 18972 22986 19024 22992
rect 18616 22710 18644 22986
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 18616 22094 18644 22646
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 18616 22066 18736 22094
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18432 20466 18460 20878
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 18616 20466 18644 20742
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18432 19990 18460 20402
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18420 19984 18472 19990
rect 18420 19926 18472 19932
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18064 18902 18092 19654
rect 18052 18896 18104 18902
rect 18052 18838 18104 18844
rect 18248 17626 18276 19790
rect 18340 18680 18368 19858
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18432 19310 18460 19790
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18432 18816 18460 19246
rect 18524 18970 18552 20334
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18432 18788 18552 18816
rect 18420 18692 18472 18698
rect 18340 18652 18420 18680
rect 18420 18634 18472 18640
rect 18432 18290 18460 18634
rect 18524 18290 18552 18788
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18432 17746 18460 18226
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18512 17672 18564 17678
rect 18248 17620 18512 17626
rect 18248 17614 18564 17620
rect 18248 17598 18552 17614
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18156 17202 18184 17478
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18052 16176 18104 16182
rect 18052 16118 18104 16124
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17604 12406 17724 12434
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17604 2582 17632 12406
rect 17788 6866 17816 15370
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 15162 18000 15302
rect 18064 15162 18092 16118
rect 18616 16114 18644 20402
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 18340 15026 18368 15846
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 17972 12238 18000 13942
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12850 18552 13126
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18524 4282 18552 4558
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 17696 3738 17724 4082
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 17972 2650 18000 3470
rect 18248 3194 18276 3470
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 18340 2446 18368 3334
rect 18524 2650 18552 4082
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18616 2446 18644 4966
rect 18708 2854 18736 22066
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 18984 21486 19012 21558
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18892 21146 18920 21422
rect 18880 21140 18932 21146
rect 18880 21082 18932 21088
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18800 19446 18828 20198
rect 18788 19440 18840 19446
rect 18788 19382 18840 19388
rect 18984 15706 19012 21422
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18892 12238 18920 12582
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18800 3058 18828 4422
rect 18892 3194 18920 5170
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18984 4146 19012 4558
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18880 3188 18932 3194
rect 18880 3130 18932 3136
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 19168 2774 19196 22510
rect 19260 20942 19288 24126
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19352 22778 19380 23598
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19260 19174 19288 19654
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19444 18850 19472 22986
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19996 22642 20024 24754
rect 19616 22636 19668 22642
rect 19616 22578 19668 22584
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 19628 22030 19656 22578
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 20088 20346 20116 45526
rect 20180 34066 20208 46922
rect 20260 38276 20312 38282
rect 20260 38218 20312 38224
rect 20272 38010 20300 38218
rect 20260 38004 20312 38010
rect 20260 37946 20312 37952
rect 20260 36168 20312 36174
rect 20260 36110 20312 36116
rect 20272 35222 20300 36110
rect 20260 35216 20312 35222
rect 20260 35158 20312 35164
rect 20168 34060 20220 34066
rect 20168 34002 20220 34008
rect 20260 33924 20312 33930
rect 20260 33866 20312 33872
rect 20168 32836 20220 32842
rect 20168 32778 20220 32784
rect 20180 32570 20208 32778
rect 20168 32564 20220 32570
rect 20168 32506 20220 32512
rect 20272 29646 20300 33866
rect 20364 31278 20392 46990
rect 20548 39098 20576 47058
rect 20640 46510 20668 49200
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 21284 46034 21312 49200
rect 25228 46368 25280 46374
rect 25228 46310 25280 46316
rect 25240 46034 25268 46310
rect 25424 46034 25452 49286
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49200 27150 50000
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49314 31014 50000
rect 30760 49286 31014 49314
rect 25792 46442 25820 49200
rect 25780 46436 25832 46442
rect 25780 46378 25832 46384
rect 27080 46034 27108 49200
rect 28368 47054 28396 49200
rect 29276 47252 29328 47258
rect 29276 47194 29328 47200
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 29288 46578 29316 47194
rect 29656 47054 29684 49200
rect 30760 47122 30788 49286
rect 30902 49200 31014 49286
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49200 40030 50000
rect 40562 49200 40674 50000
rect 41206 49314 41318 50000
rect 40788 49286 41318 49314
rect 30748 47116 30800 47122
rect 30748 47058 30800 47064
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 30104 47048 30156 47054
rect 30104 46990 30156 46996
rect 29920 46912 29972 46918
rect 29920 46854 29972 46860
rect 29276 46572 29328 46578
rect 29276 46514 29328 46520
rect 27620 46504 27672 46510
rect 27620 46446 27672 46452
rect 27632 46170 27660 46446
rect 27620 46164 27672 46170
rect 27620 46106 27672 46112
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 25228 46028 25280 46034
rect 25228 45970 25280 45976
rect 25412 46028 25464 46034
rect 25412 45970 25464 45976
rect 27068 46028 27120 46034
rect 27068 45970 27120 45976
rect 27620 46028 27672 46034
rect 27620 45970 27672 45976
rect 20904 45960 20956 45966
rect 20904 45902 20956 45908
rect 20916 45490 20944 45902
rect 21088 45892 21140 45898
rect 21088 45834 21140 45840
rect 25412 45892 25464 45898
rect 25412 45834 25464 45840
rect 20996 45824 21048 45830
rect 20996 45766 21048 45772
rect 20904 45484 20956 45490
rect 20904 45426 20956 45432
rect 20536 39092 20588 39098
rect 20536 39034 20588 39040
rect 20628 38888 20680 38894
rect 20628 38830 20680 38836
rect 20536 37868 20588 37874
rect 20536 37810 20588 37816
rect 20548 37618 20576 37810
rect 20640 37806 20668 38830
rect 21008 37874 21036 45766
rect 21100 45082 21128 45834
rect 21088 45076 21140 45082
rect 21088 45018 21140 45024
rect 25424 45014 25452 45834
rect 25780 45416 25832 45422
rect 25780 45358 25832 45364
rect 25412 45008 25464 45014
rect 25412 44950 25464 44956
rect 25792 44878 25820 45358
rect 21824 44872 21876 44878
rect 21824 44814 21876 44820
rect 25780 44872 25832 44878
rect 25780 44814 25832 44820
rect 21836 44402 21864 44814
rect 24676 44736 24728 44742
rect 24676 44678 24728 44684
rect 24688 44470 24716 44678
rect 24676 44464 24728 44470
rect 24676 44406 24728 44412
rect 21824 44396 21876 44402
rect 21824 44338 21876 44344
rect 21836 41414 21864 44338
rect 24492 44328 24544 44334
rect 24492 44270 24544 44276
rect 23480 43784 23532 43790
rect 23480 43726 23532 43732
rect 21652 41386 21864 41414
rect 21272 38412 21324 38418
rect 21272 38354 21324 38360
rect 20996 37868 21048 37874
rect 20996 37810 21048 37816
rect 21284 37806 21312 38354
rect 21548 37868 21600 37874
rect 21548 37810 21600 37816
rect 20628 37800 20680 37806
rect 20628 37742 20680 37748
rect 21272 37800 21324 37806
rect 21272 37742 21324 37748
rect 20548 37590 20668 37618
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20548 37126 20576 37198
rect 20536 37120 20588 37126
rect 20536 37062 20588 37068
rect 20536 36100 20588 36106
rect 20536 36042 20588 36048
rect 20548 35290 20576 36042
rect 20640 35834 20668 37590
rect 21284 37262 21312 37742
rect 21364 37664 21416 37670
rect 21364 37606 21416 37612
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 20628 35828 20680 35834
rect 20628 35770 20680 35776
rect 20720 35624 20772 35630
rect 20720 35566 20772 35572
rect 20536 35284 20588 35290
rect 20536 35226 20588 35232
rect 20732 34610 20760 35566
rect 20812 35488 20864 35494
rect 20812 35430 20864 35436
rect 20824 35086 20852 35430
rect 20916 35222 20944 37198
rect 21284 35630 21312 37198
rect 21272 35624 21324 35630
rect 21272 35566 21324 35572
rect 20904 35216 20956 35222
rect 20904 35158 20956 35164
rect 20996 35148 21048 35154
rect 20996 35090 21048 35096
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20904 34740 20956 34746
rect 20904 34682 20956 34688
rect 20720 34604 20772 34610
rect 20720 34546 20772 34552
rect 20732 33658 20760 34546
rect 20720 33652 20772 33658
rect 20720 33594 20772 33600
rect 20536 33516 20588 33522
rect 20536 33458 20588 33464
rect 20444 32768 20496 32774
rect 20444 32710 20496 32716
rect 20456 32434 20484 32710
rect 20548 32434 20576 33458
rect 20626 32464 20682 32473
rect 20444 32428 20496 32434
rect 20444 32370 20496 32376
rect 20536 32428 20588 32434
rect 20626 32399 20682 32408
rect 20536 32370 20588 32376
rect 20352 31272 20404 31278
rect 20352 31214 20404 31220
rect 20548 30326 20576 32370
rect 20640 32366 20668 32399
rect 20628 32360 20680 32366
rect 20628 32302 20680 32308
rect 20720 32360 20772 32366
rect 20720 32302 20772 32308
rect 20732 31754 20760 32302
rect 20732 31726 20852 31754
rect 20628 31340 20680 31346
rect 20628 31282 20680 31288
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20640 30870 20668 31282
rect 20628 30864 20680 30870
rect 20628 30806 20680 30812
rect 20732 30666 20760 31282
rect 20720 30660 20772 30666
rect 20720 30602 20772 30608
rect 20536 30320 20588 30326
rect 20536 30262 20588 30268
rect 20720 30320 20772 30326
rect 20720 30262 20772 30268
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20260 29640 20312 29646
rect 20260 29582 20312 29588
rect 20272 29238 20300 29582
rect 20260 29232 20312 29238
rect 20260 29174 20312 29180
rect 20364 28762 20392 30194
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20456 29646 20484 29990
rect 20444 29640 20496 29646
rect 20548 29628 20576 30262
rect 20732 29646 20760 30262
rect 20720 29640 20772 29646
rect 20548 29600 20668 29628
rect 20444 29582 20496 29588
rect 20456 29306 20484 29582
rect 20536 29504 20588 29510
rect 20536 29446 20588 29452
rect 20444 29300 20496 29306
rect 20444 29242 20496 29248
rect 20548 29170 20576 29446
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20352 28756 20404 28762
rect 20352 28698 20404 28704
rect 20364 27878 20392 28698
rect 20640 28082 20668 29600
rect 20720 29582 20772 29588
rect 20732 28558 20760 29582
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 20720 28416 20772 28422
rect 20720 28358 20772 28364
rect 20732 28218 20760 28358
rect 20720 28212 20772 28218
rect 20720 28154 20772 28160
rect 20536 28076 20588 28082
rect 20536 28018 20588 28024
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 20352 27872 20404 27878
rect 20352 27814 20404 27820
rect 20364 27674 20392 27814
rect 20352 27668 20404 27674
rect 20352 27610 20404 27616
rect 20260 26988 20312 26994
rect 20260 26930 20312 26936
rect 20272 26042 20300 26930
rect 20364 26874 20392 27610
rect 20548 27538 20576 28018
rect 20536 27532 20588 27538
rect 20536 27474 20588 27480
rect 20548 26994 20576 27474
rect 20824 27418 20852 31726
rect 20916 31142 20944 34682
rect 21008 34474 21036 35090
rect 21180 35080 21232 35086
rect 21180 35022 21232 35028
rect 20996 34468 21048 34474
rect 20996 34410 21048 34416
rect 21008 33862 21036 34410
rect 20996 33856 21048 33862
rect 20996 33798 21048 33804
rect 21088 33380 21140 33386
rect 21088 33322 21140 33328
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 21008 30938 21036 31282
rect 20996 30932 21048 30938
rect 20996 30874 21048 30880
rect 20994 30288 21050 30297
rect 20994 30223 21050 30232
rect 20904 28620 20956 28626
rect 20904 28562 20956 28568
rect 20916 27538 20944 28562
rect 20904 27532 20956 27538
rect 20904 27474 20956 27480
rect 20720 27396 20772 27402
rect 20824 27390 20944 27418
rect 20720 27338 20772 27344
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20364 26846 20484 26874
rect 20732 26858 20760 27338
rect 20812 26920 20864 26926
rect 20812 26862 20864 26868
rect 20456 26790 20484 26846
rect 20720 26852 20772 26858
rect 20720 26794 20772 26800
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 20824 26382 20852 26862
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20260 26036 20312 26042
rect 20260 25978 20312 25984
rect 20260 25696 20312 25702
rect 20260 25638 20312 25644
rect 20272 25226 20300 25638
rect 20260 25220 20312 25226
rect 20260 25162 20312 25168
rect 20352 24608 20404 24614
rect 20352 24550 20404 24556
rect 20364 24138 20392 24550
rect 20352 24132 20404 24138
rect 20352 24074 20404 24080
rect 20824 23662 20852 26318
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 20536 23112 20588 23118
rect 20534 23080 20536 23089
rect 20720 23112 20772 23118
rect 20588 23080 20590 23089
rect 20720 23054 20772 23060
rect 20534 23015 20590 23024
rect 20732 22438 20760 23054
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20180 21690 20208 21966
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20180 20942 20208 21626
rect 20272 21622 20300 22374
rect 20732 21978 20760 22374
rect 20824 22098 20852 23462
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20732 21962 20852 21978
rect 20732 21956 20864 21962
rect 20732 21950 20812 21956
rect 20812 21898 20864 21904
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20352 21072 20404 21078
rect 20352 21014 20404 21020
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20180 20466 20208 20878
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20088 20318 20208 20346
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19996 19718 20024 19790
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19260 18822 19472 18850
rect 19260 17762 19288 18822
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19352 18222 19380 18702
rect 19444 18426 19472 18702
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19352 17882 19380 18158
rect 19996 17882 20024 19654
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 20088 18426 20116 18634
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 19260 17734 19380 17762
rect 19352 16590 19380 17734
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19260 14414 19288 16050
rect 19352 15502 19380 16390
rect 19444 16250 19472 17206
rect 19996 16590 20024 17818
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 20180 16454 20208 20318
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20272 18290 20300 19926
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20272 17610 20300 18226
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19260 13462 19288 14350
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19352 13530 19380 14010
rect 19444 14006 19472 14214
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 19996 13326 20024 15438
rect 20364 15026 20392 21014
rect 20456 20942 20484 21286
rect 20444 20936 20496 20942
rect 20444 20878 20496 20884
rect 20456 19854 20484 20878
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20548 18970 20576 19314
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20536 18760 20588 18766
rect 20536 18702 20588 18708
rect 20548 18426 20576 18702
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20732 17746 20760 18022
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20824 17610 20852 19110
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 20272 14414 20300 14894
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20180 13394 20208 13670
rect 20732 13394 20760 14758
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19352 3534 19380 4490
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4146 19472 4422
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 20088 4282 20116 4558
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20076 3664 20128 3670
rect 20076 3606 20128 3612
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19076 2746 19196 2774
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18708 870 18920 898
rect 18708 800 18736 870
rect 3528 734 3740 762
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 18892 762 18920 870
rect 19076 762 19104 2746
rect 19352 800 19380 3130
rect 19996 3058 20024 3470
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 20088 1714 20116 3606
rect 20180 3602 20208 3878
rect 20536 3664 20588 3670
rect 20536 3606 20588 3612
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 20548 3194 20576 3606
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20640 2990 20668 5510
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20824 4826 20852 5170
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20732 3738 20760 4558
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20824 2990 20852 3334
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 20732 2514 20760 2790
rect 20916 2650 20944 27390
rect 21008 26246 21036 30223
rect 21100 27470 21128 33322
rect 21192 32434 21220 35022
rect 21272 33992 21324 33998
rect 21272 33934 21324 33940
rect 21284 33658 21312 33934
rect 21272 33652 21324 33658
rect 21272 33594 21324 33600
rect 21376 33538 21404 37606
rect 21560 36786 21588 37810
rect 21548 36780 21600 36786
rect 21548 36722 21600 36728
rect 21456 33992 21508 33998
rect 21454 33960 21456 33969
rect 21508 33960 21510 33969
rect 21454 33895 21510 33904
rect 21284 33510 21404 33538
rect 21180 32428 21232 32434
rect 21180 32370 21232 32376
rect 21180 31680 21232 31686
rect 21180 31622 21232 31628
rect 21192 30734 21220 31622
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 21284 30598 21312 33510
rect 21364 32836 21416 32842
rect 21364 32778 21416 32784
rect 21376 32026 21404 32778
rect 21456 32292 21508 32298
rect 21456 32234 21508 32240
rect 21364 32020 21416 32026
rect 21364 31962 21416 31968
rect 21272 30592 21324 30598
rect 21272 30534 21324 30540
rect 21284 30433 21312 30534
rect 21270 30424 21326 30433
rect 21270 30359 21326 30368
rect 21376 30190 21404 31962
rect 21468 31754 21496 32234
rect 21456 31748 21508 31754
rect 21456 31690 21508 31696
rect 21560 30297 21588 36722
rect 21546 30288 21602 30297
rect 21546 30223 21602 30232
rect 21272 30184 21324 30190
rect 21272 30126 21324 30132
rect 21364 30184 21416 30190
rect 21364 30126 21416 30132
rect 21180 29572 21232 29578
rect 21180 29514 21232 29520
rect 21192 29170 21220 29514
rect 21284 29510 21312 30126
rect 21272 29504 21324 29510
rect 21272 29446 21324 29452
rect 21376 29170 21404 30126
rect 21548 30116 21600 30122
rect 21548 30058 21600 30064
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 21364 29164 21416 29170
rect 21364 29106 21416 29112
rect 21180 28960 21232 28966
rect 21180 28902 21232 28908
rect 21192 28626 21220 28902
rect 21180 28620 21232 28626
rect 21180 28562 21232 28568
rect 21560 27878 21588 30058
rect 21180 27872 21232 27878
rect 21180 27814 21232 27820
rect 21548 27872 21600 27878
rect 21548 27814 21600 27820
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 21100 26994 21128 27406
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 20996 26240 21048 26246
rect 20996 26182 21048 26188
rect 20996 25968 21048 25974
rect 20996 25910 21048 25916
rect 21008 25498 21036 25910
rect 20996 25492 21048 25498
rect 20996 25434 21048 25440
rect 21008 25294 21036 25434
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 20996 24336 21048 24342
rect 20996 24278 21048 24284
rect 21008 22642 21036 24278
rect 21192 23526 21220 27814
rect 21652 26874 21680 41386
rect 22008 38820 22060 38826
rect 22008 38762 22060 38768
rect 22020 37670 22048 38762
rect 23204 38344 23256 38350
rect 23204 38286 23256 38292
rect 23216 38010 23244 38286
rect 23296 38208 23348 38214
rect 23296 38150 23348 38156
rect 22376 38004 22428 38010
rect 22376 37946 22428 37952
rect 23204 38004 23256 38010
rect 23204 37946 23256 37952
rect 22284 37868 22336 37874
rect 22284 37810 22336 37816
rect 22008 37664 22060 37670
rect 22008 37606 22060 37612
rect 21916 36100 21968 36106
rect 21916 36042 21968 36048
rect 21824 33312 21876 33318
rect 21824 33254 21876 33260
rect 21732 32972 21784 32978
rect 21732 32914 21784 32920
rect 21744 32366 21772 32914
rect 21836 32910 21864 33254
rect 21824 32904 21876 32910
rect 21824 32846 21876 32852
rect 21732 32360 21784 32366
rect 21732 32302 21784 32308
rect 21824 32224 21876 32230
rect 21824 32166 21876 32172
rect 21732 32020 21784 32026
rect 21732 31962 21784 31968
rect 21744 31210 21772 31962
rect 21836 31890 21864 32166
rect 21824 31884 21876 31890
rect 21824 31826 21876 31832
rect 21732 31204 21784 31210
rect 21732 31146 21784 31152
rect 21928 30870 21956 36042
rect 22100 34536 22152 34542
rect 22100 34478 22152 34484
rect 22112 34202 22140 34478
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 22296 33998 22324 37810
rect 22388 35086 22416 37946
rect 23308 37942 23336 38150
rect 23296 37936 23348 37942
rect 23296 37878 23348 37884
rect 22652 37256 22704 37262
rect 22652 37198 22704 37204
rect 22664 36922 22692 37198
rect 22928 37120 22980 37126
rect 22928 37062 22980 37068
rect 23112 37120 23164 37126
rect 23112 37062 23164 37068
rect 22940 36922 22968 37062
rect 22652 36916 22704 36922
rect 22652 36858 22704 36864
rect 22928 36916 22980 36922
rect 22928 36858 22980 36864
rect 23124 36786 23152 37062
rect 23388 36916 23440 36922
rect 23388 36858 23440 36864
rect 23112 36780 23164 36786
rect 23112 36722 23164 36728
rect 22560 36304 22612 36310
rect 22558 36272 22560 36281
rect 22612 36272 22614 36281
rect 23124 36242 23152 36722
rect 23400 36582 23428 36858
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 23386 36408 23442 36417
rect 23386 36343 23442 36352
rect 22558 36207 22614 36216
rect 23112 36236 23164 36242
rect 23112 36178 23164 36184
rect 23400 36038 23428 36343
rect 23492 36156 23520 43726
rect 23756 38752 23808 38758
rect 23756 38694 23808 38700
rect 23768 37806 23796 38694
rect 23940 38412 23992 38418
rect 23940 38354 23992 38360
rect 23756 37800 23808 37806
rect 23756 37742 23808 37748
rect 23952 36718 23980 38354
rect 23664 36712 23716 36718
rect 23940 36712 23992 36718
rect 23716 36660 23888 36666
rect 23664 36654 23888 36660
rect 23992 36660 24164 36666
rect 23940 36654 24164 36660
rect 23676 36638 23888 36654
rect 23952 36638 24164 36654
rect 23572 36576 23624 36582
rect 23572 36518 23624 36524
rect 23584 36394 23612 36518
rect 23584 36378 23704 36394
rect 23584 36372 23716 36378
rect 23584 36366 23664 36372
rect 23664 36314 23716 36320
rect 23572 36304 23624 36310
rect 23624 36252 23704 36258
rect 23572 36246 23704 36252
rect 23584 36230 23704 36246
rect 23572 36168 23624 36174
rect 23492 36128 23572 36156
rect 23572 36110 23624 36116
rect 23388 36032 23440 36038
rect 23388 35974 23440 35980
rect 22376 35080 22428 35086
rect 22376 35022 22428 35028
rect 22284 33992 22336 33998
rect 22284 33934 22336 33940
rect 22284 33040 22336 33046
rect 22284 32982 22336 32988
rect 22192 32768 22244 32774
rect 22192 32710 22244 32716
rect 22204 31822 22232 32710
rect 22296 32337 22324 32982
rect 22388 32434 22416 35022
rect 22652 35012 22704 35018
rect 22652 34954 22704 34960
rect 22560 34944 22612 34950
rect 22560 34886 22612 34892
rect 22572 34678 22600 34886
rect 22560 34672 22612 34678
rect 22560 34614 22612 34620
rect 22664 34241 22692 34954
rect 23584 34746 23612 36110
rect 23572 34740 23624 34746
rect 23572 34682 23624 34688
rect 23572 34400 23624 34406
rect 23572 34342 23624 34348
rect 22650 34232 22706 34241
rect 22650 34167 22652 34176
rect 22704 34167 22706 34176
rect 22652 34138 22704 34144
rect 23584 33998 23612 34342
rect 22744 33992 22796 33998
rect 22744 33934 22796 33940
rect 23572 33992 23624 33998
rect 23572 33934 23624 33940
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22560 33856 22612 33862
rect 22560 33798 22612 33804
rect 22480 33658 22508 33798
rect 22468 33652 22520 33658
rect 22468 33594 22520 33600
rect 22480 33114 22508 33594
rect 22572 33318 22600 33798
rect 22560 33312 22612 33318
rect 22560 33254 22612 33260
rect 22468 33108 22520 33114
rect 22468 33050 22520 33056
rect 22560 32904 22612 32910
rect 22560 32846 22612 32852
rect 22572 32570 22600 32846
rect 22756 32774 22784 33934
rect 23584 33522 23612 33934
rect 23572 33516 23624 33522
rect 23572 33458 23624 33464
rect 23388 33448 23440 33454
rect 23676 33402 23704 36230
rect 23756 36032 23808 36038
rect 23756 35974 23808 35980
rect 23768 35766 23796 35974
rect 23756 35760 23808 35766
rect 23756 35702 23808 35708
rect 23440 33396 23704 33402
rect 23388 33390 23704 33396
rect 23400 33374 23704 33390
rect 22744 32768 22796 32774
rect 22744 32710 22796 32716
rect 22560 32564 22612 32570
rect 22560 32506 22612 32512
rect 22376 32428 22428 32434
rect 22376 32370 22428 32376
rect 22282 32328 22338 32337
rect 22282 32263 22338 32272
rect 22192 31816 22244 31822
rect 22192 31758 22244 31764
rect 22100 31748 22152 31754
rect 22100 31690 22152 31696
rect 22008 31408 22060 31414
rect 22112 31362 22140 31690
rect 22060 31356 22140 31362
rect 22008 31350 22140 31356
rect 22020 31334 22140 31350
rect 21916 30864 21968 30870
rect 21916 30806 21968 30812
rect 22112 30802 22140 31334
rect 22100 30796 22152 30802
rect 22100 30738 22152 30744
rect 22388 30734 22416 32370
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 22376 30728 22428 30734
rect 22376 30670 22428 30676
rect 21928 30326 21956 30670
rect 22008 30660 22060 30666
rect 22008 30602 22060 30608
rect 21916 30320 21968 30326
rect 21916 30262 21968 30268
rect 21928 29850 21956 30262
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 22020 29646 22048 30602
rect 22190 30424 22246 30433
rect 22190 30359 22246 30368
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 21732 29028 21784 29034
rect 21732 28970 21784 28976
rect 21824 29028 21876 29034
rect 21824 28970 21876 28976
rect 21272 26852 21324 26858
rect 21272 26794 21324 26800
rect 21560 26846 21680 26874
rect 21284 26042 21312 26794
rect 21456 26376 21508 26382
rect 21456 26318 21508 26324
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 21468 25906 21496 26318
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 21362 23216 21418 23225
rect 21362 23151 21364 23160
rect 21416 23151 21418 23160
rect 21364 23122 21416 23128
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 21008 21622 21036 22578
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 20996 21616 21048 21622
rect 20996 21558 21048 21564
rect 21100 20942 21128 21898
rect 21560 21894 21588 26846
rect 21640 26376 21692 26382
rect 21640 26318 21692 26324
rect 21652 25498 21680 26318
rect 21640 25492 21692 25498
rect 21640 25434 21692 25440
rect 21744 22094 21772 28970
rect 21836 28762 21864 28970
rect 22020 28966 22048 29582
rect 22100 29572 22152 29578
rect 22100 29514 22152 29520
rect 22112 29170 22140 29514
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22008 28960 22060 28966
rect 22008 28902 22060 28908
rect 21824 28756 21876 28762
rect 21824 28698 21876 28704
rect 21916 28212 21968 28218
rect 21916 28154 21968 28160
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 21836 27606 21864 28018
rect 21824 27600 21876 27606
rect 21824 27542 21876 27548
rect 21836 27062 21864 27542
rect 21824 27056 21876 27062
rect 21824 26998 21876 27004
rect 21928 26518 21956 28154
rect 21916 26512 21968 26518
rect 21916 26454 21968 26460
rect 21824 26376 21876 26382
rect 21824 26318 21876 26324
rect 21836 25974 21864 26318
rect 21928 26058 21956 26454
rect 22204 26246 22232 30359
rect 22388 29646 22416 30670
rect 22572 30122 22600 32506
rect 22756 32230 22784 32710
rect 23204 32496 23256 32502
rect 23204 32438 23256 32444
rect 23216 32298 23244 32438
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23204 32292 23256 32298
rect 23204 32234 23256 32240
rect 22744 32224 22796 32230
rect 22744 32166 22796 32172
rect 23216 31822 23244 32234
rect 23400 32026 23428 32370
rect 23572 32224 23624 32230
rect 23572 32166 23624 32172
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 23204 31816 23256 31822
rect 23204 31758 23256 31764
rect 22744 31408 22796 31414
rect 22744 31350 22796 31356
rect 22756 30938 22784 31350
rect 22744 30932 22796 30938
rect 22744 30874 22796 30880
rect 23112 30864 23164 30870
rect 23112 30806 23164 30812
rect 22560 30116 22612 30122
rect 22560 30058 22612 30064
rect 22376 29640 22428 29646
rect 22376 29582 22428 29588
rect 22560 29504 22612 29510
rect 22560 29446 22612 29452
rect 22572 28490 22600 29446
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22664 28762 22692 29106
rect 22652 28756 22704 28762
rect 22652 28698 22704 28704
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22928 28416 22980 28422
rect 22928 28358 22980 28364
rect 22652 28212 22704 28218
rect 22652 28154 22704 28160
rect 22284 26308 22336 26314
rect 22284 26250 22336 26256
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 21928 26030 22048 26058
rect 21824 25968 21876 25974
rect 21824 25910 21876 25916
rect 21916 25900 21968 25906
rect 21916 25842 21968 25848
rect 21928 25294 21956 25842
rect 22020 25430 22048 26030
rect 22204 25786 22232 26182
rect 22296 26042 22324 26250
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22376 26036 22428 26042
rect 22376 25978 22428 25984
rect 22284 25832 22336 25838
rect 22204 25780 22284 25786
rect 22204 25774 22336 25780
rect 22204 25758 22324 25774
rect 22008 25424 22060 25430
rect 22008 25366 22060 25372
rect 22192 25424 22244 25430
rect 22192 25366 22244 25372
rect 21916 25288 21968 25294
rect 21916 25230 21968 25236
rect 21928 24410 21956 25230
rect 22204 24818 22232 25366
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 21916 24404 21968 24410
rect 21916 24346 21968 24352
rect 22020 24274 22048 24550
rect 22008 24268 22060 24274
rect 22008 24210 22060 24216
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22296 23866 22324 24006
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22112 23032 22140 23666
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22296 23186 22324 23462
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22192 23044 22244 23050
rect 22112 23004 22192 23032
rect 21744 22066 21956 22094
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21192 20534 21220 20742
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21180 20528 21232 20534
rect 21180 20470 21232 20476
rect 21192 19854 21220 20470
rect 21376 20398 21404 20538
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21008 16658 21036 16730
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 21008 12434 21036 16594
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21192 14278 21220 14758
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21008 12406 21220 12434
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 21008 2446 21036 3538
rect 21100 2582 21128 5646
rect 21192 2650 21220 12406
rect 21376 11762 21404 20334
rect 21560 12850 21588 21830
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21836 18970 21864 19790
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 21732 12844 21784 12850
rect 21732 12786 21784 12792
rect 21744 12434 21772 12786
rect 21652 12406 21772 12434
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21652 10674 21680 12406
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21744 11150 21772 11290
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21376 4622 21404 4966
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21652 4146 21680 10610
rect 21836 8294 21864 14418
rect 21928 12434 21956 22066
rect 22112 20534 22140 23004
rect 22192 22986 22244 22992
rect 22388 21486 22416 25978
rect 22664 25226 22692 28154
rect 22940 28082 22968 28358
rect 23124 28218 23152 30806
rect 23112 28212 23164 28218
rect 23112 28154 23164 28160
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22756 27674 22784 27814
rect 22744 27668 22796 27674
rect 22744 27610 22796 27616
rect 23400 27606 23428 31962
rect 23480 31680 23532 31686
rect 23480 31622 23532 31628
rect 23492 28626 23520 31622
rect 23584 31226 23612 32166
rect 23676 31754 23704 33374
rect 23768 32774 23796 35702
rect 23860 33046 23888 36638
rect 23940 36576 23992 36582
rect 23940 36518 23992 36524
rect 23952 36417 23980 36518
rect 23938 36408 23994 36417
rect 23938 36343 23994 36352
rect 24136 35834 24164 36638
rect 24124 35828 24176 35834
rect 24124 35770 24176 35776
rect 23940 35488 23992 35494
rect 23940 35430 23992 35436
rect 23848 33040 23900 33046
rect 23848 32982 23900 32988
rect 23952 32910 23980 35430
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24412 33386 24440 33934
rect 24400 33380 24452 33386
rect 24400 33322 24452 33328
rect 24308 32972 24360 32978
rect 24308 32914 24360 32920
rect 23940 32904 23992 32910
rect 23992 32864 24072 32892
rect 23940 32846 23992 32852
rect 23756 32768 23808 32774
rect 23756 32710 23808 32716
rect 24044 31822 24072 32864
rect 24320 32570 24348 32914
rect 24308 32564 24360 32570
rect 24308 32506 24360 32512
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 24032 31816 24084 31822
rect 24032 31758 24084 31764
rect 23676 31726 23888 31754
rect 23584 31198 23704 31226
rect 23572 31136 23624 31142
rect 23572 31078 23624 31084
rect 23584 30666 23612 31078
rect 23572 30660 23624 30666
rect 23572 30602 23624 30608
rect 23676 29646 23704 31198
rect 23860 30326 23888 31726
rect 23848 30320 23900 30326
rect 23848 30262 23900 30268
rect 23860 30054 23888 30262
rect 23848 30048 23900 30054
rect 23848 29990 23900 29996
rect 23664 29640 23716 29646
rect 23664 29582 23716 29588
rect 23480 28620 23532 28626
rect 23480 28562 23532 28568
rect 23676 28490 23704 29582
rect 23860 29102 23888 29990
rect 23848 29096 23900 29102
rect 23848 29038 23900 29044
rect 23756 28620 23808 28626
rect 23756 28562 23808 28568
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 23388 27600 23440 27606
rect 23388 27542 23440 27548
rect 23204 26376 23256 26382
rect 23204 26318 23256 26324
rect 22836 26240 22888 26246
rect 22836 26182 22888 26188
rect 22848 25226 22876 26182
rect 23216 25906 23244 26318
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23204 25900 23256 25906
rect 23204 25842 23256 25848
rect 22652 25220 22704 25226
rect 22652 25162 22704 25168
rect 22836 25220 22888 25226
rect 22836 25162 22888 25168
rect 22664 24954 22692 25162
rect 22652 24948 22704 24954
rect 22652 24890 22704 24896
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22204 19378 22232 20810
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22296 19514 22324 20334
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22204 18766 22232 19314
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22008 16516 22060 16522
rect 22008 16458 22060 16464
rect 22020 15706 22048 16458
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 22020 15026 22048 15642
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22112 15026 22140 15438
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 21928 12406 22048 12434
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21928 10810 21956 11018
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 22020 10690 22048 12406
rect 21928 10662 22048 10690
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 21836 4146 21864 4422
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 21928 4049 21956 10662
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 21914 4040 21970 4049
rect 21914 3975 21970 3984
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21376 3058 21404 3878
rect 22020 3194 22048 4558
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22112 3126 22140 14962
rect 22296 14346 22324 19246
rect 22284 14340 22336 14346
rect 22284 14282 22336 14288
rect 22296 13870 22324 14282
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22388 6798 22416 19722
rect 22480 16574 22508 24754
rect 22836 24676 22888 24682
rect 22836 24618 22888 24624
rect 22848 22642 22876 24618
rect 23020 23656 23072 23662
rect 23020 23598 23072 23604
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22940 23322 22968 23462
rect 22928 23316 22980 23322
rect 22928 23258 22980 23264
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 22572 22166 22600 22510
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 22560 22160 22612 22166
rect 22612 22108 22692 22114
rect 22560 22102 22692 22108
rect 22572 22086 22692 22102
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22572 19310 22600 21422
rect 22664 19786 22692 22086
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22848 19174 22876 22170
rect 23032 21146 23060 23598
rect 23020 21140 23072 21146
rect 23020 21082 23072 21088
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 23032 18970 23060 19246
rect 23020 18964 23072 18970
rect 23020 18906 23072 18912
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22664 18426 22692 18634
rect 22652 18420 22704 18426
rect 22652 18362 22704 18368
rect 22928 18352 22980 18358
rect 22928 18294 22980 18300
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22756 17610 22784 18022
rect 22940 17610 22968 18294
rect 22744 17604 22796 17610
rect 22744 17546 22796 17552
rect 22928 17604 22980 17610
rect 22928 17546 22980 17552
rect 22480 16546 22692 16574
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22376 5228 22428 5234
rect 22376 5170 22428 5176
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22204 3194 22232 3946
rect 22388 3670 22416 5170
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22480 4622 22508 4966
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 22376 3664 22428 3670
rect 22376 3606 22428 3612
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 22572 3058 22600 3470
rect 22664 3466 22692 16546
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 22928 14612 22980 14618
rect 22928 14554 22980 14560
rect 22940 14482 22968 14554
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22940 13938 22968 14418
rect 23032 14414 23060 14758
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22756 4826 22784 5170
rect 22744 4820 22796 4826
rect 22744 4762 22796 4768
rect 22848 4010 22876 13806
rect 22836 4004 22888 4010
rect 22836 3946 22888 3952
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 22652 3460 22704 3466
rect 22652 3402 22704 3408
rect 22756 3126 22784 3878
rect 23124 3738 23152 25842
rect 23216 22438 23244 25842
rect 23400 24682 23428 27542
rect 23768 27538 23796 28562
rect 23756 27532 23808 27538
rect 23756 27474 23808 27480
rect 23664 27396 23716 27402
rect 23664 27338 23716 27344
rect 23676 26586 23704 27338
rect 24044 27062 24072 31758
rect 24228 31686 24256 32370
rect 24504 31754 24532 44270
rect 24584 44192 24636 44198
rect 24584 44134 24636 44140
rect 24596 43858 24624 44134
rect 24584 43852 24636 43858
rect 24584 43794 24636 43800
rect 25792 41614 25820 44814
rect 27632 41682 27660 45970
rect 27620 41676 27672 41682
rect 27620 41618 27672 41624
rect 25780 41608 25832 41614
rect 25780 41550 25832 41556
rect 26424 41608 26476 41614
rect 26424 41550 26476 41556
rect 26436 40662 26464 41550
rect 29932 41414 29960 46854
rect 29840 41386 29960 41414
rect 26424 40656 26476 40662
rect 26424 40598 26476 40604
rect 27436 40452 27488 40458
rect 27436 40394 27488 40400
rect 25044 38888 25096 38894
rect 25044 38830 25096 38836
rect 25056 38554 25084 38830
rect 25044 38548 25096 38554
rect 25044 38490 25096 38496
rect 24676 38276 24728 38282
rect 24676 38218 24728 38224
rect 24688 37670 24716 38218
rect 24676 37664 24728 37670
rect 24676 37606 24728 37612
rect 24688 34610 24716 37606
rect 25780 37188 25832 37194
rect 25780 37130 25832 37136
rect 27068 37188 27120 37194
rect 27068 37130 27120 37136
rect 25792 36922 25820 37130
rect 27080 36922 27108 37130
rect 27252 37120 27304 37126
rect 27252 37062 27304 37068
rect 25320 36916 25372 36922
rect 25320 36858 25372 36864
rect 25780 36916 25832 36922
rect 25780 36858 25832 36864
rect 27068 36916 27120 36922
rect 27068 36858 27120 36864
rect 24860 36780 24912 36786
rect 24860 36722 24912 36728
rect 24952 36780 25004 36786
rect 24952 36722 25004 36728
rect 24872 36174 24900 36722
rect 24860 36168 24912 36174
rect 24860 36110 24912 36116
rect 24768 36032 24820 36038
rect 24768 35974 24820 35980
rect 24780 35698 24808 35974
rect 24768 35692 24820 35698
rect 24768 35634 24820 35640
rect 24780 34678 24808 35634
rect 24872 35630 24900 36110
rect 24964 36106 24992 36722
rect 25044 36644 25096 36650
rect 25044 36586 25096 36592
rect 25056 36242 25084 36586
rect 25044 36236 25096 36242
rect 25044 36178 25096 36184
rect 24952 36100 25004 36106
rect 24952 36042 25004 36048
rect 24860 35624 24912 35630
rect 24860 35566 24912 35572
rect 24872 34746 24900 35566
rect 25228 35012 25280 35018
rect 25228 34954 25280 34960
rect 24860 34740 24912 34746
rect 24860 34682 24912 34688
rect 25044 34740 25096 34746
rect 25044 34682 25096 34688
rect 24768 34672 24820 34678
rect 24768 34614 24820 34620
rect 24676 34604 24728 34610
rect 24676 34546 24728 34552
rect 24860 34400 24912 34406
rect 24860 34342 24912 34348
rect 24872 34202 24900 34342
rect 24860 34196 24912 34202
rect 24860 34138 24912 34144
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 24676 33856 24728 33862
rect 24676 33798 24728 33804
rect 24584 32768 24636 32774
rect 24584 32710 24636 32716
rect 24596 31822 24624 32710
rect 24584 31816 24636 31822
rect 24584 31758 24636 31764
rect 24320 31726 24532 31754
rect 24216 31680 24268 31686
rect 24216 31622 24268 31628
rect 24216 29776 24268 29782
rect 24216 29718 24268 29724
rect 24228 29510 24256 29718
rect 24216 29504 24268 29510
rect 24216 29446 24268 29452
rect 24228 28490 24256 29446
rect 24216 28484 24268 28490
rect 24216 28426 24268 28432
rect 24032 27056 24084 27062
rect 24032 26998 24084 27004
rect 23664 26580 23716 26586
rect 23664 26522 23716 26528
rect 23480 25356 23532 25362
rect 23480 25298 23532 25304
rect 23492 24818 23520 25298
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23768 24886 23796 25094
rect 23756 24880 23808 24886
rect 23756 24822 23808 24828
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23388 24676 23440 24682
rect 23388 24618 23440 24624
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 23676 23730 23704 24006
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23584 23050 23612 23462
rect 23572 23044 23624 23050
rect 23572 22986 23624 22992
rect 24216 22636 24268 22642
rect 24216 22578 24268 22584
rect 23204 22432 23256 22438
rect 23204 22374 23256 22380
rect 23216 18290 23244 22374
rect 23940 22092 23992 22098
rect 23940 22034 23992 22040
rect 23952 21554 23980 22034
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23400 20262 23428 20878
rect 24228 20466 24256 22578
rect 24320 22094 24348 31726
rect 24584 31476 24636 31482
rect 24584 31418 24636 31424
rect 24596 30258 24624 31418
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24400 28552 24452 28558
rect 24400 28494 24452 28500
rect 24412 28218 24440 28494
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24400 28212 24452 28218
rect 24400 28154 24452 28160
rect 24504 25294 24532 28358
rect 24596 26450 24624 30194
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 24492 23520 24544 23526
rect 24492 23462 24544 23468
rect 24504 23186 24532 23462
rect 24492 23180 24544 23186
rect 24492 23122 24544 23128
rect 24320 22066 24440 22094
rect 24412 20890 24440 22066
rect 24412 20862 24532 20890
rect 24400 20800 24452 20806
rect 24400 20742 24452 20748
rect 24412 20534 24440 20742
rect 24400 20528 24452 20534
rect 24400 20470 24452 20476
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 23400 19825 23428 19858
rect 24400 19848 24452 19854
rect 23386 19816 23442 19825
rect 24400 19790 24452 19796
rect 23386 19751 23442 19760
rect 24412 18970 24440 19790
rect 24400 18964 24452 18970
rect 24400 18906 24452 18912
rect 24400 18760 24452 18766
rect 24400 18702 24452 18708
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24228 18358 24256 18566
rect 24216 18352 24268 18358
rect 24216 18294 24268 18300
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 24412 17882 24440 18702
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24412 17270 24440 17818
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 24400 17264 24452 17270
rect 24400 17206 24452 17212
rect 23480 17060 23532 17066
rect 23480 17002 23532 17008
rect 23492 16590 23520 17002
rect 23676 16590 23704 17206
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23492 15570 23520 16526
rect 23480 15564 23532 15570
rect 23480 15506 23532 15512
rect 23676 15502 23704 16526
rect 23768 16522 23796 17070
rect 24504 16658 24532 20862
rect 24584 18216 24636 18222
rect 24584 18158 24636 18164
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 23756 16516 23808 16522
rect 23756 16458 23808 16464
rect 23768 16114 23796 16458
rect 24596 16182 24624 18158
rect 24584 16176 24636 16182
rect 24584 16118 24636 16124
rect 23756 16108 23808 16114
rect 23756 16050 23808 16056
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24412 15706 24440 16050
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23400 15094 23428 15302
rect 23768 15162 23796 15506
rect 23848 15428 23900 15434
rect 23848 15370 23900 15376
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23768 14346 23796 14962
rect 23756 14340 23808 14346
rect 23756 14282 23808 14288
rect 23768 14074 23796 14282
rect 23860 14278 23888 15370
rect 23952 15094 23980 15642
rect 24492 15156 24544 15162
rect 24492 15098 24544 15104
rect 23940 15088 23992 15094
rect 23940 15030 23992 15036
rect 24504 14618 24532 15098
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24032 14340 24084 14346
rect 24032 14282 24084 14288
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23860 12850 23888 14214
rect 24044 13938 24072 14282
rect 24504 13938 24532 14554
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23216 4622 23244 4966
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 21088 2576 21140 2582
rect 21088 2518 21140 2524
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 19996 1686 20116 1714
rect 19996 800 20024 1686
rect 20640 800 20668 2314
rect 21928 800 21956 2994
rect 22468 2984 22520 2990
rect 23032 2972 23060 3674
rect 23216 3534 23244 4422
rect 23388 3664 23440 3670
rect 23388 3606 23440 3612
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23112 2984 23164 2990
rect 23032 2944 23112 2972
rect 22468 2926 22520 2932
rect 23112 2926 23164 2932
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22112 2446 22140 2858
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22480 1578 22508 2926
rect 23400 2922 23428 3606
rect 23388 2916 23440 2922
rect 23388 2858 23440 2864
rect 23492 2802 23520 5170
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 23860 4146 23888 4422
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23952 3602 23980 3878
rect 23940 3596 23992 3602
rect 23940 3538 23992 3544
rect 23216 2774 23520 2802
rect 22480 1550 22600 1578
rect 22572 800 22600 1550
rect 23216 800 23244 2774
rect 24044 2378 24072 13874
rect 24596 13274 24624 16118
rect 24504 13246 24624 13274
rect 24504 4690 24532 13246
rect 24688 6914 24716 33798
rect 24780 33046 24808 33934
rect 24872 33674 24900 34138
rect 25056 34134 25084 34682
rect 25240 34202 25268 34954
rect 25332 34406 25360 36858
rect 25688 36848 25740 36854
rect 25688 36790 25740 36796
rect 25700 35698 25728 36790
rect 26148 36780 26200 36786
rect 26148 36722 26200 36728
rect 26056 36712 26108 36718
rect 26056 36654 26108 36660
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 25976 36378 26004 36518
rect 25780 36372 25832 36378
rect 25780 36314 25832 36320
rect 25964 36372 26016 36378
rect 25964 36314 26016 36320
rect 25792 36258 25820 36314
rect 25792 36230 25912 36258
rect 25884 36174 25912 36230
rect 26068 36174 26096 36654
rect 25872 36168 25924 36174
rect 25872 36110 25924 36116
rect 26056 36168 26108 36174
rect 26056 36110 26108 36116
rect 25688 35692 25740 35698
rect 25688 35634 25740 35640
rect 25964 35488 26016 35494
rect 25964 35430 26016 35436
rect 25976 35018 26004 35430
rect 25964 35012 26016 35018
rect 25964 34954 26016 34960
rect 25596 34944 25648 34950
rect 25596 34886 25648 34892
rect 25608 34610 25636 34886
rect 25596 34604 25648 34610
rect 25596 34546 25648 34552
rect 25412 34536 25464 34542
rect 25412 34478 25464 34484
rect 25320 34400 25372 34406
rect 25320 34342 25372 34348
rect 25228 34196 25280 34202
rect 25228 34138 25280 34144
rect 25044 34128 25096 34134
rect 25044 34070 25096 34076
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 24872 33646 24992 33674
rect 24964 33590 24992 33646
rect 24952 33584 25004 33590
rect 24952 33526 25004 33532
rect 24952 33312 25004 33318
rect 24952 33254 25004 33260
rect 24768 33040 24820 33046
rect 24768 32982 24820 32988
rect 24780 32774 24808 32982
rect 24768 32768 24820 32774
rect 24768 32710 24820 32716
rect 24964 32434 24992 33254
rect 25056 32473 25084 33934
rect 25332 33590 25360 34342
rect 25320 33584 25372 33590
rect 25320 33526 25372 33532
rect 25136 32836 25188 32842
rect 25136 32778 25188 32784
rect 25042 32464 25098 32473
rect 24952 32428 25004 32434
rect 25042 32399 25098 32408
rect 24952 32370 25004 32376
rect 24768 31884 24820 31890
rect 24768 31826 24820 31832
rect 24780 31482 24808 31826
rect 24860 31816 24912 31822
rect 24860 31758 24912 31764
rect 24768 31476 24820 31482
rect 24768 31418 24820 31424
rect 24768 31340 24820 31346
rect 24768 31282 24820 31288
rect 24780 24750 24808 31282
rect 24872 30802 24900 31758
rect 24860 30796 24912 30802
rect 24860 30738 24912 30744
rect 24964 29782 24992 32370
rect 25148 30734 25176 32778
rect 25332 32450 25360 33526
rect 25424 33454 25452 34478
rect 25608 34474 25636 34546
rect 25596 34468 25648 34474
rect 25596 34410 25648 34416
rect 25608 34066 25636 34410
rect 25596 34060 25648 34066
rect 25596 34002 25648 34008
rect 25964 33992 26016 33998
rect 25964 33934 26016 33940
rect 25976 33658 26004 33934
rect 25964 33652 26016 33658
rect 25964 33594 26016 33600
rect 25596 33516 25648 33522
rect 25596 33458 25648 33464
rect 25412 33448 25464 33454
rect 25412 33390 25464 33396
rect 25240 32422 25360 32450
rect 25240 32230 25268 32422
rect 25320 32360 25372 32366
rect 25608 32337 25636 33458
rect 26160 33114 26188 36722
rect 27264 36038 27292 37062
rect 27252 36032 27304 36038
rect 27252 35974 27304 35980
rect 27264 35850 27292 35974
rect 27172 35822 27292 35850
rect 26424 35760 26476 35766
rect 26424 35702 26476 35708
rect 26240 35012 26292 35018
rect 26240 34954 26292 34960
rect 26252 34241 26280 34954
rect 26238 34232 26294 34241
rect 26238 34167 26294 34176
rect 26148 33108 26200 33114
rect 26148 33050 26200 33056
rect 26436 32502 26464 35702
rect 26884 34740 26936 34746
rect 26884 34682 26936 34688
rect 26896 33998 26924 34682
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 26976 33992 27028 33998
rect 26976 33934 27028 33940
rect 26884 33448 26936 33454
rect 26884 33390 26936 33396
rect 26792 32972 26844 32978
rect 26792 32914 26844 32920
rect 26608 32904 26660 32910
rect 26608 32846 26660 32852
rect 26424 32496 26476 32502
rect 26424 32438 26476 32444
rect 26424 32360 26476 32366
rect 25320 32302 25372 32308
rect 25594 32328 25650 32337
rect 25228 32224 25280 32230
rect 25228 32166 25280 32172
rect 25332 31278 25360 32302
rect 26424 32302 26476 32308
rect 25594 32263 25650 32272
rect 25608 31958 25636 32263
rect 25688 32224 25740 32230
rect 25688 32166 25740 32172
rect 25596 31952 25648 31958
rect 25596 31894 25648 31900
rect 25320 31272 25372 31278
rect 25320 31214 25372 31220
rect 25136 30728 25188 30734
rect 25136 30670 25188 30676
rect 25148 30054 25176 30670
rect 25596 30320 25648 30326
rect 25596 30262 25648 30268
rect 25504 30252 25556 30258
rect 25504 30194 25556 30200
rect 25136 30048 25188 30054
rect 25136 29990 25188 29996
rect 24952 29776 25004 29782
rect 24952 29718 25004 29724
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24872 24818 24900 25638
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 24860 24812 24912 24818
rect 24860 24754 24912 24760
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24780 22030 24808 24142
rect 24872 23730 24900 24142
rect 24860 23724 24912 23730
rect 24860 23666 24912 23672
rect 24860 23044 24912 23050
rect 24860 22986 24912 22992
rect 24872 22574 24900 22986
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24780 20874 24808 21286
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24872 20806 24900 21490
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24872 18222 24900 18634
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24872 16590 24900 16934
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24872 15162 24900 15370
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24964 8362 24992 24346
rect 25056 12714 25084 25230
rect 25148 24410 25176 29990
rect 25516 29850 25544 30194
rect 25504 29844 25556 29850
rect 25504 29786 25556 29792
rect 25516 29170 25544 29786
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 25608 28994 25636 30262
rect 25700 29102 25728 32166
rect 26148 31816 26200 31822
rect 26148 31758 26200 31764
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 25792 30326 25820 31214
rect 26160 30394 26188 31758
rect 26436 31686 26464 32302
rect 26424 31680 26476 31686
rect 26424 31622 26476 31628
rect 26148 30388 26200 30394
rect 26148 30330 26200 30336
rect 25780 30320 25832 30326
rect 25780 30262 25832 30268
rect 26056 30184 26108 30190
rect 26056 30126 26108 30132
rect 25872 30048 25924 30054
rect 25872 29990 25924 29996
rect 25884 29646 25912 29990
rect 26068 29646 26096 30126
rect 26148 30116 26200 30122
rect 26148 30058 26200 30064
rect 26160 29850 26188 30058
rect 26148 29844 26200 29850
rect 26148 29786 26200 29792
rect 25872 29640 25924 29646
rect 25872 29582 25924 29588
rect 26056 29640 26108 29646
rect 26056 29582 26108 29588
rect 26148 29640 26200 29646
rect 26148 29582 26200 29588
rect 25688 29096 25740 29102
rect 25688 29038 25740 29044
rect 25608 28966 25912 28994
rect 25412 28960 25464 28966
rect 25412 28902 25464 28908
rect 25424 28762 25452 28902
rect 25412 28756 25464 28762
rect 25412 28698 25464 28704
rect 25780 28552 25832 28558
rect 25780 28494 25832 28500
rect 25228 28484 25280 28490
rect 25228 28426 25280 28432
rect 25240 28082 25268 28426
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25412 28076 25464 28082
rect 25412 28018 25464 28024
rect 25240 27878 25268 28018
rect 25228 27872 25280 27878
rect 25228 27814 25280 27820
rect 25240 24954 25268 27814
rect 25424 27538 25452 28018
rect 25596 28008 25648 28014
rect 25596 27950 25648 27956
rect 25412 27532 25464 27538
rect 25412 27474 25464 27480
rect 25608 27334 25636 27950
rect 25792 27946 25820 28494
rect 25884 28014 25912 28966
rect 26160 28218 26188 29582
rect 26424 29028 26476 29034
rect 26424 28970 26476 28976
rect 26436 28558 26464 28970
rect 26620 28558 26648 32846
rect 26700 31136 26752 31142
rect 26700 31078 26752 31084
rect 26712 30666 26740 31078
rect 26700 30660 26752 30666
rect 26700 30602 26752 30608
rect 26424 28552 26476 28558
rect 26424 28494 26476 28500
rect 26608 28552 26660 28558
rect 26608 28494 26660 28500
rect 26700 28552 26752 28558
rect 26700 28494 26752 28500
rect 26240 28416 26292 28422
rect 26240 28358 26292 28364
rect 26148 28212 26200 28218
rect 26148 28154 26200 28160
rect 25872 28008 25924 28014
rect 25872 27950 25924 27956
rect 25780 27940 25832 27946
rect 25780 27882 25832 27888
rect 25792 27470 25820 27882
rect 25884 27470 25912 27950
rect 25780 27464 25832 27470
rect 25780 27406 25832 27412
rect 25872 27464 25924 27470
rect 25872 27406 25924 27412
rect 25596 27328 25648 27334
rect 25596 27270 25648 27276
rect 25688 27328 25740 27334
rect 25688 27270 25740 27276
rect 25608 26926 25636 27270
rect 25700 26994 25728 27270
rect 26252 26994 26280 28358
rect 26516 27668 26568 27674
rect 26516 27610 26568 27616
rect 26528 27538 26556 27610
rect 26516 27532 26568 27538
rect 26516 27474 26568 27480
rect 26620 27062 26648 28494
rect 26712 28218 26740 28494
rect 26700 28212 26752 28218
rect 26700 28154 26752 28160
rect 26700 27464 26752 27470
rect 26700 27406 26752 27412
rect 26608 27056 26660 27062
rect 26608 26998 26660 27004
rect 25688 26988 25740 26994
rect 25688 26930 25740 26936
rect 26240 26988 26292 26994
rect 26240 26930 26292 26936
rect 25596 26920 25648 26926
rect 26056 26920 26108 26926
rect 25596 26862 25648 26868
rect 25976 26880 26056 26908
rect 25228 24948 25280 24954
rect 25228 24890 25280 24896
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 25516 22642 25544 24074
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 25596 23044 25648 23050
rect 25596 22986 25648 22992
rect 25608 22710 25636 22986
rect 25700 22710 25728 23666
rect 25596 22704 25648 22710
rect 25596 22646 25648 22652
rect 25688 22704 25740 22710
rect 25688 22646 25740 22652
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25700 22506 25728 22646
rect 25688 22500 25740 22506
rect 25688 22442 25740 22448
rect 25976 21350 26004 26880
rect 26056 26862 26108 26868
rect 26252 26518 26280 26930
rect 26712 26858 26740 27406
rect 26700 26852 26752 26858
rect 26700 26794 26752 26800
rect 26424 26784 26476 26790
rect 26424 26726 26476 26732
rect 26240 26512 26292 26518
rect 26240 26454 26292 26460
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 26068 25226 26096 25638
rect 26056 25220 26108 25226
rect 26056 25162 26108 25168
rect 26436 25158 26464 26726
rect 26712 25498 26740 26794
rect 26700 25492 26752 25498
rect 26700 25434 26752 25440
rect 26424 25152 26476 25158
rect 26424 25094 26476 25100
rect 26148 23724 26200 23730
rect 26148 23666 26200 23672
rect 26240 23724 26292 23730
rect 26240 23666 26292 23672
rect 26160 23118 26188 23666
rect 26252 23186 26280 23666
rect 26240 23180 26292 23186
rect 26240 23122 26292 23128
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 26252 23050 26280 23122
rect 26240 23044 26292 23050
rect 26240 22986 26292 22992
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 26344 22658 26372 22918
rect 26148 22636 26200 22642
rect 26068 22596 26148 22624
rect 26068 22506 26096 22596
rect 26148 22578 26200 22584
rect 26252 22630 26372 22658
rect 26252 22574 26280 22630
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26056 22500 26108 22506
rect 26056 22442 26108 22448
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 26620 22030 26648 22374
rect 26608 22024 26660 22030
rect 26608 21966 26660 21972
rect 26700 21548 26752 21554
rect 26700 21490 26752 21496
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25332 19922 25360 21286
rect 26712 21146 26740 21490
rect 26700 21140 26752 21146
rect 26700 21082 26752 21088
rect 26712 20942 26740 21082
rect 26700 20936 26752 20942
rect 26700 20878 26752 20884
rect 26148 20800 26200 20806
rect 26148 20742 26200 20748
rect 26056 20392 26108 20398
rect 26056 20334 26108 20340
rect 25780 20256 25832 20262
rect 25780 20198 25832 20204
rect 25792 19990 25820 20198
rect 25780 19984 25832 19990
rect 25780 19926 25832 19932
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25596 18828 25648 18834
rect 25596 18770 25648 18776
rect 25608 17746 25636 18770
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 25240 17338 25268 17614
rect 25228 17332 25280 17338
rect 25228 17274 25280 17280
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25228 14408 25280 14414
rect 25228 14350 25280 14356
rect 25240 14074 25268 14350
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 24952 8356 25004 8362
rect 24952 8298 25004 8304
rect 24596 6886 24716 6914
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 24492 3460 24544 3466
rect 24492 3402 24544 3408
rect 24032 2372 24084 2378
rect 24032 2314 24084 2320
rect 24504 800 24532 3402
rect 24596 3398 24624 6886
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24688 3126 24716 4966
rect 24952 4072 25004 4078
rect 24952 4014 25004 4020
rect 24860 4004 24912 4010
rect 24860 3946 24912 3952
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24676 3120 24728 3126
rect 24676 3062 24728 3068
rect 24780 2514 24808 3878
rect 24872 3534 24900 3946
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 24964 2650 24992 4014
rect 25424 3602 25452 16594
rect 25964 15088 26016 15094
rect 25964 15030 26016 15036
rect 25872 12776 25924 12782
rect 25872 12718 25924 12724
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25412 3596 25464 3602
rect 25412 3538 25464 3544
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 25516 2582 25544 3878
rect 25884 3738 25912 12718
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25608 2582 25636 3402
rect 25976 3126 26004 15030
rect 25964 3120 26016 3126
rect 25964 3062 26016 3068
rect 26068 2922 26096 20334
rect 26160 20058 26188 20742
rect 26148 20052 26200 20058
rect 26148 19994 26200 20000
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26252 17610 26280 18566
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 26148 15088 26200 15094
rect 26148 15030 26200 15036
rect 26160 14550 26188 15030
rect 26148 14544 26200 14550
rect 26148 14486 26200 14492
rect 26056 2916 26108 2922
rect 26056 2858 26108 2864
rect 26804 2650 26832 32914
rect 26896 32910 26924 33390
rect 26988 33386 27016 33934
rect 27068 33856 27120 33862
rect 27068 33798 27120 33804
rect 27080 33522 27108 33798
rect 27068 33516 27120 33522
rect 27068 33458 27120 33464
rect 26976 33380 27028 33386
rect 26976 33322 27028 33328
rect 26884 32904 26936 32910
rect 26884 32846 26936 32852
rect 27068 32904 27120 32910
rect 27172 32892 27200 35822
rect 27252 34944 27304 34950
rect 27252 34886 27304 34892
rect 27264 34134 27292 34886
rect 27252 34128 27304 34134
rect 27252 34070 27304 34076
rect 27252 33856 27304 33862
rect 27252 33798 27304 33804
rect 27264 33454 27292 33798
rect 27252 33448 27304 33454
rect 27252 33390 27304 33396
rect 27120 32864 27200 32892
rect 27252 32904 27304 32910
rect 27068 32846 27120 32852
rect 27252 32846 27304 32852
rect 27068 31204 27120 31210
rect 27068 31146 27120 31152
rect 27080 30938 27108 31146
rect 27068 30932 27120 30938
rect 27068 30874 27120 30880
rect 27080 29850 27108 30874
rect 27068 29844 27120 29850
rect 27068 29786 27120 29792
rect 26976 28076 27028 28082
rect 27080 28064 27108 29786
rect 27264 29034 27292 32846
rect 27344 32836 27396 32842
rect 27344 32778 27396 32784
rect 27356 30326 27384 32778
rect 27344 30320 27396 30326
rect 27344 30262 27396 30268
rect 27356 29646 27384 30262
rect 27344 29640 27396 29646
rect 27344 29582 27396 29588
rect 27252 29028 27304 29034
rect 27252 28970 27304 28976
rect 27264 28558 27292 28970
rect 27252 28552 27304 28558
rect 27252 28494 27304 28500
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 27264 28150 27292 28358
rect 27252 28144 27304 28150
rect 27252 28086 27304 28092
rect 27028 28036 27108 28064
rect 26976 28018 27028 28024
rect 26988 27674 27016 28018
rect 27448 27985 27476 40394
rect 28448 37256 28500 37262
rect 28448 37198 28500 37204
rect 27896 37188 27948 37194
rect 27896 37130 27948 37136
rect 27908 36786 27936 37130
rect 28460 36854 28488 37198
rect 28632 37120 28684 37126
rect 28632 37062 28684 37068
rect 28644 36854 28672 37062
rect 28448 36848 28500 36854
rect 28448 36790 28500 36796
rect 28632 36848 28684 36854
rect 28632 36790 28684 36796
rect 27896 36780 27948 36786
rect 27896 36722 27948 36728
rect 27712 36644 27764 36650
rect 27712 36586 27764 36592
rect 27724 35494 27752 36586
rect 27816 36310 27844 36341
rect 27804 36304 27856 36310
rect 27802 36272 27804 36281
rect 27856 36272 27858 36281
rect 27802 36207 27858 36216
rect 27816 36174 27844 36207
rect 27804 36168 27856 36174
rect 27804 36110 27856 36116
rect 27908 35766 27936 36722
rect 28172 36712 28224 36718
rect 28172 36654 28224 36660
rect 27988 36576 28040 36582
rect 27988 36518 28040 36524
rect 28000 36174 28028 36518
rect 28184 36378 28212 36654
rect 28172 36372 28224 36378
rect 28172 36314 28224 36320
rect 28460 36174 28488 36790
rect 28816 36576 28868 36582
rect 28816 36518 28868 36524
rect 27988 36168 28040 36174
rect 27988 36110 28040 36116
rect 28448 36168 28500 36174
rect 28448 36110 28500 36116
rect 28172 36100 28224 36106
rect 28172 36042 28224 36048
rect 28080 36032 28132 36038
rect 28080 35974 28132 35980
rect 27896 35760 27948 35766
rect 27896 35702 27948 35708
rect 27712 35488 27764 35494
rect 27712 35430 27764 35436
rect 27528 35284 27580 35290
rect 27528 35226 27580 35232
rect 27540 34066 27568 35226
rect 27908 35154 27936 35702
rect 27896 35148 27948 35154
rect 27896 35090 27948 35096
rect 27804 35080 27856 35086
rect 27804 35022 27856 35028
rect 27620 34604 27672 34610
rect 27620 34546 27672 34552
rect 27712 34604 27764 34610
rect 27712 34546 27764 34552
rect 27632 34202 27660 34546
rect 27620 34196 27672 34202
rect 27620 34138 27672 34144
rect 27528 34060 27580 34066
rect 27528 34002 27580 34008
rect 27540 32026 27568 34002
rect 27620 33992 27672 33998
rect 27724 33969 27752 34546
rect 27620 33934 27672 33940
rect 27710 33960 27766 33969
rect 27632 33658 27660 33934
rect 27710 33895 27766 33904
rect 27620 33652 27672 33658
rect 27620 33594 27672 33600
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 27724 31754 27752 33895
rect 27816 33658 27844 35022
rect 27804 33652 27856 33658
rect 27804 33594 27856 33600
rect 27908 33114 27936 35090
rect 28092 34950 28120 35974
rect 28184 35290 28212 36042
rect 28356 35624 28408 35630
rect 28356 35566 28408 35572
rect 28264 35488 28316 35494
rect 28264 35430 28316 35436
rect 28172 35284 28224 35290
rect 28172 35226 28224 35232
rect 28172 35080 28224 35086
rect 28172 35022 28224 35028
rect 28080 34944 28132 34950
rect 28080 34886 28132 34892
rect 27988 34672 28040 34678
rect 27988 34614 28040 34620
rect 28000 34134 28028 34614
rect 28092 34610 28120 34886
rect 28080 34604 28132 34610
rect 28080 34546 28132 34552
rect 28184 34202 28212 35022
rect 28276 34950 28304 35430
rect 28264 34944 28316 34950
rect 28264 34886 28316 34892
rect 28172 34196 28224 34202
rect 28172 34138 28224 34144
rect 27988 34128 28040 34134
rect 27988 34070 28040 34076
rect 28276 33998 28304 34886
rect 28368 34610 28396 35566
rect 28356 34604 28408 34610
rect 28356 34546 28408 34552
rect 28724 34536 28776 34542
rect 28724 34478 28776 34484
rect 28264 33992 28316 33998
rect 28264 33934 28316 33940
rect 27896 33108 27948 33114
rect 27896 33050 27948 33056
rect 27908 32978 27936 33050
rect 27896 32972 27948 32978
rect 27896 32914 27948 32920
rect 27632 31726 27752 31754
rect 27632 31142 27660 31726
rect 27712 31680 27764 31686
rect 27712 31622 27764 31628
rect 27724 31346 27752 31622
rect 27712 31340 27764 31346
rect 27712 31282 27764 31288
rect 27620 31136 27672 31142
rect 27620 31078 27672 31084
rect 27908 30802 27936 32914
rect 28172 32768 28224 32774
rect 28172 32710 28224 32716
rect 27988 32428 28040 32434
rect 27988 32370 28040 32376
rect 28000 31754 28028 32370
rect 28184 32230 28212 32710
rect 28276 32366 28304 33934
rect 28356 32564 28408 32570
rect 28356 32506 28408 32512
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28172 32224 28224 32230
rect 28172 32166 28224 32172
rect 28368 31958 28396 32506
rect 28172 31952 28224 31958
rect 28172 31894 28224 31900
rect 28356 31952 28408 31958
rect 28356 31894 28408 31900
rect 28184 31822 28212 31894
rect 28368 31822 28396 31894
rect 28172 31816 28224 31822
rect 28172 31758 28224 31764
rect 28356 31816 28408 31822
rect 28356 31758 28408 31764
rect 27988 31748 28040 31754
rect 27988 31690 28040 31696
rect 28000 31414 28028 31690
rect 27988 31408 28040 31414
rect 27988 31350 28040 31356
rect 28080 31340 28132 31346
rect 28080 31282 28132 31288
rect 28092 30870 28120 31282
rect 28172 31272 28224 31278
rect 28172 31214 28224 31220
rect 28184 30938 28212 31214
rect 28632 31136 28684 31142
rect 28632 31078 28684 31084
rect 28172 30932 28224 30938
rect 28172 30874 28224 30880
rect 28080 30864 28132 30870
rect 28080 30806 28132 30812
rect 27896 30796 27948 30802
rect 27896 30738 27948 30744
rect 28184 30666 28212 30874
rect 28644 30734 28672 31078
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 27712 30660 27764 30666
rect 27712 30602 27764 30608
rect 28172 30660 28224 30666
rect 28172 30602 28224 30608
rect 27724 29850 27752 30602
rect 28184 30326 28212 30602
rect 28356 30592 28408 30598
rect 28356 30534 28408 30540
rect 28172 30320 28224 30326
rect 28172 30262 28224 30268
rect 27712 29844 27764 29850
rect 27712 29786 27764 29792
rect 28368 29646 28396 30534
rect 28644 30394 28672 30670
rect 28632 30388 28684 30394
rect 28632 30330 28684 30336
rect 28540 30252 28592 30258
rect 28540 30194 28592 30200
rect 28356 29640 28408 29646
rect 28552 29628 28580 30194
rect 28644 30122 28672 30330
rect 28632 30116 28684 30122
rect 28632 30058 28684 30064
rect 28632 29640 28684 29646
rect 28552 29600 28632 29628
rect 28356 29582 28408 29588
rect 28632 29582 28684 29588
rect 28368 28558 28396 29582
rect 28356 28552 28408 28558
rect 28356 28494 28408 28500
rect 28644 28490 28672 29582
rect 28632 28484 28684 28490
rect 28632 28426 28684 28432
rect 27988 28144 28040 28150
rect 27988 28086 28040 28092
rect 27434 27976 27490 27985
rect 27434 27911 27490 27920
rect 26976 27668 27028 27674
rect 26976 27610 27028 27616
rect 26988 25362 27016 27610
rect 27448 26042 27476 27911
rect 27896 27328 27948 27334
rect 27896 27270 27948 27276
rect 27908 26994 27936 27270
rect 28000 27130 28028 28086
rect 28170 27840 28226 27849
rect 28170 27775 28226 27784
rect 28184 27470 28212 27775
rect 28368 27662 28580 27690
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 27988 27124 28040 27130
rect 27988 27066 28040 27072
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 27436 26036 27488 26042
rect 27436 25978 27488 25984
rect 26976 25356 27028 25362
rect 26976 25298 27028 25304
rect 26976 24064 27028 24070
rect 26976 24006 27028 24012
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 26988 23730 27016 24006
rect 27356 23798 27384 24006
rect 27252 23792 27304 23798
rect 27252 23734 27304 23740
rect 27344 23792 27396 23798
rect 27344 23734 27396 23740
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 27264 23066 27292 23734
rect 27342 23216 27398 23225
rect 27342 23151 27344 23160
rect 27396 23151 27398 23160
rect 27344 23122 27396 23128
rect 26976 23044 27028 23050
rect 26976 22986 27028 22992
rect 27264 23038 27568 23066
rect 26988 22506 27016 22986
rect 27264 22642 27292 23038
rect 27540 22982 27568 23038
rect 27436 22976 27488 22982
rect 27436 22918 27488 22924
rect 27528 22976 27580 22982
rect 27528 22918 27580 22924
rect 28264 22976 28316 22982
rect 28264 22918 28316 22924
rect 27448 22710 27476 22918
rect 27436 22704 27488 22710
rect 27436 22646 27488 22652
rect 27712 22704 27764 22710
rect 27712 22646 27764 22652
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 26976 22500 27028 22506
rect 26976 22442 27028 22448
rect 26884 22432 26936 22438
rect 27528 22432 27580 22438
rect 26884 22374 26936 22380
rect 27264 22380 27528 22386
rect 27264 22374 27580 22380
rect 26896 22030 26924 22374
rect 27264 22358 27568 22374
rect 27264 22166 27292 22358
rect 27252 22160 27304 22166
rect 27252 22102 27304 22108
rect 27632 22098 27660 22578
rect 27620 22092 27672 22098
rect 27620 22034 27672 22040
rect 26884 22024 26936 22030
rect 26884 21966 26936 21972
rect 27252 22024 27304 22030
rect 27252 21966 27304 21972
rect 26896 21010 26924 21966
rect 26976 21888 27028 21894
rect 26976 21830 27028 21836
rect 26988 21690 27016 21830
rect 27264 21690 27292 21966
rect 26976 21684 27028 21690
rect 26976 21626 27028 21632
rect 27252 21684 27304 21690
rect 27252 21626 27304 21632
rect 26884 21004 26936 21010
rect 26884 20946 26936 20952
rect 26988 20466 27016 21626
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 27436 21004 27488 21010
rect 27436 20946 27488 20952
rect 27252 20936 27304 20942
rect 27252 20878 27304 20884
rect 26976 20460 27028 20466
rect 26976 20402 27028 20408
rect 26884 19780 26936 19786
rect 26884 19722 26936 19728
rect 26896 19514 26924 19722
rect 26884 19508 26936 19514
rect 26884 19450 26936 19456
rect 26896 18834 26924 19450
rect 26884 18828 26936 18834
rect 26884 18770 26936 18776
rect 26896 17882 26924 18770
rect 26988 18766 27016 20402
rect 27068 20256 27120 20262
rect 27068 20198 27120 20204
rect 27080 19854 27108 20198
rect 27264 19854 27292 20878
rect 27068 19848 27120 19854
rect 27068 19790 27120 19796
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27344 19848 27396 19854
rect 27344 19790 27396 19796
rect 27264 19514 27292 19790
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 27264 18970 27292 19450
rect 27356 19378 27384 19790
rect 27448 19718 27476 20946
rect 27540 20058 27568 21422
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27632 19854 27660 20402
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 27436 19712 27488 19718
rect 27436 19654 27488 19660
rect 27448 19394 27476 19654
rect 27448 19378 27568 19394
rect 27344 19372 27396 19378
rect 27448 19372 27580 19378
rect 27448 19366 27528 19372
rect 27344 19314 27396 19320
rect 27528 19314 27580 19320
rect 27252 18964 27304 18970
rect 27252 18906 27304 18912
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 26988 18306 27016 18702
rect 27356 18698 27384 19314
rect 27344 18692 27396 18698
rect 27344 18634 27396 18640
rect 26988 18278 27108 18306
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26884 17876 26936 17882
rect 26884 17818 26936 17824
rect 26988 17338 27016 18158
rect 27080 17678 27108 18278
rect 27356 18086 27384 18634
rect 27540 18630 27568 19314
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27344 18080 27396 18086
rect 27344 18022 27396 18028
rect 27068 17672 27120 17678
rect 27068 17614 27120 17620
rect 26976 17332 27028 17338
rect 26976 17274 27028 17280
rect 27068 15632 27120 15638
rect 27068 15574 27120 15580
rect 27080 4554 27108 15574
rect 27724 6914 27752 22646
rect 28276 22574 28304 22918
rect 28368 22710 28396 27662
rect 28552 27606 28580 27662
rect 28448 27600 28500 27606
rect 28446 27568 28448 27577
rect 28540 27600 28592 27606
rect 28500 27568 28502 27577
rect 28540 27542 28592 27548
rect 28446 27503 28502 27512
rect 28540 27464 28592 27470
rect 28644 27452 28672 28426
rect 28592 27424 28672 27452
rect 28540 27406 28592 27412
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 28460 27062 28488 27270
rect 28552 27130 28580 27406
rect 28540 27124 28592 27130
rect 28540 27066 28592 27072
rect 28448 27056 28500 27062
rect 28448 26998 28500 27004
rect 28632 23112 28684 23118
rect 28632 23054 28684 23060
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 28644 22642 28672 23054
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28264 22568 28316 22574
rect 28264 22510 28316 22516
rect 28080 21004 28132 21010
rect 28080 20946 28132 20952
rect 27804 20800 27856 20806
rect 27804 20742 27856 20748
rect 27816 20466 27844 20742
rect 28092 20534 28120 20946
rect 28080 20528 28132 20534
rect 28080 20470 28132 20476
rect 27804 20460 27856 20466
rect 27804 20402 27856 20408
rect 28172 19168 28224 19174
rect 28172 19110 28224 19116
rect 28184 18766 28212 19110
rect 28172 18760 28224 18766
rect 28172 18702 28224 18708
rect 28264 18624 28316 18630
rect 28264 18566 28316 18572
rect 28276 18426 28304 18566
rect 28264 18420 28316 18426
rect 28264 18362 28316 18368
rect 27988 18352 28040 18358
rect 27988 18294 28040 18300
rect 28000 17882 28028 18294
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 28460 17202 28488 22578
rect 28736 22094 28764 34478
rect 28828 34406 28856 36518
rect 29184 36304 29236 36310
rect 29184 36246 29236 36252
rect 28908 35488 28960 35494
rect 28908 35430 28960 35436
rect 28920 34678 28948 35430
rect 29092 35012 29144 35018
rect 29092 34954 29144 34960
rect 28908 34672 28960 34678
rect 28908 34614 28960 34620
rect 29000 34536 29052 34542
rect 29000 34478 29052 34484
rect 28816 34400 28868 34406
rect 28816 34342 28868 34348
rect 28828 33998 28856 34342
rect 29012 33998 29040 34478
rect 29104 34134 29132 34954
rect 29092 34128 29144 34134
rect 29092 34070 29144 34076
rect 28816 33992 28868 33998
rect 28816 33934 28868 33940
rect 29000 33992 29052 33998
rect 29000 33934 29052 33940
rect 28828 33522 28856 33934
rect 28816 33516 28868 33522
rect 28816 33458 28868 33464
rect 29012 33318 29040 33934
rect 29000 33312 29052 33318
rect 29000 33254 29052 33260
rect 28816 31816 28868 31822
rect 28816 31758 28868 31764
rect 28828 31210 28856 31758
rect 28908 31340 28960 31346
rect 28908 31282 28960 31288
rect 28816 31204 28868 31210
rect 28816 31146 28868 31152
rect 28816 30932 28868 30938
rect 28816 30874 28868 30880
rect 28828 30258 28856 30874
rect 28920 30598 28948 31282
rect 28908 30592 28960 30598
rect 28908 30534 28960 30540
rect 28816 30252 28868 30258
rect 28816 30194 28868 30200
rect 29000 29640 29052 29646
rect 28920 29588 29000 29594
rect 28920 29582 29052 29588
rect 28920 29566 29040 29582
rect 28920 29102 28948 29566
rect 29000 29504 29052 29510
rect 29000 29446 29052 29452
rect 28908 29096 28960 29102
rect 28908 29038 28960 29044
rect 29012 29034 29040 29446
rect 29196 29170 29224 36246
rect 29644 36032 29696 36038
rect 29644 35974 29696 35980
rect 29656 35766 29684 35974
rect 29644 35760 29696 35766
rect 29644 35702 29696 35708
rect 29368 34468 29420 34474
rect 29368 34410 29420 34416
rect 29276 34060 29328 34066
rect 29276 34002 29328 34008
rect 29288 33590 29316 34002
rect 29380 33590 29408 34410
rect 29276 33584 29328 33590
rect 29276 33526 29328 33532
rect 29368 33584 29420 33590
rect 29368 33526 29420 33532
rect 29644 33312 29696 33318
rect 29644 33254 29696 33260
rect 29656 32910 29684 33254
rect 29644 32904 29696 32910
rect 29644 32846 29696 32852
rect 29736 32360 29788 32366
rect 29736 32302 29788 32308
rect 29644 32224 29696 32230
rect 29644 32166 29696 32172
rect 29276 32020 29328 32026
rect 29276 31962 29328 31968
rect 29288 31414 29316 31962
rect 29656 31822 29684 32166
rect 29748 31958 29776 32302
rect 29736 31952 29788 31958
rect 29736 31894 29788 31900
rect 29840 31906 29868 41386
rect 30012 34944 30064 34950
rect 30012 34886 30064 34892
rect 30024 34678 30052 34886
rect 30012 34672 30064 34678
rect 30012 34614 30064 34620
rect 30012 34536 30064 34542
rect 30012 34478 30064 34484
rect 30024 34066 30052 34478
rect 30012 34060 30064 34066
rect 30012 34002 30064 34008
rect 30024 33658 30052 34002
rect 30012 33652 30064 33658
rect 30012 33594 30064 33600
rect 30024 32910 30052 33594
rect 30012 32904 30064 32910
rect 30012 32846 30064 32852
rect 30012 32768 30064 32774
rect 30012 32710 30064 32716
rect 30024 32434 30052 32710
rect 29920 32428 29972 32434
rect 29920 32370 29972 32376
rect 30012 32428 30064 32434
rect 30012 32370 30064 32376
rect 29932 32026 29960 32370
rect 29920 32020 29972 32026
rect 29920 31962 29972 31968
rect 29840 31878 30052 31906
rect 29644 31816 29696 31822
rect 29644 31758 29696 31764
rect 29828 31816 29880 31822
rect 29828 31758 29880 31764
rect 29276 31408 29328 31414
rect 29276 31350 29328 31356
rect 29184 29164 29236 29170
rect 29184 29106 29236 29112
rect 29000 29028 29052 29034
rect 29000 28970 29052 28976
rect 28906 27976 28962 27985
rect 28906 27911 28908 27920
rect 28960 27911 28962 27920
rect 28908 27882 28960 27888
rect 29012 27878 29040 28970
rect 29092 28552 29144 28558
rect 29092 28494 29144 28500
rect 29196 28506 29224 29106
rect 29460 29096 29512 29102
rect 29460 29038 29512 29044
rect 29000 27872 29052 27878
rect 28906 27840 28962 27849
rect 29000 27814 29052 27820
rect 28906 27775 28962 27784
rect 28816 27600 28868 27606
rect 28814 27568 28816 27577
rect 28868 27568 28870 27577
rect 28920 27554 28948 27775
rect 29104 27674 29132 28494
rect 29196 28478 29316 28506
rect 29184 28416 29236 28422
rect 29184 28358 29236 28364
rect 29196 28082 29224 28358
rect 29184 28076 29236 28082
rect 29184 28018 29236 28024
rect 29092 27668 29144 27674
rect 29092 27610 29144 27616
rect 28920 27538 28994 27554
rect 28920 27532 29006 27538
rect 28920 27526 28954 27532
rect 28814 27503 28870 27512
rect 28954 27474 29006 27480
rect 28908 27328 28960 27334
rect 28828 27288 28908 27316
rect 28828 26994 28856 27288
rect 28908 27270 28960 27276
rect 29104 26994 29132 27610
rect 29288 27606 29316 28478
rect 29276 27600 29328 27606
rect 29276 27542 29328 27548
rect 29368 27328 29420 27334
rect 29368 27270 29420 27276
rect 29380 27062 29408 27270
rect 29368 27056 29420 27062
rect 29368 26998 29420 27004
rect 28816 26988 28868 26994
rect 28816 26930 28868 26936
rect 29092 26988 29144 26994
rect 29092 26930 29144 26936
rect 28816 24200 28868 24206
rect 28816 24142 28868 24148
rect 28828 23662 28856 24142
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 29000 23656 29052 23662
rect 29000 23598 29052 23604
rect 28828 22982 28856 23598
rect 28908 23112 28960 23118
rect 28906 23080 28908 23089
rect 28960 23080 28962 23089
rect 28906 23015 28962 23024
rect 28816 22976 28868 22982
rect 28816 22918 28868 22924
rect 29012 22506 29040 23598
rect 29000 22500 29052 22506
rect 29000 22442 29052 22448
rect 29012 22098 29040 22442
rect 28736 22066 28948 22094
rect 28540 21956 28592 21962
rect 28540 21898 28592 21904
rect 28552 21690 28580 21898
rect 28540 21684 28592 21690
rect 28540 21626 28592 21632
rect 28632 20528 28684 20534
rect 28632 20470 28684 20476
rect 28644 20058 28672 20470
rect 28632 20052 28684 20058
rect 28632 19994 28684 20000
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 27632 6886 27752 6914
rect 27068 4548 27120 4554
rect 27068 4490 27120 4496
rect 27252 4548 27304 4554
rect 27252 4490 27304 4496
rect 27264 3466 27292 4490
rect 27252 3460 27304 3466
rect 27252 3402 27304 3408
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 26792 2644 26844 2650
rect 26792 2586 26844 2592
rect 25504 2576 25556 2582
rect 25504 2518 25556 2524
rect 25596 2576 25648 2582
rect 25596 2518 25648 2524
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25148 800 25176 2450
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26436 800 26464 2382
rect 27080 800 27108 2994
rect 27264 2854 27292 3402
rect 27632 3126 27660 6886
rect 28460 4146 28488 17138
rect 28448 4140 28500 4146
rect 28448 4082 28500 4088
rect 28920 3670 28948 22066
rect 29000 22092 29052 22098
rect 29000 22034 29052 22040
rect 29092 18080 29144 18086
rect 29092 18022 29144 18028
rect 29104 17202 29132 18022
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 27620 3120 27672 3126
rect 27620 3062 27672 3068
rect 27252 2848 27304 2854
rect 27252 2790 27304 2796
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 28368 800 28396 2314
rect 29472 2310 29500 29038
rect 29552 27872 29604 27878
rect 29552 27814 29604 27820
rect 29564 27538 29592 27814
rect 29552 27532 29604 27538
rect 29552 27474 29604 27480
rect 29736 24132 29788 24138
rect 29736 24074 29788 24080
rect 29748 23322 29776 24074
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 29552 22976 29604 22982
rect 29552 22918 29604 22924
rect 29564 22642 29592 22918
rect 29552 22636 29604 22642
rect 29552 22578 29604 22584
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 29564 20602 29592 20878
rect 29552 20596 29604 20602
rect 29552 20538 29604 20544
rect 29644 17604 29696 17610
rect 29644 17546 29696 17552
rect 29656 16794 29684 17546
rect 29644 16788 29696 16794
rect 29644 16730 29696 16736
rect 29550 3632 29606 3641
rect 29550 3567 29552 3576
rect 29604 3567 29606 3576
rect 29552 3538 29604 3544
rect 29736 3460 29788 3466
rect 29736 3402 29788 3408
rect 29748 2650 29776 3402
rect 29736 2644 29788 2650
rect 29736 2586 29788 2592
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 29460 2304 29512 2310
rect 29460 2246 29512 2252
rect 29656 800 29684 2382
rect 29840 2378 29868 31758
rect 29920 23656 29972 23662
rect 29920 23598 29972 23604
rect 29932 22710 29960 23598
rect 29920 22704 29972 22710
rect 29920 22646 29972 22652
rect 30024 17610 30052 31878
rect 30116 31278 30144 46990
rect 31668 46368 31720 46374
rect 31668 46310 31720 46316
rect 31680 46034 31708 46310
rect 32232 46034 32260 49200
rect 38028 47410 38056 49200
rect 37292 47382 38056 47410
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 34520 46368 34572 46374
rect 34520 46310 34572 46316
rect 31668 46028 31720 46034
rect 31668 45970 31720 45976
rect 32220 46028 32272 46034
rect 32220 45970 32272 45976
rect 32220 45892 32272 45898
rect 32220 45834 32272 45840
rect 32232 45626 32260 45834
rect 32220 45620 32272 45626
rect 32220 45562 32272 45568
rect 32128 45484 32180 45490
rect 32128 45426 32180 45432
rect 31300 35692 31352 35698
rect 31300 35634 31352 35640
rect 31208 35488 31260 35494
rect 31208 35430 31260 35436
rect 31220 35018 31248 35430
rect 30472 35012 30524 35018
rect 30472 34954 30524 34960
rect 31208 35012 31260 35018
rect 31208 34954 31260 34960
rect 30196 34944 30248 34950
rect 30196 34886 30248 34892
rect 30208 34610 30236 34886
rect 30484 34746 30512 34954
rect 30472 34740 30524 34746
rect 30472 34682 30524 34688
rect 30196 34604 30248 34610
rect 30196 34546 30248 34552
rect 31116 34604 31168 34610
rect 31116 34546 31168 34552
rect 30208 34066 30236 34546
rect 31128 34202 31156 34546
rect 31116 34196 31168 34202
rect 31116 34138 31168 34144
rect 30196 34060 30248 34066
rect 30196 34002 30248 34008
rect 30288 33516 30340 33522
rect 30288 33458 30340 33464
rect 30300 32774 30328 33458
rect 30564 32836 30616 32842
rect 30564 32778 30616 32784
rect 30288 32768 30340 32774
rect 30288 32710 30340 32716
rect 30300 32502 30328 32710
rect 30576 32570 30604 32778
rect 30564 32564 30616 32570
rect 30564 32506 30616 32512
rect 30288 32496 30340 32502
rect 30288 32438 30340 32444
rect 31312 32434 31340 35634
rect 31392 32836 31444 32842
rect 31392 32778 31444 32784
rect 31404 32570 31432 32778
rect 31392 32564 31444 32570
rect 31392 32506 31444 32512
rect 30196 32428 30248 32434
rect 30196 32370 30248 32376
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 30208 32042 30236 32370
rect 30208 32014 30328 32042
rect 30196 31952 30248 31958
rect 30196 31894 30248 31900
rect 30208 31482 30236 31894
rect 30196 31476 30248 31482
rect 30196 31418 30248 31424
rect 30104 31272 30156 31278
rect 30104 31214 30156 31220
rect 30104 31136 30156 31142
rect 30104 31078 30156 31084
rect 30116 30598 30144 31078
rect 30104 30592 30156 30598
rect 30104 30534 30156 30540
rect 30116 30258 30144 30534
rect 30300 30258 30328 32014
rect 31024 31136 31076 31142
rect 31024 31078 31076 31084
rect 30472 30660 30524 30666
rect 30472 30602 30524 30608
rect 30484 30394 30512 30602
rect 30472 30388 30524 30394
rect 30472 30330 30524 30336
rect 30380 30320 30432 30326
rect 30380 30262 30432 30268
rect 30104 30252 30156 30258
rect 30104 30194 30156 30200
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30300 29646 30328 30194
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 30392 29170 30420 30262
rect 31036 30258 31064 31078
rect 31116 30660 31168 30666
rect 31116 30602 31168 30608
rect 31024 30252 31076 30258
rect 31024 30194 31076 30200
rect 31128 29850 31156 30602
rect 31116 29844 31168 29850
rect 31116 29786 31168 29792
rect 30840 29640 30892 29646
rect 30840 29582 30892 29588
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30196 28960 30248 28966
rect 30196 28902 30248 28908
rect 30208 28626 30236 28902
rect 30196 28620 30248 28626
rect 30196 28562 30248 28568
rect 30852 28082 30880 29582
rect 31668 29164 31720 29170
rect 31668 29106 31720 29112
rect 31680 28694 31708 29106
rect 31668 28688 31720 28694
rect 31668 28630 31720 28636
rect 30932 28484 30984 28490
rect 30932 28426 30984 28432
rect 30944 28218 30972 28426
rect 30932 28212 30984 28218
rect 30932 28154 30984 28160
rect 30840 28076 30892 28082
rect 30840 28018 30892 28024
rect 30852 27470 30880 28018
rect 30840 27464 30892 27470
rect 30840 27406 30892 27412
rect 30380 27328 30432 27334
rect 30380 27270 30432 27276
rect 30392 27062 30420 27270
rect 30380 27056 30432 27062
rect 30380 26998 30432 27004
rect 32140 26926 32168 45426
rect 34532 43858 34560 46310
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34520 43852 34572 43858
rect 34520 43794 34572 43800
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 32220 27668 32272 27674
rect 32220 27610 32272 27616
rect 32128 26920 32180 26926
rect 32128 26862 32180 26868
rect 32232 21010 32260 27610
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 37292 23798 37320 47382
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 38120 46578 38148 46990
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 37740 46504 37792 46510
rect 37740 46446 37792 46452
rect 38384 46504 38436 46510
rect 38384 46446 38436 46452
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 37280 23792 37332 23798
rect 37280 23734 37332 23740
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 32220 21004 32272 21010
rect 32220 20946 32272 20952
rect 30564 20868 30616 20874
rect 30564 20810 30616 20816
rect 30576 20602 30604 20810
rect 30564 20596 30616 20602
rect 30564 20538 30616 20544
rect 30104 20528 30156 20534
rect 30104 20470 30156 20476
rect 30012 17604 30064 17610
rect 30012 17546 30064 17552
rect 30116 16114 30144 20470
rect 30472 20460 30524 20466
rect 30472 20402 30524 20408
rect 30484 19990 30512 20402
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 30472 19984 30524 19990
rect 30472 19926 30524 19932
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 30656 17604 30708 17610
rect 30656 17546 30708 17552
rect 30668 17066 30696 17546
rect 30932 17128 30984 17134
rect 30932 17070 30984 17076
rect 30656 17060 30708 17066
rect 30656 17002 30708 17008
rect 30196 16516 30248 16522
rect 30196 16458 30248 16464
rect 30208 16250 30236 16458
rect 30196 16244 30248 16250
rect 30196 16186 30248 16192
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 30472 13252 30524 13258
rect 30472 13194 30524 13200
rect 29828 2372 29880 2378
rect 29828 2314 29880 2320
rect 18892 734 19104 762
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30484 762 30512 13194
rect 30944 8022 30972 17070
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 30932 8016 30984 8022
rect 30932 7958 30984 7964
rect 33876 8016 33928 8022
rect 33876 7958 33928 7964
rect 33784 4072 33836 4078
rect 33784 4014 33836 4020
rect 33796 3534 33824 4014
rect 33784 3528 33836 3534
rect 33784 3470 33836 3476
rect 32956 3460 33008 3466
rect 32956 3402 33008 3408
rect 32220 3392 32272 3398
rect 32220 3334 32272 3340
rect 30760 870 30972 898
rect 30760 762 30788 870
rect 30944 800 30972 870
rect 32232 800 32260 3334
rect 32968 3058 32996 3402
rect 33888 3398 33916 7958
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35900 4140 35952 4146
rect 35900 4082 35952 4088
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35912 3534 35940 4082
rect 37752 3534 37780 46446
rect 38396 46170 38424 46446
rect 39960 46374 39988 49200
rect 40788 47410 40816 49286
rect 41206 49200 41318 49286
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 43782 49200 43894 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49200 46470 50000
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 40052 47382 40816 47410
rect 39948 46368 40000 46374
rect 39948 46310 40000 46316
rect 38384 46164 38436 46170
rect 38384 46106 38436 46112
rect 38292 46096 38344 46102
rect 38292 46038 38344 46044
rect 38304 45966 38332 46038
rect 38292 45960 38344 45966
rect 38292 45902 38344 45908
rect 38304 23254 38332 45902
rect 40052 24138 40080 47382
rect 40408 46980 40460 46986
rect 40408 46922 40460 46928
rect 40420 28626 40448 46922
rect 41328 46368 41380 46374
rect 41328 46310 41380 46316
rect 41340 46034 41368 46310
rect 41892 46034 41920 49200
rect 42536 46442 42564 49200
rect 42616 47048 42668 47054
rect 42616 46990 42668 46996
rect 42628 46594 42656 46990
rect 42628 46566 42748 46594
rect 42616 46504 42668 46510
rect 42616 46446 42668 46452
rect 42524 46436 42576 46442
rect 42524 46378 42576 46384
rect 41328 46028 41380 46034
rect 41328 45970 41380 45976
rect 41880 46028 41932 46034
rect 41880 45970 41932 45976
rect 41512 45892 41564 45898
rect 41512 45834 41564 45840
rect 41524 45558 41552 45834
rect 41696 45824 41748 45830
rect 41696 45766 41748 45772
rect 41512 45552 41564 45558
rect 41512 45494 41564 45500
rect 41708 45490 41736 45766
rect 42628 45626 42656 46446
rect 42616 45620 42668 45626
rect 42616 45562 42668 45568
rect 41052 45484 41104 45490
rect 41052 45426 41104 45432
rect 41696 45484 41748 45490
rect 41696 45426 41748 45432
rect 41064 45354 41092 45426
rect 42432 45416 42484 45422
rect 42432 45358 42484 45364
rect 42616 45416 42668 45422
rect 42616 45358 42668 45364
rect 41052 45348 41104 45354
rect 41052 45290 41104 45296
rect 42444 44946 42472 45358
rect 42432 44940 42484 44946
rect 42432 44882 42484 44888
rect 42628 44402 42656 45358
rect 42616 44396 42668 44402
rect 42616 44338 42668 44344
rect 42720 44334 42748 46566
rect 43180 45422 43208 49200
rect 43260 46980 43312 46986
rect 43260 46922 43312 46928
rect 42800 45416 42852 45422
rect 42800 45358 42852 45364
rect 43168 45416 43220 45422
rect 43168 45358 43220 45364
rect 42812 45082 42840 45358
rect 43272 45082 43300 46922
rect 43824 45966 43852 49200
rect 44180 46096 44232 46102
rect 44180 46038 44232 46044
rect 43812 45960 43864 45966
rect 43812 45902 43864 45908
rect 43996 45824 44048 45830
rect 43996 45766 44048 45772
rect 42800 45076 42852 45082
rect 42800 45018 42852 45024
rect 43260 45076 43312 45082
rect 43260 45018 43312 45024
rect 43168 44872 43220 44878
rect 43168 44814 43220 44820
rect 42708 44328 42760 44334
rect 42708 44270 42760 44276
rect 41420 33312 41472 33318
rect 41420 33254 41472 33260
rect 41432 32298 41460 33254
rect 41420 32292 41472 32298
rect 41420 32234 41472 32240
rect 40408 28620 40460 28626
rect 40408 28562 40460 28568
rect 40776 24336 40828 24342
rect 40776 24278 40828 24284
rect 40040 24132 40092 24138
rect 40040 24074 40092 24080
rect 40788 23866 40816 24278
rect 40776 23860 40828 23866
rect 40776 23802 40828 23808
rect 40788 23730 40816 23802
rect 41340 23730 41460 23746
rect 40776 23724 40828 23730
rect 40776 23666 40828 23672
rect 41340 23724 41472 23730
rect 41340 23718 41420 23724
rect 41340 23526 41368 23718
rect 41420 23666 41472 23672
rect 41328 23520 41380 23526
rect 41328 23462 41380 23468
rect 38292 23248 38344 23254
rect 38292 23190 38344 23196
rect 41340 23118 41368 23462
rect 41328 23112 41380 23118
rect 41328 23054 41380 23060
rect 43180 22234 43208 44814
rect 44008 35154 44036 45766
rect 44192 44402 44220 46038
rect 44468 44878 44496 49200
rect 45112 47122 45140 49200
rect 45100 47116 45152 47122
rect 45100 47058 45152 47064
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45204 46594 45232 46990
rect 45468 46980 45520 46986
rect 45468 46922 45520 46928
rect 45204 46566 45324 46594
rect 45192 46504 45244 46510
rect 45192 46446 45244 46452
rect 44916 46368 44968 46374
rect 44916 46310 44968 46316
rect 44456 44872 44508 44878
rect 44456 44814 44508 44820
rect 44180 44396 44232 44402
rect 44180 44338 44232 44344
rect 44732 39976 44784 39982
rect 44732 39918 44784 39924
rect 43996 35148 44048 35154
rect 43996 35090 44048 35096
rect 44180 34060 44232 34066
rect 44180 34002 44232 34008
rect 44192 31822 44220 34002
rect 44180 31816 44232 31822
rect 44180 31758 44232 31764
rect 43168 22228 43220 22234
rect 43168 22170 43220 22176
rect 40224 17536 40276 17542
rect 40224 17478 40276 17484
rect 39764 16992 39816 16998
rect 39764 16934 39816 16940
rect 39776 16658 39804 16934
rect 40236 16658 40264 17478
rect 39764 16652 39816 16658
rect 39764 16594 39816 16600
rect 40224 16652 40276 16658
rect 40224 16594 40276 16600
rect 40408 16516 40460 16522
rect 40408 16458 40460 16464
rect 39672 4548 39724 4554
rect 39672 4490 39724 4496
rect 38476 4140 38528 4146
rect 38476 4082 38528 4088
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 37740 3528 37792 3534
rect 37740 3470 37792 3476
rect 36176 3460 36228 3466
rect 36176 3402 36228 3408
rect 33140 3392 33192 3398
rect 33140 3334 33192 3340
rect 33876 3392 33928 3398
rect 33876 3334 33928 3340
rect 33152 3126 33180 3334
rect 36188 3194 36216 3402
rect 35808 3188 35860 3194
rect 35808 3130 35860 3136
rect 36176 3188 36228 3194
rect 36176 3130 36228 3136
rect 33140 3120 33192 3126
rect 33140 3062 33192 3068
rect 32956 3052 33008 3058
rect 32956 2994 33008 3000
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 33520 800 33548 2926
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35820 2514 35848 3130
rect 38488 3058 38516 4082
rect 39580 3936 39632 3942
rect 39580 3878 39632 3884
rect 39120 3732 39172 3738
rect 39120 3674 39172 3680
rect 39132 3097 39160 3674
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 39118 3088 39174 3097
rect 36084 3052 36136 3058
rect 36084 2994 36136 3000
rect 38476 3052 38528 3058
rect 39118 3023 39174 3032
rect 38476 2994 38528 3000
rect 35808 2508 35860 2514
rect 35808 2450 35860 2456
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35452 800 35480 2382
rect 36096 800 36124 2994
rect 39224 2650 39252 3470
rect 39212 2644 39264 2650
rect 39212 2586 39264 2592
rect 39592 2446 39620 3878
rect 39684 3466 39712 4490
rect 39856 4140 39908 4146
rect 39856 4082 39908 4088
rect 39672 3460 39724 3466
rect 39672 3402 39724 3408
rect 39764 3460 39816 3466
rect 39764 3402 39816 3408
rect 39776 2990 39804 3402
rect 39868 3194 39896 4082
rect 39960 3726 40172 3754
rect 39960 3602 39988 3726
rect 39948 3596 40000 3602
rect 39948 3538 40000 3544
rect 40040 3596 40092 3602
rect 40040 3538 40092 3544
rect 40052 3482 40080 3538
rect 39960 3454 40080 3482
rect 39856 3188 39908 3194
rect 39856 3130 39908 3136
rect 39764 2984 39816 2990
rect 39764 2926 39816 2932
rect 39856 2984 39908 2990
rect 39856 2926 39908 2932
rect 39672 2848 39724 2854
rect 39868 2802 39896 2926
rect 39724 2796 39896 2802
rect 39672 2790 39896 2796
rect 39684 2774 39896 2790
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 39580 2440 39632 2446
rect 39580 2382 39632 2388
rect 38028 800 38056 2382
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 39316 800 39344 2314
rect 39960 800 39988 3454
rect 40144 3194 40172 3726
rect 40132 3188 40184 3194
rect 40132 3130 40184 3136
rect 40130 3088 40186 3097
rect 40130 3023 40186 3032
rect 40144 2854 40172 3023
rect 40132 2848 40184 2854
rect 40132 2790 40184 2796
rect 40420 2650 40448 16458
rect 44744 12434 44772 39918
rect 44928 35894 44956 46310
rect 45100 45280 45152 45286
rect 45100 45222 45152 45228
rect 45112 45014 45140 45222
rect 45204 45082 45232 46446
rect 45192 45076 45244 45082
rect 45192 45018 45244 45024
rect 45100 45008 45152 45014
rect 45100 44950 45152 44956
rect 45296 43314 45324 46566
rect 45376 46504 45428 46510
rect 45376 46446 45428 46452
rect 45388 44538 45416 46446
rect 45480 44538 45508 46922
rect 45756 45966 45784 49200
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 46296 45960 46348 45966
rect 46296 45902 46348 45908
rect 45744 45824 45796 45830
rect 45744 45766 45796 45772
rect 45376 44532 45428 44538
rect 45376 44474 45428 44480
rect 45468 44532 45520 44538
rect 45468 44474 45520 44480
rect 45284 43308 45336 43314
rect 45284 43250 45336 43256
rect 45756 38962 45784 45766
rect 45836 45484 45888 45490
rect 45836 45426 45888 45432
rect 45848 45082 45876 45426
rect 45928 45280 45980 45286
rect 45928 45222 45980 45228
rect 45836 45076 45888 45082
rect 45836 45018 45888 45024
rect 45744 38956 45796 38962
rect 45744 38898 45796 38904
rect 45652 38820 45704 38826
rect 45652 38762 45704 38768
rect 45664 35894 45692 38762
rect 45836 38344 45888 38350
rect 45836 38286 45888 38292
rect 44928 35866 45140 35894
rect 45664 35866 45784 35894
rect 45008 26444 45060 26450
rect 45008 26386 45060 26392
rect 44744 12406 44956 12434
rect 44732 5092 44784 5098
rect 44732 5034 44784 5040
rect 44744 4690 44772 5034
rect 44732 4684 44784 4690
rect 44732 4626 44784 4632
rect 43812 4616 43864 4622
rect 43812 4558 43864 4564
rect 43720 4480 43772 4486
rect 43720 4422 43772 4428
rect 40592 4276 40644 4282
rect 40592 4218 40644 4224
rect 40500 4140 40552 4146
rect 40500 4082 40552 4088
rect 40512 3738 40540 4082
rect 40500 3732 40552 3738
rect 40500 3674 40552 3680
rect 40604 3126 40632 4218
rect 43732 4214 43760 4422
rect 41052 4208 41104 4214
rect 41052 4150 41104 4156
rect 43720 4208 43772 4214
rect 43720 4150 43772 4156
rect 41064 4010 41092 4150
rect 41696 4072 41748 4078
rect 41696 4014 41748 4020
rect 41052 4004 41104 4010
rect 41052 3946 41104 3952
rect 41512 3936 41564 3942
rect 41512 3878 41564 3884
rect 41524 3602 41552 3878
rect 40684 3596 40736 3602
rect 40684 3538 40736 3544
rect 41512 3596 41564 3602
rect 41512 3538 41564 3544
rect 40592 3120 40644 3126
rect 40592 3062 40644 3068
rect 40696 2990 40724 3538
rect 41708 3466 41736 4014
rect 42892 3936 42944 3942
rect 42892 3878 42944 3884
rect 41696 3460 41748 3466
rect 41696 3402 41748 3408
rect 42708 3460 42760 3466
rect 42708 3402 42760 3408
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40408 2644 40460 2650
rect 40408 2586 40460 2592
rect 41708 2514 41736 3402
rect 42524 3392 42576 3398
rect 42524 3334 42576 3340
rect 41696 2508 41748 2514
rect 41696 2450 41748 2456
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40604 800 40632 2314
rect 41248 800 41276 2382
rect 42536 800 42564 3334
rect 42720 3058 42748 3402
rect 42904 3126 42932 3878
rect 42892 3120 42944 3126
rect 42892 3062 42944 3068
rect 43168 3120 43220 3126
rect 43168 3062 43220 3068
rect 42708 3052 42760 3058
rect 42708 2994 42760 3000
rect 43180 800 43208 3062
rect 43824 800 43852 4558
rect 44928 4146 44956 12406
rect 44916 4140 44968 4146
rect 44916 4082 44968 4088
rect 44928 3505 44956 4082
rect 45020 4078 45048 26386
rect 45112 17270 45140 35866
rect 45560 34128 45612 34134
rect 45560 34070 45612 34076
rect 45572 31754 45600 34070
rect 45572 31726 45692 31754
rect 45558 28656 45614 28665
rect 45558 28591 45614 28600
rect 45572 27674 45600 28591
rect 45560 27668 45612 27674
rect 45560 27610 45612 27616
rect 45560 24880 45612 24886
rect 45560 24822 45612 24828
rect 45376 24744 45428 24750
rect 45376 24686 45428 24692
rect 45388 23866 45416 24686
rect 45572 23905 45600 24822
rect 45558 23896 45614 23905
rect 45376 23860 45428 23866
rect 45558 23831 45614 23840
rect 45376 23802 45428 23808
rect 45192 20256 45244 20262
rect 45192 20198 45244 20204
rect 45204 19990 45232 20198
rect 45192 19984 45244 19990
rect 45192 19926 45244 19932
rect 45204 19446 45232 19926
rect 45560 19916 45612 19922
rect 45560 19858 45612 19864
rect 45192 19440 45244 19446
rect 45192 19382 45244 19388
rect 45572 19378 45600 19858
rect 45560 19372 45612 19378
rect 45560 19314 45612 19320
rect 45100 17264 45152 17270
rect 45100 17206 45152 17212
rect 45192 17128 45244 17134
rect 45192 17070 45244 17076
rect 45204 15434 45232 17070
rect 45468 16992 45520 16998
rect 45468 16934 45520 16940
rect 45480 15745 45508 16934
rect 45664 16590 45692 31726
rect 45756 25294 45784 35866
rect 45848 27130 45876 38286
rect 45836 27124 45888 27130
rect 45836 27066 45888 27072
rect 45836 26988 45888 26994
rect 45836 26930 45888 26936
rect 45848 26382 45876 26930
rect 45836 26376 45888 26382
rect 45836 26318 45888 26324
rect 45848 25906 45876 26318
rect 45836 25900 45888 25906
rect 45836 25842 45888 25848
rect 45848 25430 45876 25842
rect 45836 25424 45888 25430
rect 45836 25366 45888 25372
rect 45744 25288 45796 25294
rect 45744 25230 45796 25236
rect 45756 23594 45784 25230
rect 45744 23588 45796 23594
rect 45744 23530 45796 23536
rect 45836 22636 45888 22642
rect 45836 22578 45888 22584
rect 45744 20256 45796 20262
rect 45744 20198 45796 20204
rect 45756 19922 45784 20198
rect 45744 19916 45796 19922
rect 45744 19858 45796 19864
rect 45848 19666 45876 22578
rect 45940 20466 45968 45222
rect 46020 44804 46072 44810
rect 46020 44746 46072 44752
rect 46032 31890 46060 44746
rect 46308 44402 46336 45902
rect 46400 45558 46428 49200
rect 46846 47696 46902 47705
rect 46846 47631 46902 47640
rect 46860 46510 46888 47631
rect 46848 46504 46900 46510
rect 46848 46446 46900 46452
rect 47044 46034 47072 49200
rect 47688 47054 47716 49200
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47860 46572 47912 46578
rect 47860 46514 47912 46520
rect 47872 46345 47900 46514
rect 47858 46336 47914 46345
rect 47858 46271 47914 46280
rect 47032 46028 47084 46034
rect 47032 45970 47084 45976
rect 46480 45892 46532 45898
rect 46480 45834 46532 45840
rect 46492 45626 46520 45834
rect 48134 45656 48190 45665
rect 46480 45620 46532 45626
rect 48134 45591 48190 45600
rect 46480 45562 46532 45568
rect 46388 45552 46440 45558
rect 46388 45494 46440 45500
rect 46480 45484 46532 45490
rect 47308 45484 47360 45490
rect 46532 45444 46612 45472
rect 46480 45426 46532 45432
rect 46296 44396 46348 44402
rect 46296 44338 46348 44344
rect 46584 41138 46612 45444
rect 47308 45426 47360 45432
rect 46940 45416 46992 45422
rect 46940 45358 46992 45364
rect 46756 45348 46808 45354
rect 46756 45290 46808 45296
rect 46572 41132 46624 41138
rect 46572 41074 46624 41080
rect 46112 40520 46164 40526
rect 46112 40462 46164 40468
rect 46124 40050 46152 40462
rect 46204 40452 46256 40458
rect 46204 40394 46256 40400
rect 46112 40044 46164 40050
rect 46112 39986 46164 39992
rect 46216 35894 46244 40394
rect 46480 39840 46532 39846
rect 46480 39782 46532 39788
rect 46492 39506 46520 39782
rect 46480 39500 46532 39506
rect 46480 39442 46532 39448
rect 46124 35866 46244 35894
rect 46020 31884 46072 31890
rect 46020 31826 46072 31832
rect 46020 26376 46072 26382
rect 46020 26318 46072 26324
rect 45928 20460 45980 20466
rect 45928 20402 45980 20408
rect 45848 19638 45968 19666
rect 45744 19372 45796 19378
rect 45744 19314 45796 19320
rect 45756 18766 45784 19314
rect 45744 18760 45796 18766
rect 45744 18702 45796 18708
rect 45652 16584 45704 16590
rect 45652 16526 45704 16532
rect 45466 15736 45522 15745
rect 45466 15671 45522 15680
rect 45192 15428 45244 15434
rect 45192 15370 45244 15376
rect 45204 15026 45232 15370
rect 45192 15020 45244 15026
rect 45192 14962 45244 14968
rect 45652 14952 45704 14958
rect 45652 14894 45704 14900
rect 45664 14618 45692 14894
rect 45652 14612 45704 14618
rect 45652 14554 45704 14560
rect 45376 13388 45428 13394
rect 45376 13330 45428 13336
rect 45192 13252 45244 13258
rect 45192 13194 45244 13200
rect 45204 12850 45232 13194
rect 45388 12850 45416 13330
rect 45192 12844 45244 12850
rect 45192 12786 45244 12792
rect 45376 12844 45428 12850
rect 45376 12786 45428 12792
rect 45100 9988 45152 9994
rect 45100 9930 45152 9936
rect 45008 4072 45060 4078
rect 45008 4014 45060 4020
rect 44914 3496 44970 3505
rect 44914 3431 44970 3440
rect 45008 2848 45060 2854
rect 45008 2790 45060 2796
rect 45020 1850 45048 2790
rect 45112 2514 45140 9930
rect 45204 4554 45232 12786
rect 45756 12442 45784 18702
rect 45940 16794 45968 19638
rect 46032 17746 46060 26318
rect 46124 19242 46152 35866
rect 46296 32904 46348 32910
rect 46296 32846 46348 32852
rect 46308 32434 46336 32846
rect 46296 32428 46348 32434
rect 46296 32370 46348 32376
rect 46584 31754 46612 41074
rect 46768 40050 46796 45290
rect 46952 43194 46980 45358
rect 47032 44804 47084 44810
rect 47032 44746 47084 44752
rect 47044 43314 47072 44746
rect 47320 44402 47348 45426
rect 47676 45280 47728 45286
rect 47676 45222 47728 45228
rect 47400 45076 47452 45082
rect 47400 45018 47452 45024
rect 47308 44396 47360 44402
rect 47308 44338 47360 44344
rect 47032 43308 47084 43314
rect 47032 43250 47084 43256
rect 46952 43166 47072 43194
rect 46940 41540 46992 41546
rect 46940 41482 46992 41488
rect 46952 41274 46980 41482
rect 46940 41268 46992 41274
rect 46940 41210 46992 41216
rect 46756 40044 46808 40050
rect 46756 39986 46808 39992
rect 46768 31754 46796 39986
rect 47044 38962 47072 43166
rect 47124 42220 47176 42226
rect 47124 42162 47176 42168
rect 47032 38956 47084 38962
rect 47032 38898 47084 38904
rect 46940 38752 46992 38758
rect 46940 38694 46992 38700
rect 46952 38418 46980 38694
rect 46940 38412 46992 38418
rect 46940 38354 46992 38360
rect 47032 37664 47084 37670
rect 47032 37606 47084 37612
rect 47044 37126 47072 37606
rect 47032 37120 47084 37126
rect 47032 37062 47084 37068
rect 47136 35894 47164 42162
rect 47320 41414 47348 44338
rect 47412 41970 47440 45018
rect 47688 44946 47716 45222
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 47676 44940 47728 44946
rect 47676 44882 47728 44888
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 47584 44736 47636 44742
rect 47584 44678 47636 44684
rect 47596 42226 47624 44678
rect 47676 44192 47728 44198
rect 47676 44134 47728 44140
rect 47688 43858 47716 44134
rect 48240 43858 48268 44911
rect 47676 43852 47728 43858
rect 47676 43794 47728 43800
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 47768 43104 47820 43110
rect 47768 43046 47820 43052
rect 47780 42770 47808 43046
rect 47768 42764 47820 42770
rect 47768 42706 47820 42712
rect 47676 42628 47728 42634
rect 47676 42570 47728 42576
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 47688 42362 47716 42570
rect 47676 42356 47728 42362
rect 47676 42298 47728 42304
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 47584 42220 47636 42226
rect 48134 42191 48190 42200
rect 47584 42162 47636 42168
rect 47412 41942 47624 41970
rect 47320 41386 47532 41414
rect 47308 38956 47360 38962
rect 47308 38898 47360 38904
rect 47044 35866 47164 35894
rect 47044 33946 47072 35866
rect 47124 34944 47176 34950
rect 47124 34886 47176 34892
rect 47136 34066 47164 34886
rect 47216 34400 47268 34406
rect 47216 34342 47268 34348
rect 47124 34060 47176 34066
rect 47124 34002 47176 34008
rect 47044 33918 47164 33946
rect 47228 33930 47256 34342
rect 46400 31726 46612 31754
rect 46676 31726 46796 31754
rect 46296 28552 46348 28558
rect 46296 28494 46348 28500
rect 46204 27124 46256 27130
rect 46204 27066 46256 27072
rect 46216 25106 46244 27066
rect 46308 25294 46336 28494
rect 46400 26450 46428 31726
rect 46676 26874 46704 31726
rect 46846 31376 46902 31385
rect 46846 31311 46902 31320
rect 46754 30016 46810 30025
rect 46754 29951 46810 29960
rect 46492 26846 46704 26874
rect 46388 26444 46440 26450
rect 46388 26386 46440 26392
rect 46388 26308 46440 26314
rect 46388 26250 46440 26256
rect 46400 26042 46428 26250
rect 46388 26036 46440 26042
rect 46388 25978 46440 25984
rect 46296 25288 46348 25294
rect 46348 25236 46428 25242
rect 46296 25230 46428 25236
rect 46308 25214 46428 25230
rect 46216 25078 46336 25106
rect 46204 24948 46256 24954
rect 46204 24890 46256 24896
rect 46216 20058 46244 24890
rect 46308 20806 46336 25078
rect 46400 21026 46428 25214
rect 46492 21418 46520 26846
rect 46768 26194 46796 29951
rect 46584 26166 46796 26194
rect 46584 23798 46612 26166
rect 46664 26036 46716 26042
rect 46664 25978 46716 25984
rect 46572 23792 46624 23798
rect 46572 23734 46624 23740
rect 46572 22568 46624 22574
rect 46570 22536 46572 22545
rect 46624 22536 46626 22545
rect 46570 22471 46626 22480
rect 46480 21412 46532 21418
rect 46480 21354 46532 21360
rect 46400 20998 46612 21026
rect 46480 20868 46532 20874
rect 46480 20810 46532 20816
rect 46296 20800 46348 20806
rect 46296 20742 46348 20748
rect 46492 20602 46520 20810
rect 46388 20596 46440 20602
rect 46388 20538 46440 20544
rect 46480 20596 46532 20602
rect 46480 20538 46532 20544
rect 46296 20528 46348 20534
rect 46296 20470 46348 20476
rect 46204 20052 46256 20058
rect 46204 19994 46256 20000
rect 46308 19938 46336 20470
rect 46216 19910 46336 19938
rect 46112 19236 46164 19242
rect 46112 19178 46164 19184
rect 46216 19122 46244 19910
rect 46296 19712 46348 19718
rect 46296 19654 46348 19660
rect 46124 19094 46244 19122
rect 46020 17740 46072 17746
rect 46020 17682 46072 17688
rect 45928 16788 45980 16794
rect 45928 16730 45980 16736
rect 46124 16674 46152 19094
rect 46308 18766 46336 19654
rect 46400 19378 46428 20538
rect 46480 20460 46532 20466
rect 46480 20402 46532 20408
rect 46388 19372 46440 19378
rect 46388 19314 46440 19320
rect 46388 19236 46440 19242
rect 46388 19178 46440 19184
rect 46296 18760 46348 18766
rect 46296 18702 46348 18708
rect 46400 18578 46428 19178
rect 46308 18550 46428 18578
rect 46204 18080 46256 18086
rect 46204 18022 46256 18028
rect 45940 16646 46152 16674
rect 45836 12640 45888 12646
rect 45836 12582 45888 12588
rect 45744 12436 45796 12442
rect 45744 12378 45796 12384
rect 45848 12322 45876 12582
rect 45756 12306 45876 12322
rect 45744 12300 45876 12306
rect 45796 12294 45876 12300
rect 45744 12242 45796 12248
rect 45652 12232 45704 12238
rect 45652 12174 45704 12180
rect 45376 12164 45428 12170
rect 45376 12106 45428 12112
rect 45388 11218 45416 12106
rect 45560 11620 45612 11626
rect 45560 11562 45612 11568
rect 45572 11354 45600 11562
rect 45560 11348 45612 11354
rect 45560 11290 45612 11296
rect 45664 11286 45692 12174
rect 45756 11762 45784 12242
rect 45744 11756 45796 11762
rect 45744 11698 45796 11704
rect 45836 11756 45888 11762
rect 45836 11698 45888 11704
rect 45848 11354 45876 11698
rect 45836 11348 45888 11354
rect 45836 11290 45888 11296
rect 45652 11280 45704 11286
rect 45652 11222 45704 11228
rect 45376 11212 45428 11218
rect 45376 11154 45428 11160
rect 45388 10810 45416 11154
rect 45376 10804 45428 10810
rect 45376 10746 45428 10752
rect 45468 10668 45520 10674
rect 45468 10610 45520 10616
rect 45376 10600 45428 10606
rect 45376 10542 45428 10548
rect 45388 4690 45416 10542
rect 45480 9994 45508 10610
rect 45560 10532 45612 10538
rect 45560 10474 45612 10480
rect 45572 10062 45600 10474
rect 45664 10266 45692 11222
rect 45652 10260 45704 10266
rect 45652 10202 45704 10208
rect 45560 10056 45612 10062
rect 45560 9998 45612 10004
rect 45468 9988 45520 9994
rect 45468 9930 45520 9936
rect 45940 9674 45968 16646
rect 46020 16584 46072 16590
rect 46020 16526 46072 16532
rect 46032 12730 46060 16526
rect 46216 15094 46244 18022
rect 46204 15088 46256 15094
rect 46204 15030 46256 15036
rect 46308 14498 46336 18550
rect 46386 18456 46442 18465
rect 46386 18391 46442 18400
rect 46400 18290 46428 18391
rect 46388 18284 46440 18290
rect 46388 18226 46440 18232
rect 46492 16250 46520 20402
rect 46480 16244 46532 16250
rect 46480 16186 46532 16192
rect 46388 15496 46440 15502
rect 46388 15438 46440 15444
rect 46400 14822 46428 15438
rect 46388 14816 46440 14822
rect 46388 14758 46440 14764
rect 46584 14550 46612 20998
rect 46676 16182 46704 25978
rect 46860 25378 46888 31311
rect 47032 27872 47084 27878
rect 47032 27814 47084 27820
rect 47044 27538 47072 27814
rect 47032 27532 47084 27538
rect 47032 27474 47084 27480
rect 46768 25350 46888 25378
rect 46768 24954 46796 25350
rect 46846 25256 46902 25265
rect 46846 25191 46902 25200
rect 46756 24948 46808 24954
rect 46756 24890 46808 24896
rect 46860 24750 46888 25191
rect 46848 24744 46900 24750
rect 46848 24686 46900 24692
rect 46848 24608 46900 24614
rect 46848 24550 46900 24556
rect 46756 23724 46808 23730
rect 46756 23666 46808 23672
rect 46768 22778 46796 23666
rect 46756 22772 46808 22778
rect 46756 22714 46808 22720
rect 46768 22094 46796 22714
rect 46860 22642 46888 24550
rect 47136 23730 47164 33918
rect 47216 33924 47268 33930
rect 47216 33866 47268 33872
rect 47320 32178 47348 38898
rect 47504 32434 47532 41386
rect 47596 37874 47624 41942
rect 47768 41676 47820 41682
rect 47768 41618 47820 41624
rect 47780 41138 47808 41618
rect 48136 41608 48188 41614
rect 48134 41576 48136 41585
rect 48188 41576 48190 41585
rect 48134 41511 48190 41520
rect 47768 41132 47820 41138
rect 47768 41074 47820 41080
rect 48042 40896 48098 40905
rect 48042 40831 48098 40840
rect 47676 40520 47728 40526
rect 47676 40462 47728 40468
rect 47688 39574 47716 40462
rect 48056 40118 48084 40831
rect 48226 40216 48282 40225
rect 48226 40151 48282 40160
rect 48044 40112 48096 40118
rect 48044 40054 48096 40060
rect 47676 39568 47728 39574
rect 47676 39510 47728 39516
rect 48134 39536 48190 39545
rect 48240 39506 48268 40151
rect 48134 39471 48190 39480
rect 48228 39500 48280 39506
rect 47768 38956 47820 38962
rect 47768 38898 47820 38904
rect 47780 38865 47808 38898
rect 47766 38856 47822 38865
rect 47766 38791 47822 38800
rect 48148 38418 48176 39471
rect 48228 39442 48280 39448
rect 48136 38412 48188 38418
rect 48136 38354 48188 38360
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 47584 37868 47636 37874
rect 47584 37810 47636 37816
rect 47492 32428 47544 32434
rect 47492 32370 47544 32376
rect 47228 32150 47348 32178
rect 47228 28082 47256 32150
rect 47306 32056 47362 32065
rect 47306 31991 47362 32000
rect 47320 31822 47348 31991
rect 47308 31816 47360 31822
rect 47308 31758 47360 31764
rect 47308 29640 47360 29646
rect 47308 29582 47360 29588
rect 47400 29640 47452 29646
rect 47400 29582 47452 29588
rect 47320 29345 47348 29582
rect 47306 29336 47362 29345
rect 47306 29271 47362 29280
rect 47412 28626 47440 29582
rect 47400 28620 47452 28626
rect 47400 28562 47452 28568
rect 47216 28076 47268 28082
rect 47216 28018 47268 28024
rect 47228 25838 47256 28018
rect 47492 26920 47544 26926
rect 47492 26862 47544 26868
rect 47216 25832 47268 25838
rect 47216 25774 47268 25780
rect 47124 23724 47176 23730
rect 47124 23666 47176 23672
rect 46940 23112 46992 23118
rect 46940 23054 46992 23060
rect 46848 22636 46900 22642
rect 46848 22578 46900 22584
rect 46952 22098 46980 23054
rect 46768 22066 46888 22094
rect 46756 21956 46808 21962
rect 46756 21898 46808 21904
rect 46664 16176 46716 16182
rect 46664 16118 46716 16124
rect 46216 14470 46336 14498
rect 46572 14544 46624 14550
rect 46572 14486 46624 14492
rect 46664 14476 46716 14482
rect 46112 13320 46164 13326
rect 46112 13262 46164 13268
rect 46124 12850 46152 13262
rect 46112 12844 46164 12850
rect 46112 12786 46164 12792
rect 46032 12702 46152 12730
rect 46020 12640 46072 12646
rect 46020 12582 46072 12588
rect 46032 11082 46060 12582
rect 46124 12434 46152 12702
rect 46216 12646 46244 14470
rect 46664 14418 46716 14424
rect 46296 14408 46348 14414
rect 46296 14350 46348 14356
rect 46308 13938 46336 14350
rect 46480 14000 46532 14006
rect 46480 13942 46532 13948
rect 46296 13932 46348 13938
rect 46296 13874 46348 13880
rect 46308 12850 46336 13874
rect 46296 12844 46348 12850
rect 46296 12786 46348 12792
rect 46204 12640 46256 12646
rect 46204 12582 46256 12588
rect 46124 12406 46244 12434
rect 46020 11076 46072 11082
rect 46020 11018 46072 11024
rect 46112 10736 46164 10742
rect 46112 10678 46164 10684
rect 46124 9722 46152 10678
rect 46216 10606 46244 12406
rect 46492 12306 46520 13942
rect 46676 13530 46704 14418
rect 46664 13524 46716 13530
rect 46664 13466 46716 13472
rect 46480 12300 46532 12306
rect 46480 12242 46532 12248
rect 46768 11626 46796 21898
rect 46860 17202 46888 22066
rect 46940 22092 46992 22098
rect 46940 22034 46992 22040
rect 47124 22092 47176 22098
rect 47124 22034 47176 22040
rect 47032 19916 47084 19922
rect 47032 19858 47084 19864
rect 47044 18290 47072 19858
rect 47032 18284 47084 18290
rect 47032 18226 47084 18232
rect 47136 17270 47164 22034
rect 47124 17264 47176 17270
rect 47124 17206 47176 17212
rect 46848 17196 46900 17202
rect 46848 17138 46900 17144
rect 47032 16652 47084 16658
rect 47032 16594 47084 16600
rect 46940 16176 46992 16182
rect 46940 16118 46992 16124
rect 46848 14816 46900 14822
rect 46848 14758 46900 14764
rect 46860 13870 46888 14758
rect 46848 13864 46900 13870
rect 46848 13806 46900 13812
rect 46952 12434 46980 16118
rect 47044 16114 47072 16594
rect 47032 16108 47084 16114
rect 47032 16050 47084 16056
rect 47228 14346 47256 25774
rect 47504 24818 47532 26862
rect 47596 26042 47624 37810
rect 47676 37664 47728 37670
rect 47676 37606 47728 37612
rect 47688 37194 47716 37606
rect 48148 37330 48176 38111
rect 48136 37324 48188 37330
rect 48136 37266 48188 37272
rect 47676 37188 47728 37194
rect 47676 37130 47728 37136
rect 48136 35080 48188 35086
rect 48136 35022 48188 35028
rect 48148 34785 48176 35022
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48136 34604 48188 34610
rect 48136 34546 48188 34552
rect 48148 34105 48176 34546
rect 48134 34096 48190 34105
rect 48134 34031 48190 34040
rect 47860 33516 47912 33522
rect 47860 33458 47912 33464
rect 47872 33425 47900 33458
rect 47858 33416 47914 33425
rect 47858 33351 47914 33360
rect 47676 32836 47728 32842
rect 47676 32778 47728 32784
rect 48136 32836 48188 32842
rect 48136 32778 48188 32784
rect 47688 32570 47716 32778
rect 48148 32745 48176 32778
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 47676 32564 47728 32570
rect 47676 32506 47728 32512
rect 47676 32428 47728 32434
rect 47676 32370 47728 32376
rect 47688 31754 47716 32370
rect 47688 31726 47808 31754
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 47688 27402 47716 27814
rect 47676 27396 47728 27402
rect 47676 27338 47728 27344
rect 47584 26036 47636 26042
rect 47584 25978 47636 25984
rect 47676 25220 47728 25226
rect 47676 25162 47728 25168
rect 47688 24818 47716 25162
rect 47492 24812 47544 24818
rect 47492 24754 47544 24760
rect 47676 24812 47728 24818
rect 47676 24754 47728 24760
rect 47306 23216 47362 23225
rect 47306 23151 47308 23160
rect 47360 23151 47362 23160
rect 47308 23122 47360 23128
rect 47504 22094 47532 24754
rect 47676 24132 47728 24138
rect 47676 24074 47728 24080
rect 47688 23866 47716 24074
rect 47676 23860 47728 23866
rect 47676 23802 47728 23808
rect 47584 23724 47636 23730
rect 47584 23666 47636 23672
rect 47412 22066 47532 22094
rect 47308 20800 47360 20806
rect 47308 20742 47360 20748
rect 47320 18834 47348 20742
rect 47412 18902 47440 22066
rect 47400 18896 47452 18902
rect 47400 18838 47452 18844
rect 47308 18828 47360 18834
rect 47308 18770 47360 18776
rect 47216 14340 47268 14346
rect 47216 14282 47268 14288
rect 47228 13938 47256 14282
rect 47216 13932 47268 13938
rect 47216 13874 47268 13880
rect 47320 13682 47348 18770
rect 47596 18290 47624 23666
rect 47780 22778 47808 31726
rect 47860 28620 47912 28626
rect 47860 28562 47912 28568
rect 47872 28218 47900 28562
rect 47860 28212 47912 28218
rect 47860 28154 47912 28160
rect 47768 22772 47820 22778
rect 47768 22714 47820 22720
rect 47768 22094 47820 22098
rect 47872 22094 47900 28154
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48042 26616 48098 26625
rect 48042 26551 48098 26560
rect 48056 26450 48084 26551
rect 48044 26444 48096 26450
rect 48044 26386 48096 26392
rect 48134 25936 48190 25945
rect 48134 25871 48190 25880
rect 48148 25362 48176 25871
rect 48136 25356 48188 25362
rect 48136 25298 48188 25304
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48148 24274 48176 24511
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 47768 22092 47900 22094
rect 47820 22066 47900 22092
rect 47768 22034 47820 22040
rect 47950 21856 48006 21865
rect 47950 21791 48006 21800
rect 47964 21622 47992 21791
rect 47952 21616 48004 21622
rect 47952 21558 48004 21564
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 47768 21004 47820 21010
rect 47768 20946 47820 20952
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 47780 20466 47808 20946
rect 47768 20460 47820 20466
rect 47768 20402 47820 20408
rect 47676 19780 47728 19786
rect 47676 19722 47728 19728
rect 48136 19780 48188 19786
rect 48136 19722 48188 19728
rect 47688 18426 47716 19722
rect 48148 19145 48176 19722
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 47676 18420 47728 18426
rect 47676 18362 47728 18368
rect 47584 18284 47636 18290
rect 47584 18226 47636 18232
rect 47400 17196 47452 17202
rect 47400 17138 47452 17144
rect 47136 13654 47348 13682
rect 46952 12406 47072 12434
rect 46756 11620 46808 11626
rect 46756 11562 46808 11568
rect 46204 10600 46256 10606
rect 46204 10542 46256 10548
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46308 10130 46336 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 45848 9646 45968 9674
rect 46112 9716 46164 9722
rect 46112 9658 46164 9664
rect 45560 8288 45612 8294
rect 45558 8256 45560 8265
rect 45612 8256 45614 8265
rect 45558 8191 45614 8200
rect 45376 4684 45428 4690
rect 45296 4644 45376 4672
rect 45192 4548 45244 4554
rect 45192 4490 45244 4496
rect 45296 4282 45324 4644
rect 45376 4626 45428 4632
rect 45744 4480 45796 4486
rect 45744 4422 45796 4428
rect 45284 4276 45336 4282
rect 45284 4218 45336 4224
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 45204 3058 45232 3470
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 45296 2582 45324 4218
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45388 3126 45416 3334
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 45284 2576 45336 2582
rect 45284 2518 45336 2524
rect 45756 2514 45784 4422
rect 45848 3738 45876 9646
rect 46846 9616 46902 9625
rect 46846 9551 46848 9560
rect 46900 9551 46902 9560
rect 46848 9522 46900 9528
rect 46846 6216 46902 6225
rect 46846 6151 46902 6160
rect 46860 5778 46888 6151
rect 46848 5772 46900 5778
rect 46848 5714 46900 5720
rect 46848 5228 46900 5234
rect 46848 5170 46900 5176
rect 46388 4820 46440 4826
rect 46388 4762 46440 4768
rect 46400 4622 46428 4762
rect 46388 4616 46440 4622
rect 46388 4558 46440 4564
rect 46480 4480 46532 4486
rect 46480 4422 46532 4428
rect 46388 4208 46440 4214
rect 46388 4150 46440 4156
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 45836 3732 45888 3738
rect 45836 3674 45888 3680
rect 45848 2514 45876 3674
rect 46308 3602 46336 3878
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 45100 2508 45152 2514
rect 45100 2450 45152 2456
rect 45744 2508 45796 2514
rect 45744 2450 45796 2456
rect 45836 2508 45888 2514
rect 45836 2450 45888 2456
rect 45468 2372 45520 2378
rect 45468 2314 45520 2320
rect 45020 1822 45140 1850
rect 45112 800 45140 1822
rect 30484 734 30788 762
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45480 354 45508 2314
rect 46400 800 46428 4150
rect 46492 3602 46520 4422
rect 46860 4185 46888 5170
rect 47044 4570 47072 12406
rect 47136 8022 47164 13654
rect 47216 13388 47268 13394
rect 47216 13330 47268 13336
rect 47228 12850 47256 13330
rect 47216 12844 47268 12850
rect 47216 12786 47268 12792
rect 47124 8016 47176 8022
rect 47124 7958 47176 7964
rect 47124 7200 47176 7206
rect 47124 7142 47176 7148
rect 47136 6866 47164 7142
rect 47124 6860 47176 6866
rect 47124 6802 47176 6808
rect 47228 5710 47256 12786
rect 47412 12434 47440 17138
rect 47412 12406 47532 12434
rect 47504 9586 47532 12406
rect 47492 9580 47544 9586
rect 47492 9522 47544 9528
rect 47308 8968 47360 8974
rect 47308 8910 47360 8916
rect 47400 8968 47452 8974
rect 47400 8910 47452 8916
rect 47320 7585 47348 8910
rect 47412 7954 47440 8910
rect 47400 7948 47452 7954
rect 47400 7890 47452 7896
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47216 5704 47268 5710
rect 47216 5646 47268 5652
rect 47216 5024 47268 5030
rect 47216 4966 47268 4972
rect 46952 4542 47072 4570
rect 47228 4554 47256 4966
rect 47216 4548 47268 4554
rect 46846 4176 46902 4185
rect 46846 4111 46902 4120
rect 46662 4040 46718 4049
rect 46662 3975 46718 3984
rect 46676 3942 46704 3975
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 46952 2990 46980 4542
rect 47216 4490 47268 4496
rect 47032 4480 47084 4486
rect 47032 4422 47084 4428
rect 46940 2984 46992 2990
rect 46940 2926 46992 2932
rect 47044 800 47072 4422
rect 47504 3670 47532 9522
rect 47596 4826 47624 18226
rect 47676 17604 47728 17610
rect 47676 17546 47728 17552
rect 48136 17604 48188 17610
rect 48136 17546 48188 17552
rect 47688 17338 47716 17546
rect 47676 17332 47728 17338
rect 47676 17274 47728 17280
rect 48148 17105 48176 17546
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 48136 16516 48188 16522
rect 48136 16458 48188 16464
rect 47688 16250 47716 16458
rect 48148 16425 48176 16458
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 47676 16244 47728 16250
rect 47676 16186 47728 16192
rect 47860 15496 47912 15502
rect 47912 15444 47992 15450
rect 47860 15438 47992 15444
rect 47872 15422 47992 15438
rect 47860 15360 47912 15366
rect 47860 15302 47912 15308
rect 47768 15088 47820 15094
rect 47768 15030 47820 15036
rect 47676 15020 47728 15026
rect 47676 14962 47728 14968
rect 47688 14414 47716 14962
rect 47780 14550 47808 15030
rect 47768 14544 47820 14550
rect 47768 14486 47820 14492
rect 47676 14408 47728 14414
rect 47676 14350 47728 14356
rect 47872 14278 47900 15302
rect 47964 14822 47992 15422
rect 47952 14816 48004 14822
rect 47952 14758 48004 14764
rect 47860 14272 47912 14278
rect 47860 14214 47912 14220
rect 47872 13870 47900 14214
rect 47964 14074 47992 14758
rect 48228 14340 48280 14346
rect 48228 14282 48280 14288
rect 47952 14068 48004 14074
rect 47952 14010 48004 14016
rect 47860 13864 47912 13870
rect 47860 13806 47912 13812
rect 47676 13320 47728 13326
rect 47676 13262 47728 13268
rect 47688 12374 47716 13262
rect 47676 12368 47728 12374
rect 47676 12310 47728 12316
rect 48134 12336 48190 12345
rect 48134 12271 48136 12280
rect 48188 12271 48190 12280
rect 48136 12242 48188 12248
rect 47768 11552 47820 11558
rect 47768 11494 47820 11500
rect 47780 11218 47808 11494
rect 47768 11212 47820 11218
rect 47768 11154 47820 11160
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 47676 9988 47728 9994
rect 47676 9930 47728 9936
rect 47688 9654 47716 9930
rect 47676 9648 47728 9654
rect 47676 9590 47728 9596
rect 47766 8936 47822 8945
rect 47766 8871 47822 8880
rect 47780 8566 47808 8871
rect 47768 8560 47820 8566
rect 47768 8502 47820 8508
rect 47676 7948 47728 7954
rect 47676 7890 47728 7896
rect 47584 4820 47636 4826
rect 47584 4762 47636 4768
rect 47492 3664 47544 3670
rect 47492 3606 47544 3612
rect 47688 3466 47716 7890
rect 48136 7404 48188 7410
rect 48136 7346 48188 7352
rect 48148 6905 48176 7346
rect 48134 6896 48190 6905
rect 48240 6866 48268 14282
rect 48134 6831 48190 6840
rect 48228 6860 48280 6866
rect 48228 6802 48280 6808
rect 48240 4690 48268 6802
rect 48320 5228 48372 5234
rect 48320 5170 48372 5176
rect 48228 4684 48280 4690
rect 48228 4626 48280 4632
rect 47768 4208 47820 4214
rect 47768 4150 47820 4156
rect 47780 3505 47808 4150
rect 47766 3496 47822 3505
rect 47676 3460 47728 3466
rect 47766 3431 47822 3440
rect 47676 3402 47728 3408
rect 47768 3052 47820 3058
rect 47768 2994 47820 3000
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47688 800 47716 2926
rect 47780 1465 47808 2994
rect 47952 2372 48004 2378
rect 47952 2314 48004 2320
rect 47766 1456 47822 1465
rect 47766 1391 47822 1400
rect 45558 776 45614 785
rect 45558 711 45614 720
rect 45572 354 45600 711
rect 45480 326 45600 354
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 47964 105 47992 2314
rect 48332 800 48360 5170
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48976 800 49004 3402
rect 47950 96 48006 105
rect 47950 31 48006 40
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1398 47640 1454 47696
rect 3422 46960 3478 47016
rect 1398 40160 1454 40216
rect 1398 33396 1400 33416
rect 1400 33396 1452 33416
rect 1452 33396 1454 33416
rect 1398 33360 1454 33396
rect 1582 35400 1638 35456
rect 1306 32680 1362 32736
rect 1858 42880 1914 42936
rect 1858 41520 1914 41576
rect 2778 46280 2834 46336
rect 1858 32000 1914 32056
rect 1398 25236 1400 25256
rect 1400 25236 1452 25256
rect 1452 25236 1454 25256
rect 1398 25200 1454 25236
rect 1398 12280 1454 12336
rect 1858 23160 1914 23216
rect 1858 17720 1914 17776
rect 1858 16360 1914 16416
rect 2226 19080 2282 19136
rect 2962 44920 3018 44976
rect 2778 36760 2834 36816
rect 3330 28600 3386 28656
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3514 43560 3570 43616
rect 3698 39480 3754 39536
rect 3606 31320 3662 31376
rect 3330 17076 3332 17096
rect 3332 17076 3384 17096
rect 3384 17076 3386 17096
rect 3330 17040 3386 17076
rect 2778 15000 2834 15056
rect 2962 7520 3018 7576
rect 3974 19760 4030 19816
rect 3974 18400 4030 18456
rect 3974 13676 3976 13696
rect 3976 13676 4028 13696
rect 4028 13676 4030 13696
rect 3974 13640 4030 13676
rect 3514 10240 3570 10296
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3514 6860 3570 6896
rect 3514 6840 3516 6860
rect 3516 6840 3568 6860
rect 3568 6840 3570 6860
rect 3422 3440 3478 3496
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3974 3576 4030 3632
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3514 1400 3570 1456
rect 2870 720 2926 776
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 17130 3460 17186 3496
rect 17130 3440 17132 3460
rect 17132 3440 17184 3460
rect 17184 3440 17186 3460
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 20626 32408 20682 32464
rect 20994 30232 21050 30288
rect 20534 23060 20536 23080
rect 20536 23060 20588 23080
rect 20588 23060 20590 23080
rect 20534 23024 20590 23060
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21454 33940 21456 33960
rect 21456 33940 21508 33960
rect 21508 33940 21510 33960
rect 21454 33904 21510 33940
rect 21270 30368 21326 30424
rect 21546 30232 21602 30288
rect 22558 36252 22560 36272
rect 22560 36252 22612 36272
rect 22612 36252 22614 36272
rect 22558 36216 22614 36252
rect 23386 36352 23442 36408
rect 22650 34196 22706 34232
rect 22650 34176 22652 34196
rect 22652 34176 22704 34196
rect 22704 34176 22706 34196
rect 22282 32272 22338 32328
rect 22190 30368 22246 30424
rect 21362 23180 21418 23216
rect 21362 23160 21364 23180
rect 21364 23160 21416 23180
rect 21416 23160 21418 23180
rect 23938 36352 23994 36408
rect 21914 3984 21970 4040
rect 23386 19760 23442 19816
rect 25042 32408 25098 32464
rect 26238 34176 26294 34232
rect 25594 32272 25650 32328
rect 27802 36252 27804 36272
rect 27804 36252 27856 36272
rect 27856 36252 27858 36272
rect 27802 36216 27858 36252
rect 27710 33904 27766 33960
rect 27434 27920 27490 27976
rect 28170 27784 28226 27840
rect 27342 23180 27398 23216
rect 27342 23160 27344 23180
rect 27344 23160 27396 23180
rect 27396 23160 27398 23180
rect 28446 27548 28448 27568
rect 28448 27548 28500 27568
rect 28500 27548 28502 27568
rect 28446 27512 28502 27548
rect 28906 27940 28962 27976
rect 28906 27920 28908 27940
rect 28908 27920 28960 27940
rect 28960 27920 28962 27940
rect 28906 27784 28962 27840
rect 28814 27548 28816 27568
rect 28816 27548 28868 27568
rect 28868 27548 28870 27568
rect 28814 27512 28870 27548
rect 28906 23060 28908 23080
rect 28908 23060 28960 23080
rect 28960 23060 28962 23080
rect 28906 23024 28962 23060
rect 29550 3596 29606 3632
rect 29550 3576 29552 3596
rect 29552 3576 29604 3596
rect 29604 3576 29606 3596
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 39118 3032 39174 3088
rect 40130 3032 40186 3088
rect 45558 28600 45614 28656
rect 45558 23840 45614 23896
rect 46846 47640 46902 47696
rect 47858 46280 47914 46336
rect 48134 45600 48190 45656
rect 45466 15680 45522 15736
rect 44914 3440 44970 3496
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 46846 31320 46902 31376
rect 46754 29960 46810 30016
rect 46570 22516 46572 22536
rect 46572 22516 46624 22536
rect 46624 22516 46626 22536
rect 46570 22480 46626 22516
rect 46386 18400 46442 18456
rect 46846 25200 46902 25256
rect 48134 41556 48136 41576
rect 48136 41556 48188 41576
rect 48188 41556 48190 41576
rect 48134 41520 48190 41556
rect 48042 40840 48098 40896
rect 48226 40160 48282 40216
rect 48134 39480 48190 39536
rect 47766 38800 47822 38856
rect 48134 38120 48190 38176
rect 47306 32000 47362 32056
rect 47306 29280 47362 29336
rect 48134 34720 48190 34776
rect 48134 34040 48190 34096
rect 47858 33360 47914 33416
rect 48134 32680 48190 32736
rect 47306 23180 47362 23216
rect 47306 23160 47308 23180
rect 47308 23160 47360 23180
rect 47360 23160 47362 23180
rect 48134 27920 48190 27976
rect 48042 26560 48098 26616
rect 48134 25880 48190 25936
rect 48134 24520 48190 24576
rect 47950 21800 48006 21856
rect 48134 21120 48190 21176
rect 48134 19080 48190 19136
rect 45558 8236 45560 8256
rect 45560 8236 45612 8256
rect 45612 8236 45614 8256
rect 45558 8200 45614 8236
rect 46846 9580 46902 9616
rect 46846 9560 46848 9580
rect 46848 9560 46900 9580
rect 46900 9560 46902 9580
rect 46846 6160 46902 6216
rect 47306 7520 47362 7576
rect 46846 4120 46902 4176
rect 46662 3984 46718 4040
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 12300 48190 12336
rect 48134 12280 48136 12300
rect 48136 12280 48188 12300
rect 48188 12280 48190 12300
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 47766 8880 47822 8936
rect 48134 6840 48190 6896
rect 47766 3440 47822 3496
rect 47766 1400 47822 1456
rect 45558 720 45614 776
rect 47950 40 48006 96
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1393 47698 1459 47701
rect 0 47696 1459 47698
rect 0 47640 1398 47696
rect 1454 47640 1459 47696
rect 0 47638 1459 47640
rect 0 47548 800 47638
rect 1393 47635 1459 47638
rect 46841 47698 46907 47701
rect 49200 47698 50000 47788
rect 46841 47696 50000 47698
rect 46841 47640 46846 47696
rect 46902 47640 50000 47696
rect 46841 47638 50000 47640
rect 46841 47635 46907 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3417 47018 3483 47021
rect 0 47016 3483 47018
rect 0 46960 3422 47016
rect 3478 46960 3483 47016
rect 0 46958 3483 46960
rect 0 46868 800 46958
rect 3417 46955 3483 46958
rect 46054 46956 46060 47020
rect 46124 47018 46130 47020
rect 49200 47018 50000 47108
rect 46124 46958 50000 47018
rect 46124 46956 46130 46958
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46188 800 46278
rect 2773 46275 2839 46278
rect 47853 46338 47919 46341
rect 49200 46338 50000 46428
rect 47853 46336 50000 46338
rect 47853 46280 47858 46336
rect 47914 46280 50000 46336
rect 47853 46278 50000 46280
rect 47853 46275 47919 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 2957 44978 3023 44981
rect 0 44976 3023 44978
rect 0 44920 2962 44976
rect 3018 44920 3023 44976
rect 0 44918 3023 44920
rect 0 44828 800 44918
rect 2957 44915 3023 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3509 43618 3575 43621
rect 0 43616 3575 43618
rect 0 43560 3514 43616
rect 3570 43560 3575 43616
rect 0 43558 3575 43560
rect 0 43468 800 43558
rect 3509 43555 3575 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1853 42938 1919 42941
rect 0 42936 1919 42938
rect 0 42880 1858 42936
rect 1914 42880 1919 42936
rect 0 42878 1919 42880
rect 0 42788 800 42878
rect 1853 42875 1919 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 48037 40898 48103 40901
rect 49200 40898 50000 40988
rect 48037 40896 50000 40898
rect 48037 40840 48042 40896
rect 48098 40840 50000 40896
rect 48037 40838 50000 40840
rect 48037 40835 48103 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1393 40218 1459 40221
rect 0 40216 1459 40218
rect 0 40160 1398 40216
rect 1454 40160 1459 40216
rect 0 40158 1459 40160
rect 0 40068 800 40158
rect 1393 40155 1459 40158
rect 48221 40218 48287 40221
rect 49200 40218 50000 40308
rect 48221 40216 50000 40218
rect 48221 40160 48226 40216
rect 48282 40160 50000 40216
rect 48221 40158 50000 40160
rect 48221 40155 48287 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3693 39538 3759 39541
rect 0 39536 3759 39538
rect 0 39480 3698 39536
rect 3754 39480 3759 39536
rect 0 39478 3759 39480
rect 0 39388 800 39478
rect 3693 39475 3759 39478
rect 48129 39538 48195 39541
rect 49200 39538 50000 39628
rect 48129 39536 50000 39538
rect 48129 39480 48134 39536
rect 48190 39480 50000 39536
rect 48129 39478 50000 39480
rect 48129 39475 48195 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47761 38858 47827 38861
rect 49200 38858 50000 38948
rect 47761 38856 50000 38858
rect 47761 38800 47766 38856
rect 47822 38800 50000 38856
rect 47761 38798 50000 38800
rect 47761 38795 47827 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 23381 36410 23447 36413
rect 23933 36410 23999 36413
rect 23381 36408 23999 36410
rect 23381 36352 23386 36408
rect 23442 36352 23938 36408
rect 23994 36352 23999 36408
rect 23381 36350 23999 36352
rect 23381 36347 23447 36350
rect 23933 36347 23999 36350
rect 22553 36274 22619 36277
rect 27797 36274 27863 36277
rect 22553 36272 27863 36274
rect 0 35988 800 36228
rect 22553 36216 22558 36272
rect 22614 36216 27802 36272
rect 27858 36216 27863 36272
rect 22553 36214 27863 36216
rect 22553 36211 22619 36214
rect 27797 36211 27863 36214
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35458 800 35548
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 22645 34234 22711 34237
rect 26233 34234 26299 34237
rect 22645 34232 26299 34234
rect 0 33948 800 34188
rect 22645 34176 22650 34232
rect 22706 34176 26238 34232
rect 26294 34176 26299 34232
rect 22645 34174 26299 34176
rect 22645 34171 22711 34174
rect 26233 34171 26299 34174
rect 48129 34098 48195 34101
rect 49200 34098 50000 34188
rect 48129 34096 50000 34098
rect 48129 34040 48134 34096
rect 48190 34040 50000 34096
rect 48129 34038 50000 34040
rect 48129 34035 48195 34038
rect 21449 33962 21515 33965
rect 27705 33962 27771 33965
rect 21449 33960 27771 33962
rect 21449 33904 21454 33960
rect 21510 33904 27710 33960
rect 27766 33904 27771 33960
rect 49200 33948 50000 34038
rect 21449 33902 27771 33904
rect 21449 33899 21515 33902
rect 27705 33899 27771 33902
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 47853 33418 47919 33421
rect 49200 33418 50000 33508
rect 47853 33416 50000 33418
rect 47853 33360 47858 33416
rect 47914 33360 50000 33416
rect 47853 33358 50000 33360
rect 47853 33355 47919 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32828
rect 1301 32738 1367 32741
rect 0 32736 1367 32738
rect 0 32680 1306 32736
rect 1362 32680 1367 32736
rect 0 32678 1367 32680
rect 0 32588 800 32678
rect 1301 32675 1367 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 49200 32588 50000 32678
rect 20621 32466 20687 32469
rect 25037 32466 25103 32469
rect 20621 32464 25103 32466
rect 20621 32408 20626 32464
rect 20682 32408 25042 32464
rect 25098 32408 25103 32464
rect 20621 32406 25103 32408
rect 20621 32403 20687 32406
rect 25037 32403 25103 32406
rect 22277 32330 22343 32333
rect 25589 32330 25655 32333
rect 22277 32328 25655 32330
rect 22277 32272 22282 32328
rect 22338 32272 25594 32328
rect 25650 32272 25655 32328
rect 22277 32270 25655 32272
rect 22277 32267 22343 32270
rect 25589 32267 25655 32270
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 1853 32058 1919 32061
rect 0 32056 1919 32058
rect 0 32000 1858 32056
rect 1914 32000 1919 32056
rect 0 31998 1919 32000
rect 0 31908 800 31998
rect 1853 31995 1919 31998
rect 47301 32058 47367 32061
rect 49200 32058 50000 32148
rect 47301 32056 50000 32058
rect 47301 32000 47306 32056
rect 47362 32000 50000 32056
rect 47301 31998 50000 32000
rect 47301 31995 47367 31998
rect 49200 31908 50000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3601 31378 3667 31381
rect 0 31376 3667 31378
rect 0 31320 3606 31376
rect 3662 31320 3667 31376
rect 0 31318 3667 31320
rect 0 31228 800 31318
rect 3601 31315 3667 31318
rect 46841 31378 46907 31381
rect 49200 31378 50000 31468
rect 46841 31376 50000 31378
rect 46841 31320 46846 31376
rect 46902 31320 50000 31376
rect 46841 31318 50000 31320
rect 46841 31315 46907 31318
rect 49200 31228 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 21265 30426 21331 30429
rect 22185 30426 22251 30429
rect 21265 30424 22251 30426
rect 21265 30368 21270 30424
rect 21326 30368 22190 30424
rect 22246 30368 22251 30424
rect 21265 30366 22251 30368
rect 21265 30363 21331 30366
rect 22185 30363 22251 30366
rect 20989 30290 21055 30293
rect 21541 30290 21607 30293
rect 20989 30288 21607 30290
rect 20989 30232 20994 30288
rect 21050 30232 21546 30288
rect 21602 30232 21607 30288
rect 20989 30230 21607 30232
rect 20989 30227 21055 30230
rect 21541 30227 21607 30230
rect 0 29868 800 30108
rect 46749 30018 46815 30021
rect 49200 30018 50000 30108
rect 46749 30016 50000 30018
rect 46749 29960 46754 30016
rect 46810 29960 50000 30016
rect 46749 29958 50000 29960
rect 46749 29955 46815 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 47301 29338 47367 29341
rect 49200 29338 50000 29428
rect 47301 29336 50000 29338
rect 47301 29280 47306 29336
rect 47362 29280 50000 29336
rect 47301 29278 50000 29280
rect 47301 29275 47367 29278
rect 49200 29188 50000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3325 28658 3391 28661
rect 0 28656 3391 28658
rect 0 28600 3330 28656
rect 3386 28600 3391 28656
rect 0 28598 3391 28600
rect 0 28508 800 28598
rect 3325 28595 3391 28598
rect 45553 28658 45619 28661
rect 49200 28658 50000 28748
rect 45553 28656 50000 28658
rect 45553 28600 45558 28656
rect 45614 28600 50000 28656
rect 45553 28598 50000 28600
rect 45553 28595 45619 28598
rect 49200 28508 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 27429 27978 27495 27981
rect 28901 27978 28967 27981
rect 27429 27976 28967 27978
rect 27429 27920 27434 27976
rect 27490 27920 28906 27976
rect 28962 27920 28967 27976
rect 27429 27918 28967 27920
rect 27429 27915 27495 27918
rect 28901 27915 28967 27918
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 28165 27842 28231 27845
rect 28901 27842 28967 27845
rect 28165 27840 28967 27842
rect 28165 27784 28170 27840
rect 28226 27784 28906 27840
rect 28962 27784 28967 27840
rect 49200 27828 50000 27918
rect 28165 27782 28967 27784
rect 28165 27779 28231 27782
rect 28901 27779 28967 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 28441 27570 28507 27573
rect 28809 27570 28875 27573
rect 28441 27568 28875 27570
rect 28441 27512 28446 27568
rect 28502 27512 28814 27568
rect 28870 27512 28875 27568
rect 28441 27510 28875 27512
rect 28441 27507 28507 27510
rect 28809 27507 28875 27510
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 48037 26618 48103 26621
rect 49200 26618 50000 26708
rect 48037 26616 50000 26618
rect 48037 26560 48042 26616
rect 48098 26560 50000 26616
rect 48037 26558 50000 26560
rect 48037 26555 48103 26558
rect 49200 26468 50000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 48129 25938 48195 25941
rect 49200 25938 50000 26028
rect 48129 25936 50000 25938
rect 48129 25880 48134 25936
rect 48190 25880 50000 25936
rect 48129 25878 50000 25880
rect 48129 25875 48195 25878
rect 49200 25788 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25108 800 25198
rect 1393 25195 1459 25198
rect 46841 25258 46907 25261
rect 49200 25258 50000 25348
rect 46841 25256 50000 25258
rect 46841 25200 46846 25256
rect 46902 25200 50000 25256
rect 46841 25198 50000 25200
rect 46841 25195 46907 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24428 800 24668
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 45553 23898 45619 23901
rect 49200 23898 50000 23988
rect 45553 23896 50000 23898
rect 45553 23840 45558 23896
rect 45614 23840 50000 23896
rect 45553 23838 50000 23840
rect 45553 23835 45619 23838
rect 49200 23748 50000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23068 800 23158
rect 1853 23155 1919 23158
rect 21357 23218 21423 23221
rect 27337 23218 27403 23221
rect 21357 23216 27403 23218
rect 21357 23160 21362 23216
rect 21418 23160 27342 23216
rect 27398 23160 27403 23216
rect 21357 23158 27403 23160
rect 21357 23155 21423 23158
rect 27337 23155 27403 23158
rect 47301 23218 47367 23221
rect 49200 23218 50000 23308
rect 47301 23216 50000 23218
rect 47301 23160 47306 23216
rect 47362 23160 50000 23216
rect 47301 23158 50000 23160
rect 47301 23155 47367 23158
rect 20529 23082 20595 23085
rect 28901 23082 28967 23085
rect 20529 23080 28967 23082
rect 20529 23024 20534 23080
rect 20590 23024 28906 23080
rect 28962 23024 28967 23080
rect 49200 23068 50000 23158
rect 20529 23022 28967 23024
rect 20529 23019 20595 23022
rect 28901 23019 28967 23022
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 46565 22538 46631 22541
rect 49200 22538 50000 22628
rect 46565 22536 50000 22538
rect 46565 22480 46570 22536
rect 46626 22480 50000 22536
rect 46565 22478 50000 22480
rect 46565 22475 46631 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21708 800 21948
rect 47945 21858 48011 21861
rect 49200 21858 50000 21948
rect 47945 21856 50000 21858
rect 47945 21800 47950 21856
rect 48006 21800 50000 21856
rect 47945 21798 50000 21800
rect 47945 21795 48011 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 49200 21028 50000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19668 800 19758
rect 3969 19755 4035 19758
rect 23381 19818 23447 19821
rect 46054 19818 46060 19820
rect 23381 19816 46060 19818
rect 23381 19760 23386 19816
rect 23442 19760 46060 19816
rect 23381 19758 46060 19760
rect 23381 19755 23447 19758
rect 46054 19756 46060 19758
rect 46124 19756 46130 19820
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3969 18458 4035 18461
rect 0 18456 4035 18458
rect 0 18400 3974 18456
rect 4030 18400 4035 18456
rect 0 18398 4035 18400
rect 0 18308 800 18398
rect 3969 18395 4035 18398
rect 46381 18458 46447 18461
rect 49200 18458 50000 18548
rect 46381 18456 50000 18458
rect 46381 18400 46386 18456
rect 46442 18400 50000 18456
rect 46381 18398 50000 18400
rect 46381 18395 46447 18398
rect 49200 18308 50000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1853 17778 1919 17781
rect 0 17776 1919 17778
rect 0 17720 1858 17776
rect 1914 17720 1919 17776
rect 0 17718 1919 17720
rect 0 17628 800 17718
rect 1853 17715 1919 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3325 17098 3391 17101
rect 0 17096 3391 17098
rect 0 17040 3330 17096
rect 3386 17040 3391 17096
rect 0 17038 3391 17040
rect 0 16948 800 17038
rect 3325 17035 3391 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16268 800 16358
rect 1853 16355 1919 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16508
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 45461 15738 45527 15741
rect 49200 15738 50000 15828
rect 45461 15736 50000 15738
rect 45461 15680 45466 15736
rect 45522 15680 50000 15736
rect 45461 15678 50000 15680
rect 45461 15675 45527 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3969 13698 4035 13701
rect 0 13696 4035 13698
rect 0 13640 3974 13696
rect 4030 13640 4035 13696
rect 0 13638 4035 13640
rect 0 13548 800 13638
rect 3969 13635 4035 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 3509 10298 3575 10301
rect 0 10296 3575 10298
rect 0 10240 3514 10296
rect 3570 10240 3575 10296
rect 0 10238 3575 10240
rect 0 10148 800 10238
rect 3509 10235 3575 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 46841 9618 46907 9621
rect 49200 9618 50000 9708
rect 46841 9616 50000 9618
rect 46841 9560 46846 9616
rect 46902 9560 50000 9616
rect 46841 9558 50000 9560
rect 46841 9555 46907 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47761 8938 47827 8941
rect 49200 8938 50000 9028
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 45553 8258 45619 8261
rect 49200 8258 50000 8348
rect 45553 8256 50000 8258
rect 45553 8200 45558 8256
rect 45614 8200 50000 8256
rect 45553 8198 50000 8200
rect 45553 8195 45619 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 2957 7578 3023 7581
rect 0 7576 3023 7578
rect 0 7520 2962 7576
rect 3018 7520 3023 7576
rect 0 7518 3023 7520
rect 0 7428 800 7518
rect 2957 7515 3023 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 3509 6898 3575 6901
rect 0 6896 3575 6898
rect 0 6840 3514 6896
rect 3570 6840 3575 6896
rect 0 6838 3575 6840
rect 0 6748 800 6838
rect 3509 6835 3575 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 46841 6218 46907 6221
rect 49200 6218 50000 6308
rect 46841 6216 50000 6218
rect 46841 6160 46846 6216
rect 46902 6160 50000 6216
rect 46841 6158 50000 6160
rect 46841 6155 46907 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 46841 4178 46907 4181
rect 49200 4178 50000 4268
rect 46841 4176 50000 4178
rect 46841 4120 46846 4176
rect 46902 4120 50000 4176
rect 46841 4118 50000 4120
rect 46841 4115 46907 4118
rect 21909 4042 21975 4045
rect 46657 4042 46723 4045
rect 21909 4040 46723 4042
rect 21909 3984 21914 4040
rect 21970 3984 46662 4040
rect 46718 3984 46723 4040
rect 49200 4028 50000 4118
rect 21909 3982 46723 3984
rect 21909 3979 21975 3982
rect 46657 3979 46723 3982
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 3969 3634 4035 3637
rect 29545 3634 29611 3637
rect 3969 3632 29611 3634
rect 0 3498 800 3588
rect 3969 3576 3974 3632
rect 4030 3576 29550 3632
rect 29606 3576 29611 3632
rect 3969 3574 29611 3576
rect 3969 3571 4035 3574
rect 29545 3571 29611 3574
rect 3417 3498 3483 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3348 800 3438
rect 3417 3435 3483 3438
rect 17125 3498 17191 3501
rect 44909 3498 44975 3501
rect 17125 3496 44975 3498
rect 17125 3440 17130 3496
rect 17186 3440 44914 3496
rect 44970 3440 44975 3496
rect 17125 3438 44975 3440
rect 17125 3435 17191 3438
rect 44909 3435 44975 3438
rect 47761 3498 47827 3501
rect 49200 3498 50000 3588
rect 47761 3496 50000 3498
rect 47761 3440 47766 3496
rect 47822 3440 50000 3496
rect 47761 3438 50000 3440
rect 47761 3435 47827 3438
rect 49200 3348 50000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 39113 3090 39179 3093
rect 40125 3090 40191 3093
rect 39113 3088 40191 3090
rect 39113 3032 39118 3088
rect 39174 3032 40130 3088
rect 40186 3032 40191 3088
rect 39113 3030 40191 3032
rect 39113 3027 39179 3030
rect 40125 3027 40191 3030
rect 0 2668 800 2908
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3509 1458 3575 1461
rect 0 1456 3575 1458
rect 0 1400 3514 1456
rect 3570 1400 3575 1456
rect 0 1398 3575 1400
rect 0 1308 800 1398
rect 3509 1395 3575 1398
rect 47761 1458 47827 1461
rect 49200 1458 50000 1548
rect 47761 1456 50000 1458
rect 47761 1400 47766 1456
rect 47822 1400 50000 1456
rect 47761 1398 50000 1400
rect 47761 1395 47827 1398
rect 49200 1308 50000 1398
rect 0 778 800 868
rect 2865 778 2931 781
rect 0 776 2931 778
rect 0 720 2870 776
rect 2926 720 2931 776
rect 0 718 2931 720
rect 0 628 800 718
rect 2865 715 2931 718
rect 45553 778 45619 781
rect 49200 778 50000 868
rect 45553 776 50000 778
rect 45553 720 45558 776
rect 45614 720 50000 776
rect 45553 718 50000 720
rect 45553 715 45619 718
rect 49200 628 50000 718
rect 47945 98 48011 101
rect 49200 98 50000 188
rect 47945 96 50000 98
rect 47945 40 47950 96
rect 48006 40 50000 96
rect 47945 38 50000 40
rect 47945 35 48011 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 46060 46956 46124 47020
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 46060 19756 46124 19820
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 46059 47020 46125 47021
rect 46059 46956 46060 47020
rect 46124 46956 46125 47020
rect 46059 46955 46125 46956
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 46062 19821 46122 46955
rect 46059 19820 46125 19821
rect 46059 19756 46060 19820
rect 46124 19756 46125 19820
rect 46059 19755 46125 19756
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 40664 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 19780 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform -1 0 25484 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 24196 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 20608 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1644511149
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_185
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_242
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1644511149
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_291
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_314
timestamp 1644511149
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1644511149
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1644511149
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1644511149
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_412
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_459
timestamp 1644511149
transform 1 0 43332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_467
timestamp 1644511149
transform 1 0 44068 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1644511149
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_95
timestamp 1644511149
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_102
timestamp 1644511149
transform 1 0 10488 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1644511149
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_133
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_156
timestamp 1644511149
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1644511149
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1644511149
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1644511149
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1644511149
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1644511149
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1644511149
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1644511149
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_254
timestamp 1644511149
transform 1 0 24472 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_271
timestamp 1644511149
transform 1 0 26036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_289
timestamp 1644511149
transform 1 0 27692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_301
timestamp 1644511149
transform 1 0 28796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_313
timestamp 1644511149
transform 1 0 29900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_325
timestamp 1644511149
transform 1 0 31004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1644511149
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_345
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_379
timestamp 1644511149
transform 1 0 35972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1644511149
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_414
timestamp 1644511149
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_439
timestamp 1644511149
transform 1 0 41492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_473
timestamp 1644511149
transform 1 0 44620 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_59
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_63
timestamp 1644511149
transform 1 0 6900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_74
timestamp 1644511149
transform 1 0 7912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1644511149
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_95
timestamp 1644511149
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_99
timestamp 1644511149
transform 1 0 10212 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_152
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1644511149
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_182
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1644511149
transform 1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_226
timestamp 1644511149
transform 1 0 21896 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_232
timestamp 1644511149
transform 1 0 22448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_236
timestamp 1644511149
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_243
timestamp 1644511149
transform 1 0 23460 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_260
timestamp 1644511149
transform 1 0 25024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_285
timestamp 1644511149
transform 1 0 27324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_297
timestamp 1644511149
transform 1 0 28428 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1644511149
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_330
timestamp 1644511149
transform 1 0 31464 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1644511149
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_346
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_350
timestamp 1644511149
transform 1 0 33304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_399
timestamp 1644511149
transform 1 0 37812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_411
timestamp 1644511149
transform 1 0 38916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1644511149
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_460
timestamp 1644511149
transform 1 0 43424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_467
timestamp 1644511149
transform 1 0 44068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1644511149
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_99
timestamp 1644511149
transform 1 0 10212 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_180
timestamp 1644511149
transform 1 0 17664 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1644511149
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_191
timestamp 1644511149
transform 1 0 18676 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_195
timestamp 1644511149
transform 1 0 19044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_202
timestamp 1644511149
transform 1 0 19688 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_210
timestamp 1644511149
transform 1 0 20424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1644511149
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_239
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1644511149
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_250
timestamp 1644511149
transform 1 0 24104 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_259
timestamp 1644511149
transform 1 0 24932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_266
timestamp 1644511149
transform 1 0 25576 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1644511149
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_424
timestamp 1644511149
transform 1 0 40112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_431
timestamp 1644511149
transform 1 0 40756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_443
timestamp 1644511149
transform 1 0 41860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_453
timestamp 1644511149
transform 1 0 42780 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_457
timestamp 1644511149
transform 1 0 43148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_482
timestamp 1644511149
transform 1 0 45448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_499
timestamp 1644511149
transform 1 0 47012 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_104
timestamp 1644511149
transform 1 0 10672 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_116
timestamp 1644511149
transform 1 0 11776 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_128
timestamp 1644511149
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_202
timestamp 1644511149
transform 1 0 19688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_216
timestamp 1644511149
transform 1 0 20976 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1644511149
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1644511149
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1644511149
transform 1 0 22908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1644511149
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_261
timestamp 1644511149
transform 1 0 25116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_283
timestamp 1644511149
transform 1 0 27140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_295
timestamp 1644511149
transform 1 0 28244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_468
timestamp 1644511149
transform 1 0 44160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_488
timestamp 1644511149
transform 1 0 46000 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_495
timestamp 1644511149
transform 1 0 46644 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_196
timestamp 1644511149
transform 1 0 19136 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_207
timestamp 1644511149
transform 1 0 20148 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1644511149
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_228
timestamp 1644511149
transform 1 0 22080 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_235
timestamp 1644511149
transform 1 0 22724 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_244
timestamp 1644511149
transform 1 0 23552 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_256
timestamp 1644511149
transform 1 0 24656 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_268
timestamp 1644511149
transform 1 0 25760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1644511149
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_64
timestamp 1644511149
transform 1 0 6992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp 1644511149
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_232
timestamp 1644511149
transform 1 0 22448 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_244
timestamp 1644511149
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1644511149
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1644511149
transform 1 0 8648 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1644511149
transform 1 0 9752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1644511149
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1644511149
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_69
timestamp 1644511149
transform 1 0 7452 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_73
timestamp 1644511149
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1644511149
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_497
timestamp 1644511149
transform 1 0 46828 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1644511149
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1644511149
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_157
timestamp 1644511149
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_161
timestamp 1644511149
transform 1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_186
timestamp 1644511149
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1644511149
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_500
timestamp 1644511149
transform 1 0 47104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_508
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_486
timestamp 1644511149
transform 1 0 45816 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_490
timestamp 1644511149
transform 1 0 46184 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_228
timestamp 1644511149
transform 1 0 22080 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_240
timestamp 1644511149
transform 1 0 23184 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_252
timestamp 1644511149
transform 1 0 24288 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_264
timestamp 1644511149
transform 1 0 25392 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_479
timestamp 1644511149
transform 1 0 45172 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_483
timestamp 1644511149
transform 1 0 45540 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1644511149
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_172
timestamp 1644511149
transform 1 0 16928 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_184
timestamp 1644511149
transform 1 0 18032 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_487
timestamp 1644511149
transform 1 0 45908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_155
timestamp 1644511149
transform 1 0 15364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_477
timestamp 1644511149
transform 1 0 44988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_500
timestamp 1644511149
transform 1 0 47104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_174
timestamp 1644511149
transform 1 0 17112 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_186
timestamp 1644511149
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1644511149
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_487
timestamp 1644511149
transform 1 0 45908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_512
timestamp 1644511149
transform 1 0 48208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_173
timestamp 1644511149
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_194
timestamp 1644511149
transform 1 0 18952 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_206
timestamp 1644511149
transform 1 0 20056 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1644511149
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_241
timestamp 1644511149
transform 1 0 23276 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_245
timestamp 1644511149
transform 1 0 23644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1644511149
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1644511149
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_482
timestamp 1644511149
transform 1 0 45448 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_492
timestamp 1644511149
transform 1 0 46368 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_499
timestamp 1644511149
transform 1 0 47012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1644511149
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_149
timestamp 1644511149
transform 1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_173
timestamp 1644511149
transform 1 0 17020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_181
timestamp 1644511149
transform 1 0 17756 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_187
timestamp 1644511149
transform 1 0 18308 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1644511149
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_201
timestamp 1644511149
transform 1 0 19596 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_232
timestamp 1644511149
transform 1 0 22448 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1644511149
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_485
timestamp 1644511149
transform 1 0 45724 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_491
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_498
timestamp 1644511149
transform 1 0 46920 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_507
timestamp 1644511149
transform 1 0 47748 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_515
timestamp 1644511149
transform 1 0 48484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1644511149
transform 1 0 13340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1644511149
transform 1 0 15548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_173
timestamp 1644511149
transform 1 0 17020 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1644511149
transform 1 0 18032 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_209
timestamp 1644511149
transform 1 0 20332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1644511149
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_248
timestamp 1644511149
transform 1 0 23920 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_255
timestamp 1644511149
transform 1 0 24564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_267
timestamp 1644511149
transform 1 0 25668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_491
timestamp 1644511149
transform 1 0 46276 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_500
timestamp 1644511149
transform 1 0 47104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_508
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1644511149
transform 1 0 14352 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_156
timestamp 1644511149
transform 1 0 15456 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1644511149
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_176
timestamp 1644511149
transform 1 0 17296 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_201
timestamp 1644511149
transform 1 0 19596 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_207
timestamp 1644511149
transform 1 0 20148 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_229
timestamp 1644511149
transform 1 0 22172 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_256
timestamp 1644511149
transform 1 0 24656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1644511149
transform 1 0 25300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_275
timestamp 1644511149
transform 1 0 26404 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_287
timestamp 1644511149
transform 1 0 27508 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1644511149
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_486
timestamp 1644511149
transform 1 0 45816 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_503
timestamp 1644511149
transform 1 0 47380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_510
timestamp 1644511149
transform 1 0 48024 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_99
timestamp 1644511149
transform 1 0 10212 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_103
timestamp 1644511149
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_154
timestamp 1644511149
transform 1 0 15272 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_160
timestamp 1644511149
transform 1 0 15824 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_192
timestamp 1644511149
transform 1 0 18768 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_204
timestamp 1644511149
transform 1 0 19872 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_213
timestamp 1644511149
transform 1 0 20700 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1644511149
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_239
timestamp 1644511149
transform 1 0 23092 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_250
timestamp 1644511149
transform 1 0 24104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_259
timestamp 1644511149
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_271
timestamp 1644511149
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_500
timestamp 1644511149
transform 1 0 47104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_510
timestamp 1644511149
transform 1 0 48024 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_114
timestamp 1644511149
transform 1 0 11592 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_126
timestamp 1644511149
transform 1 0 12696 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1644511149
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_145
timestamp 1644511149
transform 1 0 14444 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_152
timestamp 1644511149
transform 1 0 15088 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_160
timestamp 1644511149
transform 1 0 15824 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_182
timestamp 1644511149
transform 1 0 17848 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1644511149
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_237
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_244
timestamp 1644511149
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_258
timestamp 1644511149
transform 1 0 24840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_270
timestamp 1644511149
transform 1 0 25944 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_282
timestamp 1644511149
transform 1 0 27048 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_294
timestamp 1644511149
transform 1 0 28152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1644511149
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_504
timestamp 1644511149
transform 1 0 47472 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_511
timestamp 1644511149
transform 1 0 48116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_515
timestamp 1644511149
transform 1 0 48484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_177
timestamp 1644511149
transform 1 0 17388 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_185
timestamp 1644511149
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_190
timestamp 1644511149
transform 1 0 18584 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_199
timestamp 1644511149
transform 1 0 19412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_211
timestamp 1644511149
transform 1 0 20516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_265
timestamp 1644511149
transform 1 0 25484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1644511149
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_313
timestamp 1644511149
transform 1 0 29900 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_318
timestamp 1644511149
transform 1 0 30360 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_330
timestamp 1644511149
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_500
timestamp 1644511149
transform 1 0 47104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_103
timestamp 1644511149
transform 1 0 10580 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_125
timestamp 1644511149
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1644511149
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_145
timestamp 1644511149
transform 1 0 14444 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_157
timestamp 1644511149
transform 1 0 15548 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_179
timestamp 1644511149
transform 1 0 17572 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1644511149
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_207
timestamp 1644511149
transform 1 0 20148 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_228
timestamp 1644511149
transform 1 0 22080 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_240
timestamp 1644511149
transform 1 0 23184 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1644511149
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1644511149
transform 1 0 25300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_275
timestamp 1644511149
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_287
timestamp 1644511149
transform 1 0 27508 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_299
timestamp 1644511149
transform 1 0 28612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_313
timestamp 1644511149
transform 1 0 29900 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_335
timestamp 1644511149
transform 1 0 31924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_347
timestamp 1644511149
transform 1 0 33028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1644511149
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_434
timestamp 1644511149
transform 1 0 41032 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_446
timestamp 1644511149
transform 1 0 42136 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_458
timestamp 1644511149
transform 1 0 43240 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_470
timestamp 1644511149
transform 1 0 44344 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_156
timestamp 1644511149
transform 1 0 15456 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1644511149
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_173
timestamp 1644511149
transform 1 0 17020 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_206
timestamp 1644511149
transform 1 0 20056 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1644511149
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_248
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_257
timestamp 1644511149
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_265
timestamp 1644511149
transform 1 0 25484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_272
timestamp 1644511149
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_300
timestamp 1644511149
transform 1 0 28704 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_325
timestamp 1644511149
transform 1 0 31004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1644511149
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_126
timestamp 1644511149
transform 1 0 12696 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_135
timestamp 1644511149
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_146
timestamp 1644511149
transform 1 0 14536 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_158
timestamp 1644511149
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_166
timestamp 1644511149
transform 1 0 16376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_185
timestamp 1644511149
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1644511149
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_200
timestamp 1644511149
transform 1 0 19504 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_212
timestamp 1644511149
transform 1 0 20608 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_238
timestamp 1644511149
transform 1 0 23000 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1644511149
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_261
timestamp 1644511149
transform 1 0 25116 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_282
timestamp 1644511149
transform 1 0 27048 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_290
timestamp 1644511149
transform 1 0 27784 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_295
timestamp 1644511149
transform 1 0 28244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_322
timestamp 1644511149
transform 1 0 30728 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_334
timestamp 1644511149
transform 1 0 31832 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_346
timestamp 1644511149
transform 1 0 32936 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1644511149
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_483
timestamp 1644511149
transform 1 0 45540 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_487
timestamp 1644511149
transform 1 0 45908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_11
timestamp 1644511149
transform 1 0 2116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_23
timestamp 1644511149
transform 1 0 3220 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_35
timestamp 1644511149
transform 1 0 4324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1644511149
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_89
timestamp 1644511149
transform 1 0 9292 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_94
timestamp 1644511149
transform 1 0 9752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_101
timestamp 1644511149
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1644511149
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_116
timestamp 1644511149
transform 1 0 11776 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_128
timestamp 1644511149
transform 1 0 12880 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_146
timestamp 1644511149
transform 1 0 14536 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1644511149
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_176
timestamp 1644511149
transform 1 0 17296 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 1644511149
transform 1 0 18032 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_190
timestamp 1644511149
transform 1 0 18584 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_198
timestamp 1644511149
transform 1 0 19320 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_207
timestamp 1644511149
transform 1 0 20148 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 1644511149
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_229
timestamp 1644511149
transform 1 0 22172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_236
timestamp 1644511149
transform 1 0 22816 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_243
timestamp 1644511149
transform 1 0 23460 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_270
timestamp 1644511149
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1644511149
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_301
timestamp 1644511149
transform 1 0 28796 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_313
timestamp 1644511149
transform 1 0 29900 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_325
timestamp 1644511149
transform 1 0 31004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1644511149
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_489
timestamp 1644511149
transform 1 0 46092 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_493
timestamp 1644511149
transform 1 0 46460 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1644511149
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_107
timestamp 1644511149
transform 1 0 10948 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp 1644511149
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_161
timestamp 1644511149
transform 1 0 15916 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_170
timestamp 1644511149
transform 1 0 16744 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1644511149
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1644511149
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_203
timestamp 1644511149
transform 1 0 19780 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_232
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_239
timestamp 1644511149
transform 1 0 23092 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_257
timestamp 1644511149
transform 1 0 24748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_269
timestamp 1644511149
transform 1 0 25852 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_276
timestamp 1644511149
transform 1 0 26496 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_284
timestamp 1644511149
transform 1 0 27232 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_290
timestamp 1644511149
transform 1 0 27784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_297
timestamp 1644511149
transform 1 0 28428 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_305
timestamp 1644511149
transform 1 0 29164 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_485
timestamp 1644511149
transform 1 0 45724 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_508
timestamp 1644511149
transform 1 0 47840 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_91
timestamp 1644511149
transform 1 0 9476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 1644511149
transform 1 0 10212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1644511149
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1644511149
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1644511149
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_130
timestamp 1644511149
transform 1 0 13064 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_141
timestamp 1644511149
transform 1 0 14076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_153
timestamp 1644511149
transform 1 0 15180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1644511149
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_177
timestamp 1644511149
transform 1 0 17388 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_199
timestamp 1644511149
transform 1 0 19412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1644511149
transform 1 0 20148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_212
timestamp 1644511149
transform 1 0 20608 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_232
timestamp 1644511149
transform 1 0 22448 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1644511149
transform 1 0 24748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1644511149
transform 1 0 25852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1644511149
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_285
timestamp 1644511149
transform 1 0 27324 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_290
timestamp 1644511149
transform 1 0 27784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_302
timestamp 1644511149
transform 1 0 28888 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_314
timestamp 1644511149
transform 1 0 29992 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1644511149
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1644511149
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_494
timestamp 1644511149
transform 1 0 46552 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_502
timestamp 1644511149
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_99
timestamp 1644511149
transform 1 0 10212 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_111
timestamp 1644511149
transform 1 0 11316 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_116
timestamp 1644511149
transform 1 0 11776 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_128
timestamp 1644511149
transform 1 0 12880 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_148
timestamp 1644511149
transform 1 0 14720 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_156
timestamp 1644511149
transform 1 0 15456 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1644511149
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1644511149
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1644511149
transform 1 0 20056 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_214
timestamp 1644511149
transform 1 0 20792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1644511149
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_273
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_288
timestamp 1644511149
transform 1 0 27600 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_296
timestamp 1644511149
transform 1 0 28336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_487
timestamp 1644511149
transform 1 0 45908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1644511149
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_101
timestamp 1644511149
transform 1 0 10396 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1644511149
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1644511149
transform 1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1644511149
transform 1 0 14628 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_159
timestamp 1644511149
transform 1 0 15732 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_178
timestamp 1644511149
transform 1 0 17480 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_186
timestamp 1644511149
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_247
timestamp 1644511149
transform 1 0 23828 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1644511149
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_284
timestamp 1644511149
transform 1 0 27232 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_311
timestamp 1644511149
transform 1 0 29716 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_322
timestamp 1644511149
transform 1 0 30728 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1644511149
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_477
timestamp 1644511149
transform 1 0 44988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_481
timestamp 1644511149
transform 1 0 45356 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_488
timestamp 1644511149
transform 1 0 46000 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_499
timestamp 1644511149
transform 1 0 47012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_93
timestamp 1644511149
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1644511149
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_108
timestamp 1644511149
transform 1 0 11040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_116
timestamp 1644511149
transform 1 0 11776 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_128
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_144
timestamp 1644511149
transform 1 0 14352 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_201
timestamp 1644511149
transform 1 0 19596 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_213
timestamp 1644511149
transform 1 0 20700 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_231
timestamp 1644511149
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_239
timestamp 1644511149
transform 1 0 23092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1644511149
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_274
timestamp 1644511149
transform 1 0 26312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_281
timestamp 1644511149
transform 1 0 26956 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_292
timestamp 1644511149
transform 1 0 27968 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_317
timestamp 1644511149
transform 1 0 30268 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_339
timestamp 1644511149
transform 1 0 32292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_351
timestamp 1644511149
transform 1 0 33396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_65
timestamp 1644511149
transform 1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_88
timestamp 1644511149
transform 1 0 9200 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_100
timestamp 1644511149
transform 1 0 10304 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_179
timestamp 1644511149
transform 1 0 17572 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_187
timestamp 1644511149
transform 1 0 18308 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1644511149
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_215
timestamp 1644511149
transform 1 0 20884 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_245
timestamp 1644511149
transform 1 0 23644 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_251
timestamp 1644511149
transform 1 0 24196 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_264
timestamp 1644511149
transform 1 0 25392 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_289
timestamp 1644511149
transform 1 0 27692 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_300
timestamp 1644511149
transform 1 0 28704 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_312
timestamp 1644511149
transform 1 0 29808 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_324
timestamp 1644511149
transform 1 0 30912 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1644511149
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_69
timestamp 1644511149
transform 1 0 7452 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_73
timestamp 1644511149
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1644511149
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_105
timestamp 1644511149
transform 1 0 10764 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_112
timestamp 1644511149
transform 1 0 11408 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_120
timestamp 1644511149
transform 1 0 12144 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_128
timestamp 1644511149
transform 1 0 12880 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_135
timestamp 1644511149
transform 1 0 13524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_145
timestamp 1644511149
transform 1 0 14444 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_162
timestamp 1644511149
transform 1 0 16008 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_174
timestamp 1644511149
transform 1 0 17112 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_181
timestamp 1644511149
transform 1 0 17756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1644511149
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1644511149
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_206
timestamp 1644511149
transform 1 0 20056 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_216
timestamp 1644511149
transform 1 0 20976 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_240
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_261
timestamp 1644511149
transform 1 0 25116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_273
timestamp 1644511149
transform 1 0 26220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_280
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_66
timestamp 1644511149
transform 1 0 7176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_91
timestamp 1644511149
transform 1 0 9476 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_98
timestamp 1644511149
transform 1 0 10120 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1644511149
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_134
timestamp 1644511149
transform 1 0 13432 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1644511149
transform 1 0 14168 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_210
timestamp 1644511149
transform 1 0 20424 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_214
timestamp 1644511149
transform 1 0 20792 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_234
timestamp 1644511149
transform 1 0 22632 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_242
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_268
timestamp 1644511149
transform 1 0 25760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_287
timestamp 1644511149
transform 1 0 27508 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_299
timestamp 1644511149
transform 1 0 28612 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_307
timestamp 1644511149
transform 1 0 29348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_312
timestamp 1644511149
transform 1 0 29808 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_324
timestamp 1644511149
transform 1 0 30912 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_489
timestamp 1644511149
transform 1 0 46092 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_508
timestamp 1644511149
transform 1 0 47840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_74
timestamp 1644511149
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1644511149
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_88
timestamp 1644511149
transform 1 0 9200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_92
timestamp 1644511149
transform 1 0 9568 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_96
timestamp 1644511149
transform 1 0 9936 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_120
timestamp 1644511149
transform 1 0 12144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_127
timestamp 1644511149
transform 1 0 12788 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_149
timestamp 1644511149
transform 1 0 14812 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_155
timestamp 1644511149
transform 1 0 15364 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_163
timestamp 1644511149
transform 1 0 16100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_173
timestamp 1644511149
transform 1 0 17020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_181
timestamp 1644511149
transform 1 0 17756 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_206
timestamp 1644511149
transform 1 0 20056 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_210
timestamp 1644511149
transform 1 0 20424 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_223
timestamp 1644511149
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_276
timestamp 1644511149
transform 1 0 26496 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_287
timestamp 1644511149
transform 1 0 27508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_296
timestamp 1644511149
transform 1 0 28336 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_300
timestamp 1644511149
transform 1 0 28704 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_319
timestamp 1644511149
transform 1 0 30452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_331
timestamp 1644511149
transform 1 0 31556 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_343
timestamp 1644511149
transform 1 0 32660 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_355
timestamp 1644511149
transform 1 0 33764 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_90
timestamp 1644511149
transform 1 0 9384 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_102
timestamp 1644511149
transform 1 0 10488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1644511149
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_123
timestamp 1644511149
transform 1 0 12420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_148
timestamp 1644511149
transform 1 0 14720 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_156
timestamp 1644511149
transform 1 0 15456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_189
timestamp 1644511149
transform 1 0 18492 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_195
timestamp 1644511149
transform 1 0 19044 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_233
timestamp 1644511149
transform 1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_241
timestamp 1644511149
transform 1 0 23276 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_248
timestamp 1644511149
transform 1 0 23920 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_258
timestamp 1644511149
transform 1 0 24840 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_264
timestamp 1644511149
transform 1 0 25392 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_268
timestamp 1644511149
transform 1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_301
timestamp 1644511149
transform 1 0 28796 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_309
timestamp 1644511149
transform 1 0 29532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_432
timestamp 1644511149
transform 1 0 40848 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_440
timestamp 1644511149
transform 1 0 41584 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_455
timestamp 1644511149
transform 1 0 42964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_467
timestamp 1644511149
transform 1 0 44068 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_479
timestamp 1644511149
transform 1 0 45172 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_491
timestamp 1644511149
transform 1 0 46276 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_104
timestamp 1644511149
transform 1 0 10672 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_116
timestamp 1644511149
transform 1 0 11776 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_122
timestamp 1644511149
transform 1 0 12328 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_145
timestamp 1644511149
transform 1 0 14444 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_155
timestamp 1644511149
transform 1 0 15364 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_161
timestamp 1644511149
transform 1 0 15916 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_168
timestamp 1644511149
transform 1 0 16560 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_176
timestamp 1644511149
transform 1 0 17296 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_182
timestamp 1644511149
transform 1 0 17848 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_186
timestamp 1644511149
transform 1 0 18216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1644511149
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_257
timestamp 1644511149
transform 1 0 24748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_269
timestamp 1644511149
transform 1 0 25852 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_275
timestamp 1644511149
transform 1 0 26404 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_280
timestamp 1644511149
transform 1 0 26864 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_287
timestamp 1644511149
transform 1 0 27508 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_299
timestamp 1644511149
transform 1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_330
timestamp 1644511149
transform 1 0 31464 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_342
timestamp 1644511149
transform 1 0 32568 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_354
timestamp 1644511149
transform 1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1644511149
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_483
timestamp 1644511149
transform 1 0 45540 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_487
timestamp 1644511149
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_100
timestamp 1644511149
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_129
timestamp 1644511149
transform 1 0 12972 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_150
timestamp 1644511149
transform 1 0 14904 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1644511149
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_177
timestamp 1644511149
transform 1 0 17388 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_183
timestamp 1644511149
transform 1 0 17940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_195
timestamp 1644511149
transform 1 0 19044 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_200
timestamp 1644511149
transform 1 0 19504 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_204
timestamp 1644511149
transform 1 0 19872 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1644511149
transform 1 0 20240 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_233
timestamp 1644511149
transform 1 0 22540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_241
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_263
timestamp 1644511149
transform 1 0 25300 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_275
timestamp 1644511149
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_9
timestamp 1644511149
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1644511149
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_89
timestamp 1644511149
transform 1 0 9292 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_113
timestamp 1644511149
transform 1 0 11500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_125
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_131
timestamp 1644511149
transform 1 0 13156 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_144
timestamp 1644511149
transform 1 0 14352 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_156
timestamp 1644511149
transform 1 0 15456 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_162
timestamp 1644511149
transform 1 0 16008 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_170
timestamp 1644511149
transform 1 0 16744 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_182
timestamp 1644511149
transform 1 0 17848 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1644511149
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_217
timestamp 1644511149
transform 1 0 21068 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 1644511149
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_238
timestamp 1644511149
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1644511149
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_259
timestamp 1644511149
transform 1 0 24932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_283
timestamp 1644511149
transform 1 0 27140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_295
timestamp 1644511149
transform 1 0 28244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_487
timestamp 1644511149
transform 1 0 45908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_118
timestamp 1644511149
transform 1 0 11960 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_126
timestamp 1644511149
transform 1 0 12696 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_133
timestamp 1644511149
transform 1 0 13340 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_140
timestamp 1644511149
transform 1 0 13984 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_152
timestamp 1644511149
transform 1 0 15088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_156
timestamp 1644511149
transform 1 0 15456 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_189
timestamp 1644511149
transform 1 0 18492 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_197
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_204
timestamp 1644511149
transform 1 0 19872 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_211
timestamp 1644511149
transform 1 0 20516 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_234
timestamp 1644511149
transform 1 0 22632 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_246
timestamp 1644511149
transform 1 0 23736 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_257
timestamp 1644511149
transform 1 0 24748 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_268
timestamp 1644511149
transform 1 0 25760 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_476
timestamp 1644511149
transform 1 0 44896 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_500
timestamp 1644511149
transform 1 0 47104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_511
timestamp 1644511149
transform 1 0 48116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_515
timestamp 1644511149
transform 1 0 48484 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_101
timestamp 1644511149
transform 1 0 10396 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_122
timestamp 1644511149
transform 1 0 12328 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_128
timestamp 1644511149
transform 1 0 12880 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_144
timestamp 1644511149
transform 1 0 14352 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_160
timestamp 1644511149
transform 1 0 15824 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_168
timestamp 1644511149
transform 1 0 16560 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_175
timestamp 1644511149
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1644511149
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_217
timestamp 1644511149
transform 1 0 21068 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_227
timestamp 1644511149
transform 1 0 21988 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_235
timestamp 1644511149
transform 1 0 22724 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_243
timestamp 1644511149
transform 1 0 23460 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_247
timestamp 1644511149
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_269
timestamp 1644511149
transform 1 0 25852 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_274
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_286
timestamp 1644511149
transform 1 0 27416 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_298
timestamp 1644511149
transform 1 0 28520 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1644511149
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_486
timestamp 1644511149
transform 1 0 45816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_511
timestamp 1644511149
transform 1 0 48116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_515
timestamp 1644511149
transform 1 0 48484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_99
timestamp 1644511149
transform 1 0 10212 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1644511149
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_121
timestamp 1644511149
transform 1 0 12236 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_127
timestamp 1644511149
transform 1 0 12788 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_148
timestamp 1644511149
transform 1 0 14720 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_156
timestamp 1644511149
transform 1 0 15456 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_191
timestamp 1644511149
transform 1 0 18676 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_203
timestamp 1644511149
transform 1 0 19780 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_214
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1644511149
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_233
timestamp 1644511149
transform 1 0 22540 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_245
timestamp 1644511149
transform 1 0 23644 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_257
timestamp 1644511149
transform 1 0 24748 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_265
timestamp 1644511149
transform 1 0 25484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_289
timestamp 1644511149
transform 1 0 27692 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_294
timestamp 1644511149
transform 1 0 28152 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_302
timestamp 1644511149
transform 1 0 28888 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_324
timestamp 1644511149
transform 1 0 30912 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_112
timestamp 1644511149
transform 1 0 11408 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_144
timestamp 1644511149
transform 1 0 14352 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_151
timestamp 1644511149
transform 1 0 14996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_163
timestamp 1644511149
transform 1 0 16100 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_175
timestamp 1644511149
transform 1 0 17204 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_180
timestamp 1644511149
transform 1 0 17664 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 1644511149
transform 1 0 18676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_217
timestamp 1644511149
transform 1 0 21068 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_225
timestamp 1644511149
transform 1 0 21804 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_262
timestamp 1644511149
transform 1 0 25208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_273
timestamp 1644511149
transform 1 0 26220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_282
timestamp 1644511149
transform 1 0 27048 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_290
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_294
timestamp 1644511149
transform 1 0 28152 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_315
timestamp 1644511149
transform 1 0 30084 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_319
timestamp 1644511149
transform 1 0 30452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_331
timestamp 1644511149
transform 1 0 31556 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_343
timestamp 1644511149
transform 1 0 32660 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_355
timestamp 1644511149
transform 1 0 33764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1644511149
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_116
timestamp 1644511149
transform 1 0 11776 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_122
timestamp 1644511149
transform 1 0 12328 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_126
timestamp 1644511149
transform 1 0 12696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_138
timestamp 1644511149
transform 1 0 13800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_142
timestamp 1644511149
transform 1 0 14168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_177
timestamp 1644511149
transform 1 0 17388 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_198
timestamp 1644511149
transform 1 0 19320 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_207
timestamp 1644511149
transform 1 0 20148 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_216
timestamp 1644511149
transform 1 0 20976 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_229
timestamp 1644511149
transform 1 0 22172 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_241
timestamp 1644511149
transform 1 0 23276 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_259
timestamp 1644511149
transform 1 0 24932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_263
timestamp 1644511149
transform 1 0 25300 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1644511149
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_301
timestamp 1644511149
transform 1 0 28796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_310
timestamp 1644511149
transform 1 0 29624 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_322
timestamp 1644511149
transform 1 0 30728 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_326
timestamp 1644511149
transform 1 0 31096 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1644511149
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_500
timestamp 1644511149
transform 1 0 47104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_106
timestamp 1644511149
transform 1 0 10856 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_131
timestamp 1644511149
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_162
timestamp 1644511149
transform 1 0 16008 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_186
timestamp 1644511149
transform 1 0 18216 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1644511149
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_204
timestamp 1644511149
transform 1 0 19872 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_212
timestamp 1644511149
transform 1 0 20608 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_235
timestamp 1644511149
transform 1 0 22724 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1644511149
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_260
timestamp 1644511149
transform 1 0 25024 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_270
timestamp 1644511149
transform 1 0 25944 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_274
timestamp 1644511149
transform 1 0 26312 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_284
timestamp 1644511149
transform 1 0 27232 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_292
timestamp 1644511149
transform 1 0 27968 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_299
timestamp 1644511149
transform 1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_512
timestamp 1644511149
transform 1 0 48208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_136
timestamp 1644511149
transform 1 0 13616 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_140
timestamp 1644511149
transform 1 0 13984 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1644511149
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_180
timestamp 1644511149
transform 1 0 17664 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_203
timestamp 1644511149
transform 1 0 19780 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1644511149
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_230
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_242
timestamp 1644511149
transform 1 0 23368 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_254
timestamp 1644511149
transform 1 0 24472 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_262
timestamp 1644511149
transform 1 0 25208 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_270
timestamp 1644511149
transform 1 0 25944 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1644511149
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_300
timestamp 1644511149
transform 1 0 28704 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_313
timestamp 1644511149
transform 1 0 29900 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_320
timestamp 1644511149
transform 1 0 30544 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_145
timestamp 1644511149
transform 1 0 14444 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_152
timestamp 1644511149
transform 1 0 15088 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_164
timestamp 1644511149
transform 1 0 16192 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_172
timestamp 1644511149
transform 1 0 16928 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_180
timestamp 1644511149
transform 1 0 17664 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1644511149
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_218
timestamp 1644511149
transform 1 0 21160 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_228
timestamp 1644511149
transform 1 0 22080 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_235
timestamp 1644511149
transform 1 0 22724 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1644511149
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_257
timestamp 1644511149
transform 1 0 24748 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_267
timestamp 1644511149
transform 1 0 25668 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_276
timestamp 1644511149
transform 1 0 26496 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_284
timestamp 1644511149
transform 1 0 27232 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_291
timestamp 1644511149
transform 1 0 27876 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_300
timestamp 1644511149
transform 1 0 28704 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_328
timestamp 1644511149
transform 1 0 31280 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_340
timestamp 1644511149
transform 1 0 32384 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_352
timestamp 1644511149
transform 1 0 33488 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_150
timestamp 1644511149
transform 1 0 14904 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_162
timestamp 1644511149
transform 1 0 16008 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1644511149
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1644511149
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_230
timestamp 1644511149
transform 1 0 22264 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_242
timestamp 1644511149
transform 1 0 23368 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_260
timestamp 1644511149
transform 1 0 25024 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1644511149
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_285
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_294
timestamp 1644511149
transform 1 0 28152 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_307
timestamp 1644511149
transform 1 0 29348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_311
timestamp 1644511149
transform 1 0 29716 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_319
timestamp 1644511149
transform 1 0 30452 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_159
timestamp 1644511149
transform 1 0 15732 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_178
timestamp 1644511149
transform 1 0 17480 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_188
timestamp 1644511149
transform 1 0 18400 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_213
timestamp 1644511149
transform 1 0 20700 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_220
timestamp 1644511149
transform 1 0 21344 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_228
timestamp 1644511149
transform 1 0 22080 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_237
timestamp 1644511149
transform 1 0 22908 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_243
timestamp 1644511149
transform 1 0 23460 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_269
timestamp 1644511149
transform 1 0 25852 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_295
timestamp 1644511149
transform 1 0 28244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_315
timestamp 1644511149
transform 1 0 30084 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_336
timestamp 1644511149
transform 1 0 32016 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_348
timestamp 1644511149
transform 1 0 33120 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1644511149
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_14
timestamp 1644511149
transform 1 0 2392 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_26
timestamp 1644511149
transform 1 0 3496 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_38
timestamp 1644511149
transform 1 0 4600 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_50
timestamp 1644511149
transform 1 0 5704 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_143
timestamp 1644511149
transform 1 0 14260 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1644511149
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_176
timestamp 1644511149
transform 1 0 17296 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_180
timestamp 1644511149
transform 1 0 17664 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_188
timestamp 1644511149
transform 1 0 18400 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_200
timestamp 1644511149
transform 1 0 19504 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_245
timestamp 1644511149
transform 1 0 23644 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_269
timestamp 1644511149
transform 1 0 25852 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_277
timestamp 1644511149
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_289
timestamp 1644511149
transform 1 0 27692 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_297
timestamp 1644511149
transform 1 0 28428 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_320
timestamp 1644511149
transform 1 0 30544 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_163
timestamp 1644511149
transform 1 0 16100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_173
timestamp 1644511149
transform 1 0 17020 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_185
timestamp 1644511149
transform 1 0 18124 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_231
timestamp 1644511149
transform 1 0 22356 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_246
timestamp 1644511149
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_260
timestamp 1644511149
transform 1 0 25024 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_264
timestamp 1644511149
transform 1 0 25392 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_269
timestamp 1644511149
transform 1 0 25852 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_287
timestamp 1644511149
transform 1 0 27508 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_298
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1644511149
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_315
timestamp 1644511149
transform 1 0 30084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_327
timestamp 1644511149
transform 1 0 31188 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_339
timestamp 1644511149
transform 1 0 32292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_351
timestamp 1644511149
transform 1 0 33396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_9
timestamp 1644511149
transform 1 0 1932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_34
timestamp 1644511149
transform 1 0 4232 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_46
timestamp 1644511149
transform 1 0 5336 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1644511149
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_158
timestamp 1644511149
transform 1 0 15640 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1644511149
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_173
timestamp 1644511149
transform 1 0 17020 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_177
timestamp 1644511149
transform 1 0 17388 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1644511149
transform 1 0 18032 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1644511149
transform 1 0 19136 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_216
timestamp 1644511149
transform 1 0 20976 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_229
timestamp 1644511149
transform 1 0 22172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_236
timestamp 1644511149
transform 1 0 22816 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_245
timestamp 1644511149
transform 1 0 23644 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_254
timestamp 1644511149
transform 1 0 24472 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_258
timestamp 1644511149
transform 1 0 24840 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_263
timestamp 1644511149
transform 1 0 25300 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_269
timestamp 1644511149
transform 1 0 25852 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_289
timestamp 1644511149
transform 1 0 27692 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_296
timestamp 1644511149
transform 1 0 28336 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_308
timestamp 1644511149
transform 1 0 29440 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_312
timestamp 1644511149
transform 1 0 29808 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_321
timestamp 1644511149
transform 1 0 30636 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_327
timestamp 1644511149
transform 1 0 31188 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_331
timestamp 1644511149
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_508
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1644511149
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_173
timestamp 1644511149
transform 1 0 17020 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_181
timestamp 1644511149
transform 1 0 17756 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_186
timestamp 1644511149
transform 1 0 18216 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1644511149
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_205
timestamp 1644511149
transform 1 0 19964 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_216
timestamp 1644511149
transform 1 0 20976 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_228
timestamp 1644511149
transform 1 0 22080 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_237
timestamp 1644511149
transform 1 0 22908 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_285
timestamp 1644511149
transform 1 0 27324 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_293
timestamp 1644511149
transform 1 0 28060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1644511149
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_312
timestamp 1644511149
transform 1 0 29808 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_340
timestamp 1644511149
transform 1 0 32384 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_352
timestamp 1644511149
transform 1 0 33488 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_157
timestamp 1644511149
transform 1 0 15548 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_175
timestamp 1644511149
transform 1 0 17204 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_182
timestamp 1644511149
transform 1 0 17848 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_195
timestamp 1644511149
transform 1 0 19044 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_201
timestamp 1644511149
transform 1 0 19596 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_206
timestamp 1644511149
transform 1 0 20056 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_232
timestamp 1644511149
transform 1 0 22448 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_244
timestamp 1644511149
transform 1 0 23552 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_254
timestamp 1644511149
transform 1 0 24472 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_263
timestamp 1644511149
transform 1 0 25300 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_271
timestamp 1644511149
transform 1 0 26036 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_285
timestamp 1644511149
transform 1 0 27324 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_301
timestamp 1644511149
transform 1 0 28796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_310
timestamp 1644511149
transform 1 0 29624 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_512
timestamp 1644511149
transform 1 0 48208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_162
timestamp 1644511149
transform 1 0 16008 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_169
timestamp 1644511149
transform 1 0 16652 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_173
timestamp 1644511149
transform 1 0 17020 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_180
timestamp 1644511149
transform 1 0 17664 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_190
timestamp 1644511149
transform 1 0 18584 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_201
timestamp 1644511149
transform 1 0 19596 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_213
timestamp 1644511149
transform 1 0 20700 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_228
timestamp 1644511149
transform 1 0 22080 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_236
timestamp 1644511149
transform 1 0 22816 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_261
timestamp 1644511149
transform 1 0 25116 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_273
timestamp 1644511149
transform 1 0 26220 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_279
timestamp 1644511149
transform 1 0 26772 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_283
timestamp 1644511149
transform 1 0 27140 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_294
timestamp 1644511149
transform 1 0 28152 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1644511149
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_324
timestamp 1644511149
transform 1 0 30912 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_336
timestamp 1644511149
transform 1 0 32016 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_348
timestamp 1644511149
transform 1 0 33120 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1644511149
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_497
timestamp 1644511149
transform 1 0 46828 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_184
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_194
timestamp 1644511149
transform 1 0 18952 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_203
timestamp 1644511149
transform 1 0 19780 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_215
timestamp 1644511149
transform 1 0 20884 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_245
timestamp 1644511149
transform 1 0 23644 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_259
timestamp 1644511149
transform 1 0 24932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_269
timestamp 1644511149
transform 1 0 25852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1644511149
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_287
timestamp 1644511149
transform 1 0 27508 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_297
timestamp 1644511149
transform 1 0 28428 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_307
timestamp 1644511149
transform 1 0 29348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_320
timestamp 1644511149
transform 1 0 30544 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_330
timestamp 1644511149
transform 1 0 31464 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_512
timestamp 1644511149
transform 1 0 48208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_162
timestamp 1644511149
transform 1 0 16008 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_174
timestamp 1644511149
transform 1 0 17112 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_178
timestamp 1644511149
transform 1 0 17480 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_185
timestamp 1644511149
transform 1 0 18124 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_193
timestamp 1644511149
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_204
timestamp 1644511149
transform 1 0 19872 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_210
timestamp 1644511149
transform 1 0 20424 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_218
timestamp 1644511149
transform 1 0 21160 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_226
timestamp 1644511149
transform 1 0 21896 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_230
timestamp 1644511149
transform 1 0 22264 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_234
timestamp 1644511149
transform 1 0 22632 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_246
timestamp 1644511149
transform 1 0 23736 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_276
timestamp 1644511149
transform 1 0 26496 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_286
timestamp 1644511149
transform 1 0 27416 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_297
timestamp 1644511149
transform 1 0 28428 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1644511149
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_315
timestamp 1644511149
transform 1 0 30084 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_336
timestamp 1644511149
transform 1 0 32016 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_348
timestamp 1644511149
transform 1 0 33120 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1644511149
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_153
timestamp 1644511149
transform 1 0 15180 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_157
timestamp 1644511149
transform 1 0 15548 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 1644511149
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_215
timestamp 1644511149
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_245
timestamp 1644511149
transform 1 0 23644 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_251
timestamp 1644511149
transform 1 0 24196 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_258
timestamp 1644511149
transform 1 0 24840 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_266
timestamp 1644511149
transform 1 0 25576 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_271
timestamp 1644511149
transform 1 0 26036 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_287
timestamp 1644511149
transform 1 0 27508 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_308
timestamp 1644511149
transform 1 0 29440 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_320
timestamp 1644511149
transform 1 0 30544 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_326
timestamp 1644511149
transform 1 0 31096 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_330
timestamp 1644511149
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1644511149
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1644511149
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_149
timestamp 1644511149
transform 1 0 14812 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_155
timestamp 1644511149
transform 1 0 15364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_168
timestamp 1644511149
transform 1 0 16560 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_181
timestamp 1644511149
transform 1 0 17756 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_187
timestamp 1644511149
transform 1 0 18308 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_200
timestamp 1644511149
transform 1 0 19504 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_210
timestamp 1644511149
transform 1 0 20424 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_222
timestamp 1644511149
transform 1 0 21528 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_234
timestamp 1644511149
transform 1 0 22632 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_238
timestamp 1644511149
transform 1 0 23000 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_258
timestamp 1644511149
transform 1 0 24840 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_272
timestamp 1644511149
transform 1 0 26128 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_284
timestamp 1644511149
transform 1 0 27232 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_288
timestamp 1644511149
transform 1 0 27600 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_298
timestamp 1644511149
transform 1 0 28520 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1644511149
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_312
timestamp 1644511149
transform 1 0 29808 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_324
timestamp 1644511149
transform 1 0 30912 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_336
timestamp 1644511149
transform 1 0 32016 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_348
timestamp 1644511149
transform 1 0 33120 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1644511149
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_28
timestamp 1644511149
transform 1 0 3680 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1644511149
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_143
timestamp 1644511149
transform 1 0 14260 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1644511149
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_190
timestamp 1644511149
transform 1 0 18584 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_202
timestamp 1644511149
transform 1 0 19688 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1644511149
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1644511149
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_229
timestamp 1644511149
transform 1 0 22172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_236
timestamp 1644511149
transform 1 0 22816 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_240
timestamp 1644511149
transform 1 0 23184 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_250
timestamp 1644511149
transform 1 0 24104 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_256
timestamp 1644511149
transform 1 0 24656 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_262
timestamp 1644511149
transform 1 0 25208 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 1644511149
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_284
timestamp 1644511149
transform 1 0 27232 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_290
timestamp 1644511149
transform 1 0 27784 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_311
timestamp 1644511149
transform 1 0 29716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_323
timestamp 1644511149
transform 1 0 30820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1644511149
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_215
timestamp 1644511149
transform 1 0 20884 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_239
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_285
timestamp 1644511149
transform 1 0 27324 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_297
timestamp 1644511149
transform 1 0 28428 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_512
timestamp 1644511149
transform 1 0 48208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_164
timestamp 1644511149
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_172
timestamp 1644511149
transform 1 0 16928 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_178
timestamp 1644511149
transform 1 0 17480 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_188
timestamp 1644511149
transform 1 0 18400 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_203
timestamp 1644511149
transform 1 0 19780 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_210
timestamp 1644511149
transform 1 0 20424 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_229
timestamp 1644511149
transform 1 0 22172 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_257
timestamp 1644511149
transform 1 0 24748 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_269
timestamp 1644511149
transform 1 0 25852 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_277
timestamp 1644511149
transform 1 0 26588 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_500
timestamp 1644511149
transform 1 0 47104 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_173
timestamp 1644511149
transform 1 0 17020 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_183
timestamp 1644511149
transform 1 0 17940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_217
timestamp 1644511149
transform 1 0 21068 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_229
timestamp 1644511149
transform 1 0 22172 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_237
timestamp 1644511149
transform 1 0 22908 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_243
timestamp 1644511149
transform 1 0 23460 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_260
timestamp 1644511149
transform 1 0 25024 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_272
timestamp 1644511149
transform 1 0 26128 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_284
timestamp 1644511149
transform 1 0 27232 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_296
timestamp 1644511149
transform 1 0 28336 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_197
timestamp 1644511149
transform 1 0 19228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_201
timestamp 1644511149
transform 1 0 19596 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_216
timestamp 1644511149
transform 1 0 20976 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_245
timestamp 1644511149
transform 1 0 23644 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_253
timestamp 1644511149
transform 1 0 24380 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_264
timestamp 1644511149
transform 1 0 25392 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_500
timestamp 1644511149
transform 1 0 47104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_469
timestamp 1644511149
transform 1 0 44252 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_483
timestamp 1644511149
transform 1 0 45540 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_495
timestamp 1644511149
transform 1 0 46644 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_499
timestamp 1644511149
transform 1 0 47012 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_505
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_512
timestamp 1644511149
transform 1 0 48208 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_13
timestamp 1644511149
transform 1 0 2300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_25
timestamp 1644511149
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_287
timestamp 1644511149
transform 1 0 27508 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_299
timestamp 1644511149
transform 1 0 28612 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_499
timestamp 1644511149
transform 1 0 47012 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_503
timestamp 1644511149
transform 1 0 47380 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_9
timestamp 1644511149
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_13
timestamp 1644511149
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_25
timestamp 1644511149
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_37
timestamp 1644511149
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1644511149
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_500
timestamp 1644511149
transform 1 0 47104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_508
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_271
timestamp 1644511149
transform 1 0 26036 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_296
timestamp 1644511149
transform 1 0 28336 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1644511149
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_13
timestamp 1644511149
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_25
timestamp 1644511149
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_37
timestamp 1644511149
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1644511149
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_489
timestamp 1644511149
transform 1 0 46092 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_493
timestamp 1644511149
transform 1 0 46460 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_248
timestamp 1644511149
transform 1 0 23920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_274
timestamp 1644511149
transform 1 0 26312 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_286
timestamp 1644511149
transform 1 0 27416 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_298
timestamp 1644511149
transform 1 0 28520 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1644511149
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_245
timestamp 1644511149
transform 1 0 23644 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_253
timestamp 1644511149
transform 1 0 24380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_275
timestamp 1644511149
transform 1 0 26404 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_455
timestamp 1644511149
transform 1 0 42964 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_463
timestamp 1644511149
transform 1 0 43700 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_468
timestamp 1644511149
transform 1 0 44160 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_476
timestamp 1644511149
transform 1 0 44896 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_482
timestamp 1644511149
transform 1 0 45448 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_220
timestamp 1644511149
transform 1 0 21344 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_232
timestamp 1644511149
transform 1 0 22448 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_244
timestamp 1644511149
transform 1 0 23552 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_260
timestamp 1644511149
transform 1 0 25024 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_272
timestamp 1644511149
transform 1 0 26128 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_284
timestamp 1644511149
transform 1 0 27232 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_296
timestamp 1644511149
transform 1 0 28336 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_449
timestamp 1644511149
transform 1 0 42412 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_453
timestamp 1644511149
transform 1 0 42780 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_460
timestamp 1644511149
transform 1 0 43424 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_468
timestamp 1644511149
transform 1 0 44160 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_477
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_485
timestamp 1644511149
transform 1 0 45724 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_14
timestamp 1644511149
transform 1 0 2392 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_26
timestamp 1644511149
transform 1 0 3496 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_38
timestamp 1644511149
transform 1 0 4600 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_50
timestamp 1644511149
transform 1 0 5704 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_101
timestamp 1644511149
transform 1 0 10396 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_107
timestamp 1644511149
transform 1 0 10948 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_213
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_218
timestamp 1644511149
transform 1 0 21160 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_340
timestamp 1644511149
transform 1 0 32384 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_352
timestamp 1644511149
transform 1 0 33488 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_364
timestamp 1644511149
transform 1 0 34592 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_376
timestamp 1644511149
transform 1 0 35696 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1644511149
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_433
timestamp 1644511149
transform 1 0 40940 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_437
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_444
timestamp 1644511149
transform 1 0 41952 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_472
timestamp 1644511149
transform 1 0 44528 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_482
timestamp 1644511149
transform 1 0 45448 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_489
timestamp 1644511149
transform 1 0 46092 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1644511149
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_508
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1644511149
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_36
timestamp 1644511149
transform 1 0 4416 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_40
timestamp 1644511149
transform 1 0 4784 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_44
timestamp 1644511149
transform 1 0 5152 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_56
timestamp 1644511149
transform 1 0 6256 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_68
timestamp 1644511149
transform 1 0 7360 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_80
timestamp 1644511149
transform 1 0 8464 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_124
timestamp 1644511149
transform 1 0 12512 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_128
timestamp 1644511149
transform 1 0 12880 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1644511149
transform 1 0 13524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_200
timestamp 1644511149
transform 1 0 19504 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_207
timestamp 1644511149
transform 1 0 20148 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_236
timestamp 1644511149
transform 1 0 22816 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_248
timestamp 1644511149
transform 1 0 23920 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_261
timestamp 1644511149
transform 1 0 25116 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_283
timestamp 1644511149
transform 1 0 27140 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_290
timestamp 1644511149
transform 1 0 27784 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_302
timestamp 1644511149
transform 1 0 28888 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_329
timestamp 1644511149
transform 1 0 31372 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_353
timestamp 1644511149
transform 1 0 33580 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_361
timestamp 1644511149
transform 1 0 34316 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_407
timestamp 1644511149
transform 1 0 38548 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1644511149
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_458
timestamp 1644511149
transform 1 0 43240 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_464
timestamp 1644511149
transform 1 0 43792 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_7
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_14
timestamp 1644511149
transform 1 0 2392 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_26
timestamp 1644511149
transform 1 0 3496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_30
timestamp 1644511149
transform 1 0 3864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1644511149
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_101
timestamp 1644511149
transform 1 0 10396 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_106
timestamp 1644511149
transform 1 0 10856 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_132
timestamp 1644511149
transform 1 0 13248 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_157
timestamp 1644511149
transform 1 0 15548 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_165
timestamp 1644511149
transform 1 0 16284 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_266
timestamp 1644511149
transform 1 0 25576 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1644511149
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_302
timestamp 1644511149
transform 1 0 28888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_327
timestamp 1644511149
transform 1 0 31188 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_340
timestamp 1644511149
transform 1 0 32384 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_352
timestamp 1644511149
transform 1 0 33488 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_364
timestamp 1644511149
transform 1 0 34592 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_376
timestamp 1644511149
transform 1 0 35696 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_388
timestamp 1644511149
transform 1 0 36800 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_431
timestamp 1644511149
transform 1 0 40756 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_437
timestamp 1644511149
transform 1 0 41308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1644511149
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_57
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_67
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_75
timestamp 1644511149
transform 1 0 8004 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_121
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_132
timestamp 1644511149
transform 1 0 13248 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_151
timestamp 1644511149
transform 1 0 14996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_163
timestamp 1644511149
transform 1 0 16100 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_191
timestamp 1644511149
transform 1 0 18676 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_201
timestamp 1644511149
transform 1 0 19596 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_216
timestamp 1644511149
transform 1 0 20976 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_300
timestamp 1644511149
transform 1 0 28704 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_332
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_406
timestamp 1644511149
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_418
timestamp 1644511149
transform 1 0 39560 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_441
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_447
timestamp 1644511149
transform 1 0 42228 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_511
timestamp 1644511149
transform 1 0 48116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_515
timestamp 1644511149
transform 1 0 48484 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0571_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0573_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0574_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0575_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27692 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0576_
timestamp 1644511149
transform 1 0 28888 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0577_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26036 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0578_
timestamp 1644511149
transform 1 0 18124 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0579_
timestamp 1644511149
transform 1 0 18400 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0580_
timestamp 1644511149
transform 1 0 18032 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0581_
timestamp 1644511149
transform 1 0 28796 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0582_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0583_
timestamp 1644511149
transform 1 0 24380 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0584_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23828 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0585_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0586_
timestamp 1644511149
transform 1 0 19688 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0587_
timestamp 1644511149
transform 1 0 20884 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0588_
timestamp 1644511149
transform 1 0 20516 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0589_
timestamp 1644511149
transform 1 0 22172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0590_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18124 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26864 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9752 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0594_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0595_
timestamp 1644511149
transform 1 0 13064 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0596_
timestamp 1644511149
transform 1 0 15916 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0597_
timestamp 1644511149
transform 1 0 16008 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0598_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0599_
timestamp 1644511149
transform 1 0 12972 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0600_
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0601_
timestamp 1644511149
transform 1 0 15548 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19872 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0604_
timestamp 1644511149
transform 1 0 26956 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0607_
timestamp 1644511149
transform 1 0 27324 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0608_
timestamp 1644511149
transform 1 0 25208 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1644511149
transform 1 0 27968 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0610_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0611_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1644511149
transform 1 0 28520 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0613_
timestamp 1644511149
transform 1 0 27324 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1644511149
transform 1 0 28428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0615_
timestamp 1644511149
transform 1 0 27876 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0616_
timestamp 1644511149
transform 1 0 26128 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0617_
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0618_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1644511149
transform 1 0 25484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0620_
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1644511149
transform 1 0 27232 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0622_
timestamp 1644511149
transform 1 0 26128 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0623_
timestamp 1644511149
transform 1 0 25484 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0625_
timestamp 1644511149
transform 1 0 21896 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1644511149
transform 1 0 17664 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1644511149
transform 1 0 15548 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0628_
timestamp 1644511149
transform 1 0 15732 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0629_
timestamp 1644511149
transform 1 0 15456 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0630_
timestamp 1644511149
transform 1 0 16192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0631_
timestamp 1644511149
transform 1 0 16928 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0633_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0634_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0635_
timestamp 1644511149
transform 1 0 15456 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16468 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16008 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0638_
timestamp 1644511149
transform 1 0 12052 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0640_
timestamp 1644511149
transform 1 0 15364 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0643_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12696 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0645_
timestamp 1644511149
transform 1 0 11592 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0646_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12788 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1644511149
transform 1 0 11960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0648_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1644511149
transform 1 0 12420 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0651_
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0652_
timestamp 1644511149
transform 1 0 10212 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0653_
timestamp 1644511149
transform 1 0 11776 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1644511149
transform 1 0 10396 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0655_
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1644511149
transform 1 0 12512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0657_
timestamp 1644511149
transform 1 0 14720 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0658_
timestamp 1644511149
transform 1 0 11408 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0659_
timestamp 1644511149
transform 1 0 10672 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0660_
timestamp 1644511149
transform 1 0 9660 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1644511149
transform 1 0 9844 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0662_
timestamp 1644511149
transform 1 0 10580 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0663_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9568 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0665_
timestamp 1644511149
transform 1 0 9844 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0666_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9660 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0667_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1644511149
transform 1 0 10120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0669_
timestamp 1644511149
transform 1 0 8832 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0670_
timestamp 1644511149
transform 1 0 14260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0672_
timestamp 1644511149
transform 1 0 15272 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0673_
timestamp 1644511149
transform 1 0 13432 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0674_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12144 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1644511149
transform 1 0 14260 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0676_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0677_
timestamp 1644511149
transform 1 0 13064 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1644511149
transform 1 0 15180 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0679_
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0680_
timestamp 1644511149
transform 1 0 13248 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1644511149
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0682_
timestamp 1644511149
transform 1 0 12788 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0684_
timestamp 1644511149
transform 1 0 16468 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0685_
timestamp 1644511149
transform 1 0 16744 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0686_
timestamp 1644511149
transform 1 0 16836 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0687_
timestamp 1644511149
transform 1 0 14720 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0688_
timestamp 1644511149
transform 1 0 19136 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0689_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1644511149
transform 1 0 18400 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0691_
timestamp 1644511149
transform 1 0 16744 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0692_
timestamp 1644511149
transform 1 0 16468 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1644511149
transform 1 0 19320 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0694_
timestamp 1644511149
transform 1 0 17388 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1644511149
transform 1 0 18308 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0696_
timestamp 1644511149
transform 1 0 17112 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0697_
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0698_
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1644511149
transform 1 0 19136 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0700_
timestamp 1644511149
transform 1 0 17112 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1644511149
transform 1 0 18584 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0702_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18032 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0703_
timestamp 1644511149
transform 1 0 18124 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0704_
timestamp 1644511149
transform 1 0 17204 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0705_
timestamp 1644511149
transform 1 0 23000 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1644511149
transform 1 0 22540 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0707_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0708_
timestamp 1644511149
transform 1 0 19504 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1644511149
transform 1 0 23184 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0710_
timestamp 1644511149
transform 1 0 18124 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0711_
timestamp 1644511149
transform 1 0 19320 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0712_
timestamp 1644511149
transform 1 0 20332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1644511149
transform 1 0 23460 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0714_
timestamp 1644511149
transform 1 0 20424 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0715_
timestamp 1644511149
transform 1 0 20516 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21344 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1644511149
transform 1 0 22632 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0718_
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0719_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 1644511149
transform 1 0 19596 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0721_
timestamp 1644511149
transform 1 0 24932 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0722_
timestamp 1644511149
transform 1 0 23552 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21528 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0725_
timestamp 1644511149
transform 1 0 22632 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0726_
timestamp 1644511149
transform 1 0 21988 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0727_
timestamp 1644511149
transform 1 0 22448 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0728_
timestamp 1644511149
transform 1 0 21528 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0729_
timestamp 1644511149
transform 1 0 19596 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0731_
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _0732_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0733_
timestamp 1644511149
transform 1 0 23644 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0734_
timestamp 1644511149
transform 1 0 20332 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0735_
timestamp 1644511149
transform 1 0 19228 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0736_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0737_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18032 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0738_
timestamp 1644511149
transform 1 0 23184 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0739_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0740_
timestamp 1644511149
transform 1 0 17020 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0741_
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _0742_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0743_
timestamp 1644511149
transform 1 0 24104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16836 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0745_
timestamp 1644511149
transform 1 0 17112 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0746_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0747_
timestamp 1644511149
transform 1 0 21528 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0748_
timestamp 1644511149
transform 1 0 20516 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0749_
timestamp 1644511149
transform 1 0 20516 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0750_
timestamp 1644511149
transform 1 0 20792 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0751_
timestamp 1644511149
transform 1 0 26220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0752_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21712 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20608 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1644511149
transform 1 0 20700 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0755_
timestamp 1644511149
transform 1 0 27140 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0756_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20240 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _0757_
timestamp 1644511149
transform 1 0 21804 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0758_
timestamp 1644511149
transform 1 0 27048 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0759_
timestamp 1644511149
transform 1 0 24932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0760_
timestamp 1644511149
transform 1 0 24840 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0761_
timestamp 1644511149
transform 1 0 23368 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0762_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0763_
timestamp 1644511149
transform 1 0 21252 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0764_
timestamp 1644511149
transform 1 0 25300 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 1644511149
transform 1 0 24564 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0766_
timestamp 1644511149
transform 1 0 23736 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0767_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1644511149
transform 1 0 24564 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0769_
timestamp 1644511149
transform 1 0 23736 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0770_
timestamp 1644511149
transform 1 0 24748 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0771_
timestamp 1644511149
transform 1 0 23092 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0772_
timestamp 1644511149
transform 1 0 27968 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _0773_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0774_
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0775_
timestamp 1644511149
transform 1 0 25208 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0776_
timestamp 1644511149
transform 1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0777_
timestamp 1644511149
transform 1 0 25944 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0778_
timestamp 1644511149
transform 1 0 25668 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0779_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26680 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0780_
timestamp 1644511149
transform 1 0 25760 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 1644511149
transform 1 0 26864 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0782_
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0783_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0784_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0785_
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0786_
timestamp 1644511149
transform 1 0 28336 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0787_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27508 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0788_
timestamp 1644511149
transform 1 0 27600 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0789_
timestamp 1644511149
transform 1 0 18400 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0790_
timestamp 1644511149
transform 1 0 28520 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0791_
timestamp 1644511149
transform 1 0 27784 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0792_
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0793_
timestamp 1644511149
transform 1 0 29900 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0794_
timestamp 1644511149
transform 1 0 30268 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0795_
timestamp 1644511149
transform 1 0 30912 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0796_
timestamp 1644511149
transform 1 0 29992 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0797_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0798_
timestamp 1644511149
transform 1 0 29624 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0799_
timestamp 1644511149
transform 1 0 29900 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0800_
timestamp 1644511149
transform 1 0 19320 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0801_
timestamp 1644511149
transform 1 0 25300 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0802_
timestamp 1644511149
transform 1 0 25392 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0803_
timestamp 1644511149
transform 1 0 17112 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0804_
timestamp 1644511149
transform 1 0 17940 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0805_
timestamp 1644511149
transform 1 0 18584 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0806_
timestamp 1644511149
transform 1 0 19136 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 1644511149
transform 1 0 20148 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0808_
timestamp 1644511149
transform 1 0 19320 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0809_
timestamp 1644511149
transform 1 0 17296 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0810_
timestamp 1644511149
transform 1 0 16376 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0811_
timestamp 1644511149
transform 1 0 15640 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1644511149
transform 1 0 17112 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0813_
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0814_
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0815_
timestamp 1644511149
transform 1 0 17572 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0816_
timestamp 1644511149
transform 1 0 17388 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0817_
timestamp 1644511149
transform 1 0 15364 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0818_
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0819_
timestamp 1644511149
transform 1 0 20516 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0820_
timestamp 1644511149
transform 1 0 19872 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0821_
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0822_
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0823_
timestamp 1644511149
transform 1 0 16652 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0824_
timestamp 1644511149
transform 1 0 17848 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0825_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0826_
timestamp 1644511149
transform 1 0 17204 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0827_
timestamp 1644511149
transform 1 0 17112 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0828_
timestamp 1644511149
transform 1 0 15732 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0829_
timestamp 1644511149
transform 1 0 17756 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0830_
timestamp 1644511149
transform 1 0 17572 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 1644511149
transform 1 0 17112 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0832_
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0834_
timestamp 1644511149
transform 1 0 28612 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 1644511149
transform 1 0 28428 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0836_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0837_
timestamp 1644511149
transform 1 0 29072 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0838_
timestamp 1644511149
transform 1 0 28152 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0839_
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0840_
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0841_
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0842_
timestamp 1644511149
transform 1 0 28796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0843_
timestamp 1644511149
transform 1 0 27876 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0844_
timestamp 1644511149
transform 1 0 27140 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0845_
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0846_
timestamp 1644511149
transform 1 0 29900 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0847_
timestamp 1644511149
transform 1 0 30820 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0848_
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0849_
timestamp 1644511149
transform 1 0 25392 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0850_
timestamp 1644511149
transform 1 0 25300 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0851_
timestamp 1644511149
transform 1 0 26404 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0852_
timestamp 1644511149
transform 1 0 24288 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0853_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0854_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0855_
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0856_
timestamp 1644511149
transform 1 0 25576 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0857_
timestamp 1644511149
transform 1 0 25668 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1644511149
transform 1 0 23092 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0859_
timestamp 1644511149
transform 1 0 22724 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0860_
timestamp 1644511149
transform 1 0 45540 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0861_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46000 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1644511149
transform 1 0 25760 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1644511149
transform 1 0 24748 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1644511149
transform 1 0 45540 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0871_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45080 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0873_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45264 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1644511149
transform 1 0 45816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0879_
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1644511149
transform 1 0 27508 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1644511149
transform 1 0 46828 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1644511149
transform 1 0 41676 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1644511149
transform 1 0 42872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0885_
timestamp 1644511149
transform 1 0 20976 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0886_
timestamp 1644511149
transform 1 0 20516 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1644511149
transform 1 0 15640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1644511149
transform 1 0 46736 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1644511149
transform 1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 30084 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0892_
timestamp 1644511149
transform 1 0 20148 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 20424 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0898_
timestamp 1644511149
transform 1 0 19688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 7636 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 7544 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 17480 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1644511149
transform 1 0 6900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 19688 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0904_
timestamp 1644511149
transform 1 0 21804 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 23460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 30452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1644511149
transform 1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 46736 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1644511149
transform 1 0 41032 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0916_
timestamp 1644511149
transform 1 0 20976 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0917_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 7544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0923_
timestamp 1644511149
transform 1 0 21344 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1644511149
transform 1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 43148 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0929_
timestamp 1644511149
transform 1 0 20424 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 23368 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 23736 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 21068 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0935_
timestamp 1644511149
transform 1 0 20516 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 10672 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 2116 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 2116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 45172 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 38272 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0941_
timestamp 1644511149
transform 1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 21160 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 15824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0947_
timestamp 1644511149
transform 1 0 41032 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0948_
timestamp 1644511149
transform 1 0 14996 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 14168 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 13340 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 12052 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 14812 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 14720 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0954_
timestamp 1644511149
transform 1 0 29900 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 29532 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 28428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 23920 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 23184 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0960_
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 46368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 42504 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0966_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 2024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0972_
timestamp 1644511149
transform 1 0 17940 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0979_
timestamp 1644511149
transform 1 0 20424 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0980_
timestamp 1644511149
transform 1 0 19688 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _0982_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _0983_
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0984_
timestamp 1644511149
transform 1 0 45080 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0985_
timestamp 1644511149
transform 1 0 45356 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0986_
timestamp 1644511149
transform 1 0 45264 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0987_
timestamp 1644511149
transform 1 0 46736 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0988_
timestamp 1644511149
transform 1 0 47748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0989_
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0990_
timestamp 1644511149
transform 1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0991_
timestamp 1644511149
transform 1 0 23000 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0992_
timestamp 1644511149
transform 1 0 23644 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _0993_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0994_
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0995_
timestamp 1644511149
transform 1 0 46368 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0996_
timestamp 1644511149
transform 1 0 45172 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0997_
timestamp 1644511149
transform 1 0 45816 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0998_
timestamp 1644511149
transform 1 0 45540 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _0999_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45264 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1000_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45816 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__and2b_1  _1001_
timestamp 1644511149
transform 1 0 45356 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1002_
timestamp 1644511149
transform 1 0 45080 0 -1 11968
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _1003_
timestamp 1644511149
transform 1 0 45816 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1004_
timestamp 1644511149
transform 1 0 46644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1005_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46184 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1006_
timestamp 1644511149
transform 1 0 47840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1007_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46276 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1008_
timestamp 1644511149
transform 1 0 22632 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1644511149
transform 1 0 24288 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1010_
timestamp 1644511149
transform 1 0 25024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1011_
timestamp 1644511149
transform 1 0 22724 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _1012_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1013_
timestamp 1644511149
transform 1 0 24472 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1014_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _1015_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1017_
timestamp 1644511149
transform 1 0 24288 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1018_
timestamp 1644511149
transform 1 0 24748 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1019_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45356 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1020_
timestamp 1644511149
transform 1 0 44344 0 -1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1021_
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _1022_
timestamp 1644511149
transform 1 0 17112 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 23552 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1644511149
transform 1 0 25484 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1644511149
transform 1 0 24472 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1644511149
transform 1 0 27416 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1644511149
transform 1 0 27876 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1644511149
transform 1 0 31004 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform 1 0 27600 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1644511149
transform 1 0 30176 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1644511149
transform 1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1032_
timestamp 1644511149
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1644511149
transform 1 0 15088 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 15456 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1644511149
transform 1 0 15364 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1038_
timestamp 1644511149
transform 1 0 25944 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1644511149
transform 1 0 15272 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1644511149
transform 1 0 16376 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 20148 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1644511149
transform 1 0 31280 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1644511149
transform 1 0 31188 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1044_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1644511149
transform 1 0 28520 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1644511149
transform 1 0 25760 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1644511149
transform 1 0 22540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1050_
timestamp 1644511149
transform 1 0 20976 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1644511149
transform 1 0 23184 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1644511149
transform 1 0 22540 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1644511149
transform 1 0 22632 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1644511149
transform 1 0 22448 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1056_
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1644511149
transform 1 0 18400 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1644511149
transform 1 0 20240 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1061_
timestamp 1644511149
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1062_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1063_
timestamp 1644511149
transform 1 0 17848 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1644511149
transform 1 0 18308 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1065_
timestamp 1644511149
transform 1 0 19596 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1066_
timestamp 1644511149
transform 1 0 18216 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1067_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1068_
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1069_
timestamp 1644511149
transform 1 0 12972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1070_
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1071_
timestamp 1644511149
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1644511149
transform 1 0 12420 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1073_
timestamp 1644511149
transform 1 0 12696 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1074_
timestamp 1644511149
transform 1 0 11408 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1075_
timestamp 1644511149
transform 1 0 9384 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1076_
timestamp 1644511149
transform 1 0 9844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1077_
timestamp 1644511149
transform 1 0 10672 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1079_
timestamp 1644511149
transform 1 0 10120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1080_
timestamp 1644511149
transform 1 0 9292 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1082_
timestamp 1644511149
transform 1 0 10304 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1083_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1085_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1086_
timestamp 1644511149
transform 1 0 14444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1087_
timestamp 1644511149
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1088_
timestamp 1644511149
transform 1 0 16376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1089_
timestamp 1644511149
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1090_
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1091_
timestamp 1644511149
transform 1 0 26496 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1092_
timestamp 1644511149
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1093_
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 26680 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1644511149
transform 1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1096_
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1097_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1644511149
transform 1 0 20148 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22080 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1100_
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1101_
timestamp 1644511149
transform 1 0 23460 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1103_
timestamp 1644511149
transform 1 0 30176 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1644511149
transform 1 0 26404 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 1644511149
transform 1 0 29072 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 1644511149
transform 1 0 29900 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1107_
timestamp 1644511149
transform 1 0 15548 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1108_
timestamp 1644511149
transform 1 0 14352 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 1644511149
transform 1 0 14352 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 1644511149
transform 1 0 14260 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 1644511149
transform 1 0 19044 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 1644511149
transform 1 0 14168 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 1644511149
transform 1 0 14168 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1114_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1115_
timestamp 1644511149
transform 1 0 30544 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1116_
timestamp 1644511149
transform 1 0 30176 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1117_
timestamp 1644511149
transform 1 0 27876 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 1644511149
transform 1 0 27600 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 1644511149
transform 1 0 24656 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1121_
timestamp 1644511149
transform 1 0 21252 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1122_
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1123_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1124_
timestamp 1644511149
transform 1 0 19596 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1125_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 1644511149
transform 1 0 20884 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 1644511149
transform 1 0 16376 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 1644511149
transform 1 0 17480 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1131_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20884 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1133_
timestamp 1644511149
transform 1 0 17480 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1134_
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 1644511149
transform 1 0 16928 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1136_
timestamp 1644511149
transform 1 0 18400 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 1644511149
transform 1 0 17112 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1139_
timestamp 1644511149
transform 1 0 13156 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1140_
timestamp 1644511149
transform 1 0 12696 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1141_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1142_
timestamp 1644511149
transform 1 0 12052 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1143_
timestamp 1644511149
transform 1 0 9016 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1144_
timestamp 1644511149
transform 1 0 11316 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1145_
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1146_
timestamp 1644511149
transform 1 0 10304 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1147_
timestamp 1644511149
transform 1 0 9384 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1148_
timestamp 1644511149
transform 1 0 11224 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1149_
timestamp 1644511149
transform 1 0 10488 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1150_
timestamp 1644511149
transform 1 0 12880 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1151_
timestamp 1644511149
transform 1 0 13064 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1152_
timestamp 1644511149
transform 1 0 14352 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1153_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1154_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1155_
timestamp 1644511149
transform 1 0 21988 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1156_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1157_
timestamp 1644511149
transform 1 0 24564 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1644511149
transform 1 0 27232 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1159_
timestamp 1644511149
transform 1 0 27784 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 1644511149
transform 1 0 25208 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1162_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1163_
timestamp 1644511149
transform 1 0 18584 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1164__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47472 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1165__82
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1166__83
timestamp 1644511149
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1167__84
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1168__85
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1169__86
timestamp 1644511149
transform 1 0 20884 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1170__87
timestamp 1644511149
transform 1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1171__88
timestamp 1644511149
transform 1 0 25300 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1172__89
timestamp 1644511149
transform 1 0 10580 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1173__90
timestamp 1644511149
transform 1 0 25944 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1174__91
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1175__92
timestamp 1644511149
transform 1 0 2116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1176__93
timestamp 1644511149
transform 1 0 33672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1177__94
timestamp 1644511149
transform 1 0 4140 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1178__95
timestamp 1644511149
transform 1 0 1656 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1179__96
timestamp 1644511149
transform 1 0 43792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1180__97
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1181__98
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1182__99
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1183__100
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1184__101
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1185__102
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1186__103
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1187__104
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1188__105
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1189__106
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1190__107
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1191__108
timestamp 1644511149
transform 1 0 45816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1192__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1193__110
timestamp 1644511149
transform 1 0 45632 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1194__111
timestamp 1644511149
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1195__112
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1196__113
timestamp 1644511149
transform 1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1197__114
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1198__115
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1199__116
timestamp 1644511149
transform 1 0 42688 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1200__117
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1201__118
timestamp 1644511149
transform 1 0 12972 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1202__119
timestamp 1644511149
transform 1 0 6716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1203__120
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1204__121
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1205__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1206__123
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1207__124
timestamp 1644511149
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1208__125
timestamp 1644511149
transform 1 0 46184 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1209__126
timestamp 1644511149
transform 1 0 19872 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1210__127
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1211__128
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1212__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1213__130
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1214__131
timestamp 1644511149
transform 1 0 1840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1215__132
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1216__133
timestamp 1644511149
transform 1 0 7268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1217__134
timestamp 1644511149
transform 1 0 45632 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1218__135
timestamp 1644511149
transform 1 0 43884 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24472 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1220_
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1221_
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1222_
timestamp 1644511149
transform 1 0 45172 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1223_
timestamp 1644511149
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1224_
timestamp 1644511149
transform 1 0 21712 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1225_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1226_
timestamp 1644511149
transform 1 0 26404 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1227_
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1228_
timestamp 1644511149
transform 1 0 46276 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1229_
timestamp 1644511149
transform 1 0 31648 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1230_
timestamp 1644511149
transform 1 0 19964 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1231_
timestamp 1644511149
transform 1 0 46276 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1232_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1233_
timestamp 1644511149
transform 1 0 20884 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1234_
timestamp 1644511149
transform 1 0 10304 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1235_
timestamp 1644511149
transform 1 0 25208 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1236_
timestamp 1644511149
transform 1 0 10580 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1237_
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1238_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1239_
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1240_
timestamp 1644511149
transform 1 0 32936 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1241_
timestamp 1644511149
transform 1 0 3956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1242_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1243_
timestamp 1644511149
transform 1 0 42688 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1244_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1245_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1246_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1247_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1248_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1249_
timestamp 1644511149
transform 1 0 7912 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1250_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1251_
timestamp 1644511149
transform 1 0 46184 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1252_
timestamp 1644511149
transform 1 0 21804 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1253_
timestamp 1644511149
transform 1 0 10672 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1254_
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1255_
timestamp 1644511149
transform 1 0 15916 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1256_
timestamp 1644511149
transform 1 0 20516 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1257_
timestamp 1644511149
transform 1 0 14996 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1258_
timestamp 1644511149
transform 1 0 15088 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1259_
timestamp 1644511149
transform 1 0 20240 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1260_
timestamp 1644511149
transform 1 0 29992 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1261_
timestamp 1644511149
transform 1 0 15732 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1262_
timestamp 1644511149
transform 1 0 7268 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1263_
timestamp 1644511149
transform 1 0 9660 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1264_
timestamp 1644511149
transform 1 0 15640 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1265_
timestamp 1644511149
transform 1 0 7544 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1266_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1267_
timestamp 1644511149
transform 1 0 14076 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1268_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1269_
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1270_
timestamp 1644511149
transform 1 0 12972 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1271_
timestamp 1644511149
transform 1 0 12788 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1272_
timestamp 1644511149
transform 1 0 17388 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1273_
timestamp 1644511149
transform 1 0 19136 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1274_
timestamp 1644511149
transform 1 0 14260 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1275_
timestamp 1644511149
transform 1 0 21896 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1276_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1277_
timestamp 1644511149
transform 1 0 24196 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1278_
timestamp 1644511149
transform 1 0 29716 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1279_
timestamp 1644511149
transform 1 0 30360 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1280_
timestamp 1644511149
transform 1 0 29072 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1281_
timestamp 1644511149
transform 1 0 22816 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1282_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1283_
timestamp 1644511149
transform 1 0 9108 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1284_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1285_
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1286_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1644511149
transform 1 0 41308 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1644511149
transform 1 0 24564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1644511149
transform 1 0 42596 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1644511149
transform 1 0 13616 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1644511149
transform 1 0 6716 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 13524 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1644511149
transform 1 0 45172 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1309_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1310_
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1311_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1312_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1313_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1314_
timestamp 1644511149
transform 1 0 42596 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 19596 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 19688 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 26864 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1644511149
transform 1 0 47656 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 12972 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 47932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 45724 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1644511149
transform 1 0 44160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1644511149
transform 1 0 1748 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1644511149
transform 1 0 47288 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1644511149
transform 1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1644511149
transform 1 0 40020 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1644511149
transform 1 0 47840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 47656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input33
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1644511149
transform 1 0 47748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1644511149
transform 1 0 47288 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1644511149
transform 1 0 47840 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1644511149
transform 1 0 9292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1644511149
transform 1 0 12328 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1644511149
transform 1 0 20056 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 46460 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1644511149
transform 1 0 47656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 30728 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 45356 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 27324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1644511149
transform 1 0 11684 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 46184 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 46184 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1644511149
transform 1 0 47288 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1644511149
transform 1 0 46460 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1644511149
transform 1 0 47932 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 23276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 6716 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41124 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 41492 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 38456 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 39560 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 40480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 18768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 19320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 19872 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 21344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 23276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 23828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 22172 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[0\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 24840 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 29256 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 15272 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 20884 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2300 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35880 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 45908 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 45172 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 25392 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 25208 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 20608 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 25576 0 1 40256
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
