magic
tech sky130A
magscale 1 2
timestamp 1654174284
<< viali >>
rect 29929 47209 29963 47243
rect 13369 47141 13403 47175
rect 19441 47141 19475 47175
rect 47961 47141 47995 47175
rect 11713 47073 11747 47107
rect 20085 47073 20119 47107
rect 30757 47073 30791 47107
rect 44465 47073 44499 47107
rect 47041 47073 47075 47107
rect 1961 47005 1995 47039
rect 2697 47005 2731 47039
rect 3801 47005 3835 47039
rect 4813 47005 4847 47039
rect 6837 47005 6871 47039
rect 7757 47005 7791 47039
rect 9413 47005 9447 47039
rect 11989 47005 12023 47039
rect 13093 47005 13127 47039
rect 14565 47005 14599 47039
rect 16681 47005 16715 47039
rect 16957 47005 16991 47039
rect 19257 47005 19291 47039
rect 20361 47005 20395 47039
rect 25697 47005 25731 47039
rect 28641 47005 28675 47039
rect 29745 47005 29779 47039
rect 31033 47005 31067 47039
rect 38393 47005 38427 47039
rect 42625 47005 42659 47039
rect 45201 47005 45235 47039
rect 47777 47005 47811 47039
rect 4077 46937 4111 46971
rect 7941 46937 7975 46971
rect 9597 46937 9631 46971
rect 14749 46937 14783 46971
rect 40325 46937 40359 46971
rect 40509 46937 40543 46971
rect 42809 46937 42843 46971
rect 45385 46937 45419 46971
rect 2145 46869 2179 46903
rect 2881 46869 2915 46903
rect 4905 46869 4939 46903
rect 6929 46869 6963 46903
rect 28457 46869 28491 46903
rect 28457 46597 28491 46631
rect 1409 46529 1443 46563
rect 12449 46529 12483 46563
rect 28273 46529 28307 46563
rect 38117 46529 38151 46563
rect 47869 46529 47903 46563
rect 13645 46461 13679 46495
rect 13829 46461 13863 46495
rect 14289 46461 14323 46495
rect 18981 46461 19015 46495
rect 19441 46461 19475 46495
rect 19625 46461 19659 46495
rect 20637 46461 20671 46495
rect 24593 46461 24627 46495
rect 24777 46461 24811 46495
rect 25789 46461 25823 46495
rect 30113 46461 30147 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 41889 46461 41923 46495
rect 42441 46461 42475 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46857 46461 46891 46495
rect 27169 46393 27203 46427
rect 1593 46325 1627 46359
rect 2329 46325 2363 46359
rect 4445 46325 4479 46359
rect 10701 46325 10735 46359
rect 12541 46325 12575 46359
rect 22017 46325 22051 46359
rect 32321 46325 32355 46359
rect 41245 46325 41279 46359
rect 48053 46325 48087 46359
rect 13553 46121 13587 46155
rect 14197 46121 14231 46155
rect 18613 46121 18647 46155
rect 38301 46121 38335 46155
rect 1409 45985 1443 46019
rect 2789 45985 2823 46019
rect 4169 45985 4203 46019
rect 4721 45985 4755 46019
rect 10425 45985 10459 46019
rect 11069 45985 11103 46019
rect 20085 45985 20119 46019
rect 21281 45985 21315 46019
rect 25421 45985 25455 46019
rect 25881 45985 25915 46019
rect 31677 45985 31711 46019
rect 32229 45985 32263 46019
rect 41245 45985 41279 46019
rect 41889 45985 41923 46019
rect 47041 45985 47075 46019
rect 14105 45917 14139 45951
rect 18521 45917 18555 45951
rect 19441 45917 19475 45951
rect 38209 45917 38243 45951
rect 43913 45917 43947 45951
rect 45661 45917 45695 45951
rect 46305 45917 46339 45951
rect 1593 45849 1627 45883
rect 4353 45849 4387 45883
rect 10609 45849 10643 45883
rect 19533 45849 19567 45883
rect 20269 45849 20303 45883
rect 25605 45849 25639 45883
rect 31861 45849 31895 45883
rect 41429 45849 41463 45883
rect 46489 45849 46523 45883
rect 44097 45781 44131 45815
rect 45753 45781 45787 45815
rect 2329 45577 2363 45611
rect 5089 45577 5123 45611
rect 10609 45577 10643 45611
rect 32229 45577 32263 45611
rect 41429 45577 41463 45611
rect 25421 45509 25455 45543
rect 27077 45509 27111 45543
rect 45109 45509 45143 45543
rect 47685 45509 47719 45543
rect 2237 45441 2271 45475
rect 4997 45441 5031 45475
rect 10517 45441 10551 45475
rect 25329 45441 25363 45475
rect 26985 45441 27019 45475
rect 32137 45441 32171 45475
rect 41337 45441 41371 45475
rect 46213 45441 46247 45475
rect 47593 45441 47627 45475
rect 42717 45373 42751 45407
rect 42901 45373 42935 45407
rect 44097 45373 44131 45407
rect 46489 45373 46523 45407
rect 45201 45237 45235 45271
rect 42073 45033 42107 45067
rect 43177 45033 43211 45067
rect 43821 45033 43855 45067
rect 45753 45033 45787 45067
rect 45201 44965 45235 44999
rect 48145 44897 48179 44931
rect 28181 44829 28215 44863
rect 41981 44829 42015 44863
rect 43085 44829 43119 44863
rect 43729 44829 43763 44863
rect 45661 44829 45695 44863
rect 46305 44829 46339 44863
rect 46489 44761 46523 44795
rect 28273 44693 28307 44727
rect 46029 44489 46063 44523
rect 46673 44489 46707 44523
rect 28089 44421 28123 44455
rect 42901 44353 42935 44387
rect 45477 44353 45511 44387
rect 45937 44353 45971 44387
rect 46581 44353 46615 44387
rect 47593 44353 47627 44387
rect 27905 44285 27939 44319
rect 28365 44285 28399 44319
rect 38669 44285 38703 44319
rect 38853 44285 38887 44319
rect 40049 44285 40083 44319
rect 44005 44285 44039 44319
rect 47685 44149 47719 44183
rect 38853 43945 38887 43979
rect 27353 43809 27387 43843
rect 29653 43809 29687 43843
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 27169 43741 27203 43775
rect 29561 43741 29595 43775
rect 38761 43741 38795 43775
rect 45845 43741 45879 43775
rect 46305 43741 46339 43775
rect 29009 43673 29043 43707
rect 27169 43333 27203 43367
rect 1409 43265 1443 43299
rect 26249 43265 26283 43299
rect 46305 43265 46339 43299
rect 46949 43265 46983 43299
rect 26985 43197 27019 43231
rect 28825 43197 28859 43231
rect 1593 43061 1627 43095
rect 26341 43061 26375 43095
rect 47777 43061 47811 43095
rect 46305 42721 46339 42755
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 47685 42313 47719 42347
rect 27169 42245 27203 42279
rect 46857 42177 46891 42211
rect 47593 42177 47627 42211
rect 26985 42109 27019 42143
rect 28825 42109 28859 42143
rect 2053 41973 2087 42007
rect 46949 41973 46983 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46489 41633 46523 41667
rect 46305 41565 46339 41599
rect 1593 41497 1627 41531
rect 48145 41497 48179 41531
rect 2145 41225 2179 41259
rect 2053 41089 2087 41123
rect 46213 41089 46247 41123
rect 47777 41089 47811 41123
rect 46489 41021 46523 41055
rect 46305 40545 46339 40579
rect 1869 40409 1903 40443
rect 2053 40409 2087 40443
rect 46489 40409 46523 40443
rect 48145 40409 48179 40443
rect 18981 40069 19015 40103
rect 18429 40001 18463 40035
rect 43637 40001 43671 40035
rect 44373 40001 44407 40035
rect 44925 40001 44959 40035
rect 45845 40001 45879 40035
rect 47777 40001 47811 40035
rect 43729 39933 43763 39967
rect 46121 39865 46155 39899
rect 18613 39457 18647 39491
rect 22753 39457 22787 39491
rect 46305 39457 46339 39491
rect 17049 39389 17083 39423
rect 18061 39389 18095 39423
rect 19257 39389 19291 39423
rect 17325 39321 17359 39355
rect 20085 39321 20119 39355
rect 46489 39321 46523 39355
rect 48145 39321 48179 39355
rect 22201 39253 22235 39287
rect 22569 39253 22603 39287
rect 22661 39253 22695 39287
rect 23581 39049 23615 39083
rect 47685 39049 47719 39083
rect 18429 38913 18463 38947
rect 25789 38913 25823 38947
rect 30297 38913 30331 38947
rect 45661 38913 45695 38947
rect 45845 38913 45879 38947
rect 46397 38913 46431 38947
rect 47593 38913 47627 38947
rect 19165 38845 19199 38879
rect 21833 38845 21867 38879
rect 22109 38845 22143 38879
rect 46857 38845 46891 38879
rect 25605 38709 25639 38743
rect 30481 38709 30515 38743
rect 45661 38709 45695 38743
rect 18337 38505 18371 38539
rect 22845 38505 22879 38539
rect 26985 38505 27019 38539
rect 19257 38437 19291 38471
rect 19901 38369 19935 38403
rect 23489 38369 23523 38403
rect 24593 38369 24627 38403
rect 27537 38369 27571 38403
rect 45109 38369 45143 38403
rect 45477 38369 45511 38403
rect 17601 38301 17635 38335
rect 17969 38301 18003 38335
rect 18521 38301 18555 38335
rect 19625 38301 19659 38335
rect 20545 38301 20579 38335
rect 22017 38301 22051 38335
rect 26709 38301 26743 38335
rect 27353 38301 27387 38335
rect 44281 38301 44315 38335
rect 44465 38301 44499 38335
rect 45293 38301 45327 38335
rect 46029 38301 46063 38335
rect 46397 38301 46431 38335
rect 23213 38233 23247 38267
rect 24869 38233 24903 38267
rect 44373 38233 44407 38267
rect 47869 38233 47903 38267
rect 17417 38165 17451 38199
rect 19717 38165 19751 38199
rect 20637 38165 20671 38199
rect 21833 38165 21867 38199
rect 23305 38165 23339 38199
rect 26341 38165 26375 38199
rect 27445 38165 27479 38199
rect 22017 37961 22051 37995
rect 23121 37961 23155 37995
rect 24501 37961 24535 37995
rect 25237 37961 25271 37995
rect 46029 37961 46063 37995
rect 17141 37893 17175 37927
rect 21925 37825 21959 37859
rect 22753 37825 22787 37859
rect 24225 37825 24259 37859
rect 25145 37825 25179 37859
rect 26065 37825 26099 37859
rect 26985 37825 27019 37859
rect 45753 37825 45787 37859
rect 46121 37825 46155 37859
rect 46673 37825 46707 37859
rect 16865 37757 16899 37791
rect 19533 37757 19567 37791
rect 19809 37757 19843 37791
rect 22845 37757 22879 37791
rect 26157 37757 26191 37791
rect 26433 37757 26467 37791
rect 28181 37757 28215 37791
rect 28457 37757 28491 37791
rect 45569 37757 45603 37791
rect 18613 37621 18647 37655
rect 21281 37621 21315 37655
rect 27169 37621 27203 37655
rect 29929 37621 29963 37655
rect 46765 37621 46799 37655
rect 47777 37621 47811 37655
rect 28917 37417 28951 37451
rect 29653 37417 29687 37451
rect 45753 37417 45787 37451
rect 18705 37349 18739 37383
rect 20545 37349 20579 37383
rect 22109 37349 22143 37383
rect 18245 37281 18279 37315
rect 20085 37281 20119 37315
rect 22201 37281 22235 37315
rect 28549 37281 28583 37315
rect 46489 37281 46523 37315
rect 48145 37281 48179 37315
rect 2053 37213 2087 37247
rect 18337 37213 18371 37247
rect 19809 37213 19843 37247
rect 19993 37213 20027 37247
rect 20177 37213 20211 37247
rect 20361 37213 20395 37247
rect 21925 37213 21959 37247
rect 22845 37213 22879 37247
rect 28181 37213 28215 37247
rect 28365 37213 28399 37247
rect 28457 37213 28491 37247
rect 28733 37213 28767 37247
rect 29561 37213 29595 37247
rect 45661 37213 45695 37247
rect 45845 37213 45879 37247
rect 46305 37213 46339 37247
rect 22661 37145 22695 37179
rect 21741 37077 21775 37111
rect 23029 37077 23063 37111
rect 17785 36873 17819 36907
rect 21281 36873 21315 36907
rect 22477 36873 22511 36907
rect 30849 36805 30883 36839
rect 1777 36737 1811 36771
rect 17693 36737 17727 36771
rect 20729 36737 20763 36771
rect 21097 36737 21131 36771
rect 22293 36737 22327 36771
rect 23121 36737 23155 36771
rect 24317 36737 24351 36771
rect 28549 36737 28583 36771
rect 30757 36737 30791 36771
rect 1961 36669 1995 36703
rect 2789 36669 2823 36703
rect 28825 36669 28859 36703
rect 21097 36533 21131 36567
rect 23213 36533 23247 36567
rect 24409 36533 24443 36567
rect 30297 36533 30331 36567
rect 2237 36329 2271 36363
rect 16589 36193 16623 36227
rect 23489 36193 23523 36227
rect 25421 36193 25455 36227
rect 25697 36193 25731 36227
rect 2145 36125 2179 36159
rect 16313 36125 16347 36159
rect 22385 36125 22419 36159
rect 23121 36125 23155 36159
rect 23305 36125 23339 36159
rect 23397 36125 23431 36159
rect 23673 36125 23707 36159
rect 29745 36125 29779 36159
rect 29929 36125 29963 36159
rect 30021 36125 30055 36159
rect 27997 36057 28031 36091
rect 28181 36057 28215 36091
rect 18061 35989 18095 36023
rect 22569 35989 22603 36023
rect 23857 35989 23891 36023
rect 27169 35989 27203 36023
rect 29561 35989 29595 36023
rect 17325 35785 17359 35819
rect 19441 35785 19475 35819
rect 25145 35785 25179 35819
rect 27077 35785 27111 35819
rect 27721 35785 27755 35819
rect 29469 35785 29503 35819
rect 23673 35717 23707 35751
rect 1593 35649 1627 35683
rect 17233 35649 17267 35683
rect 17877 35649 17911 35683
rect 18061 35649 18095 35683
rect 18705 35649 18739 35683
rect 18889 35649 18923 35683
rect 18981 35649 19015 35683
rect 19257 35649 19291 35683
rect 22477 35649 22511 35683
rect 22569 35649 22603 35683
rect 22845 35649 22879 35683
rect 26985 35649 27019 35683
rect 27905 35649 27939 35683
rect 27997 35649 28031 35683
rect 28140 35649 28174 35683
rect 28263 35671 28297 35705
rect 28733 35649 28767 35683
rect 28917 35651 28951 35685
rect 29009 35649 29043 35683
rect 29285 35649 29319 35683
rect 29929 35649 29963 35683
rect 30941 35649 30975 35683
rect 32137 35649 32171 35683
rect 19073 35581 19107 35615
rect 23397 35581 23431 35615
rect 29101 35581 29135 35615
rect 30021 35581 30055 35615
rect 31033 35581 31067 35615
rect 30297 35513 30331 35547
rect 31309 35513 31343 35547
rect 1409 35445 1443 35479
rect 18245 35445 18279 35479
rect 22293 35445 22327 35479
rect 22753 35445 22787 35479
rect 30113 35445 30147 35479
rect 32229 35445 32263 35479
rect 18245 35241 18279 35275
rect 19625 35241 19659 35275
rect 19809 35241 19843 35275
rect 22477 35241 22511 35275
rect 23489 35241 23523 35275
rect 25421 35241 25455 35275
rect 26801 35241 26835 35275
rect 27261 35241 27295 35275
rect 28549 35241 28583 35275
rect 29009 35241 29043 35275
rect 29653 35241 29687 35275
rect 17325 35173 17359 35207
rect 23673 35173 23707 35207
rect 18337 35105 18371 35139
rect 19533 35105 19567 35139
rect 20729 35105 20763 35139
rect 25237 35105 25271 35139
rect 26525 35105 26559 35139
rect 27353 35105 27387 35139
rect 29745 35105 29779 35139
rect 31125 35105 31159 35139
rect 17509 35037 17543 35071
rect 17693 35037 17727 35071
rect 17785 35037 17819 35071
rect 18521 35037 18555 35071
rect 19257 35037 19291 35071
rect 23121 35037 23155 35071
rect 23397 35037 23431 35071
rect 25421 35037 25455 35071
rect 26617 35037 26651 35071
rect 27537 35037 27571 35071
rect 28457 35037 28491 35071
rect 28825 35037 28859 35071
rect 29837 35037 29871 35071
rect 48145 35037 48179 35071
rect 18245 34969 18279 35003
rect 21005 34969 21039 35003
rect 25145 34969 25179 35003
rect 27261 34969 27295 35003
rect 29561 34969 29595 35003
rect 31401 34969 31435 35003
rect 18705 34901 18739 34935
rect 25605 34901 25639 34935
rect 26157 34901 26191 34935
rect 27721 34901 27755 34935
rect 30021 34901 30055 34935
rect 32873 34901 32907 34935
rect 47961 34901 47995 34935
rect 18613 34697 18647 34731
rect 19533 34697 19567 34731
rect 21189 34697 21223 34731
rect 24961 34697 24995 34731
rect 28181 34697 28215 34731
rect 28733 34697 28767 34731
rect 30205 34697 30239 34731
rect 17325 34629 17359 34663
rect 18153 34629 18187 34663
rect 19073 34629 19107 34663
rect 25973 34629 26007 34663
rect 26985 34629 27019 34663
rect 17141 34561 17175 34595
rect 17417 34561 17451 34595
rect 18337 34561 18371 34595
rect 18429 34561 18463 34595
rect 19257 34561 19291 34595
rect 19349 34561 19383 34595
rect 20255 34561 20289 34595
rect 21097 34561 21131 34595
rect 22661 34561 22695 34595
rect 25145 34561 25179 34595
rect 25329 34561 25363 34595
rect 26157 34561 26191 34595
rect 27261 34561 27295 34595
rect 27905 34561 27939 34595
rect 27997 34561 28031 34595
rect 28641 34561 28675 34595
rect 28825 34561 28859 34595
rect 29837 34561 29871 34595
rect 30021 34561 30055 34595
rect 31217 34561 31251 34595
rect 31309 34561 31343 34595
rect 31585 34561 31619 34595
rect 48145 34561 48179 34595
rect 20085 34493 20119 34527
rect 22385 34493 22419 34527
rect 25421 34493 25455 34527
rect 26341 34493 26375 34527
rect 27077 34493 27111 34527
rect 28181 34493 28215 34527
rect 31493 34493 31527 34527
rect 16957 34357 16991 34391
rect 18429 34357 18463 34391
rect 19073 34357 19107 34391
rect 20453 34357 20487 34391
rect 27169 34357 27203 34391
rect 27445 34357 27479 34391
rect 31033 34357 31067 34391
rect 47961 34357 47995 34391
rect 17969 34153 18003 34187
rect 19441 34153 19475 34187
rect 21373 34153 21407 34187
rect 21741 34153 21775 34187
rect 22477 34153 22511 34187
rect 24961 34153 24995 34187
rect 31033 34153 31067 34187
rect 31401 34153 31435 34187
rect 19625 34085 19659 34119
rect 27537 34085 27571 34119
rect 15945 34017 15979 34051
rect 17417 34017 17451 34051
rect 31493 34017 31527 34051
rect 47133 34017 47167 34051
rect 47409 34017 47443 34051
rect 1593 33949 1627 33983
rect 15669 33949 15703 33983
rect 18153 33949 18187 33983
rect 18337 33949 18371 33983
rect 18429 33949 18463 33983
rect 21557 33949 21591 33983
rect 21833 33949 21867 33983
rect 23673 33949 23707 33983
rect 26065 33949 26099 33983
rect 26249 33949 26283 33983
rect 27997 33949 28031 33983
rect 28181 33949 28215 33983
rect 29929 33949 29963 33983
rect 30113 33949 30147 33983
rect 31217 33949 31251 33983
rect 31953 33949 31987 33983
rect 32137 33949 32171 33983
rect 19257 33881 19291 33915
rect 22385 33881 22419 33915
rect 24869 33881 24903 33915
rect 27353 33881 27387 33915
rect 30021 33881 30055 33915
rect 47225 33881 47259 33915
rect 1409 33813 1443 33847
rect 19457 33813 19491 33847
rect 23765 33813 23799 33847
rect 26157 33813 26191 33847
rect 28089 33813 28123 33847
rect 32045 33813 32079 33847
rect 16037 33609 16071 33643
rect 17693 33609 17727 33643
rect 18613 33609 18647 33643
rect 19257 33609 19291 33643
rect 26173 33609 26207 33643
rect 26341 33609 26375 33643
rect 28549 33609 28583 33643
rect 17417 33541 17451 33575
rect 22201 33541 22235 33575
rect 25973 33541 26007 33575
rect 26985 33541 27019 33575
rect 30941 33541 30975 33575
rect 31033 33541 31067 33575
rect 15945 33473 15979 33507
rect 17141 33473 17175 33507
rect 17325 33473 17359 33507
rect 17509 33473 17543 33507
rect 18521 33473 18555 33507
rect 18705 33473 18739 33507
rect 19165 33473 19199 33507
rect 19349 33473 19383 33507
rect 22845 33473 22879 33507
rect 25421 33473 25455 33507
rect 25513 33473 25547 33507
rect 27169 33473 27203 33507
rect 28457 33473 28491 33507
rect 29101 33473 29135 33507
rect 30665 33473 30699 33507
rect 30813 33473 30847 33507
rect 31171 33473 31205 33507
rect 32137 33473 32171 33507
rect 47777 33473 47811 33507
rect 1409 33405 1443 33439
rect 1685 33405 1719 33439
rect 23121 33405 23155 33439
rect 24593 33405 24627 33439
rect 25053 33405 25087 33439
rect 48053 33405 48087 33439
rect 22293 33269 22327 33303
rect 25237 33269 25271 33303
rect 26157 33269 26191 33303
rect 27353 33269 27387 33303
rect 29193 33269 29227 33303
rect 31309 33269 31343 33303
rect 32229 33269 32263 33303
rect 22753 33065 22787 33099
rect 25605 33065 25639 33099
rect 25697 33065 25731 33099
rect 26801 33065 26835 33099
rect 29009 33065 29043 33099
rect 32781 33065 32815 33099
rect 23121 32997 23155 33031
rect 1409 32929 1443 32963
rect 1593 32929 1627 32963
rect 27261 32929 27295 32963
rect 31033 32929 31067 32963
rect 31309 32929 31343 32963
rect 16773 32861 16807 32895
rect 17417 32861 17451 32895
rect 18521 32861 18555 32895
rect 18705 32861 18739 32895
rect 19257 32861 19291 32895
rect 21281 32861 21315 32895
rect 22937 32861 22971 32895
rect 23213 32861 23247 32895
rect 25513 32861 25547 32895
rect 25789 32861 25823 32895
rect 25973 32861 26007 32895
rect 26617 32861 26651 32895
rect 30021 32861 30055 32895
rect 46305 32861 46339 32895
rect 3249 32793 3283 32827
rect 19349 32793 19383 32827
rect 25237 32793 25271 32827
rect 26433 32793 26467 32827
rect 27537 32793 27571 32827
rect 46489 32793 46523 32827
rect 48145 32793 48179 32827
rect 16865 32725 16899 32759
rect 17509 32725 17543 32759
rect 18613 32725 18647 32759
rect 21465 32725 21499 32759
rect 30113 32725 30147 32759
rect 18429 32521 18463 32555
rect 19073 32521 19107 32555
rect 25973 32521 26007 32555
rect 27629 32521 27663 32555
rect 30849 32521 30883 32555
rect 47685 32521 47719 32555
rect 2329 32453 2363 32487
rect 20085 32453 20119 32487
rect 25145 32453 25179 32487
rect 27077 32453 27111 32487
rect 16681 32385 16715 32419
rect 19070 32385 19104 32419
rect 21097 32385 21131 32419
rect 21189 32385 21223 32419
rect 22017 32385 22051 32419
rect 22477 32385 22511 32419
rect 23213 32385 23247 32419
rect 23857 32385 23891 32419
rect 24685 32385 24719 32419
rect 24869 32385 24903 32419
rect 25053 32385 25087 32419
rect 25914 32385 25948 32419
rect 26341 32385 26375 32419
rect 26985 32385 27019 32419
rect 27169 32385 27203 32419
rect 27813 32385 27847 32419
rect 27997 32385 28031 32419
rect 28089 32385 28123 32419
rect 30665 32385 30699 32419
rect 47041 32385 47075 32419
rect 47593 32385 47627 32419
rect 2145 32317 2179 32351
rect 3249 32317 3283 32351
rect 16957 32317 16991 32351
rect 19533 32317 19567 32351
rect 22201 32317 22235 32351
rect 22293 32317 22327 32351
rect 23397 32317 23431 32351
rect 26433 32317 26467 32351
rect 30481 32317 30515 32351
rect 22109 32249 22143 32283
rect 25789 32249 25823 32283
rect 1685 32181 1719 32215
rect 18889 32181 18923 32215
rect 19441 32181 19475 32215
rect 20177 32181 20211 32215
rect 21833 32181 21867 32215
rect 23949 32181 23983 32215
rect 18061 31977 18095 32011
rect 26525 31977 26559 32011
rect 30113 31977 30147 32011
rect 17969 31909 18003 31943
rect 19257 31909 19291 31943
rect 22937 31909 22971 31943
rect 27721 31909 27755 31943
rect 28457 31909 28491 31943
rect 31217 31909 31251 31943
rect 1409 31841 1443 31875
rect 1869 31841 1903 31875
rect 17325 31841 17359 31875
rect 18153 31841 18187 31875
rect 19441 31841 19475 31875
rect 19533 31841 19567 31875
rect 19625 31841 19659 31875
rect 20545 31841 20579 31875
rect 20821 31841 20855 31875
rect 22293 31841 22327 31875
rect 22753 31841 22787 31875
rect 47317 31841 47351 31875
rect 17049 31773 17083 31807
rect 17141 31773 17175 31807
rect 17417 31773 17451 31807
rect 17877 31773 17911 31807
rect 19717 31773 19751 31807
rect 23213 31773 23247 31807
rect 25237 31773 25271 31807
rect 28273 31773 28307 31807
rect 30665 31773 30699 31807
rect 30941 31773 30975 31807
rect 31033 31773 31067 31807
rect 47593 31773 47627 31807
rect 1593 31705 1627 31739
rect 23121 31705 23155 31739
rect 27537 31705 27571 31739
rect 30021 31705 30055 31739
rect 30849 31705 30883 31739
rect 16865 31637 16899 31671
rect 2329 31433 2363 31467
rect 18429 31433 18463 31467
rect 18889 31433 18923 31467
rect 23213 31433 23247 31467
rect 23581 31433 23615 31467
rect 27905 31433 27939 31467
rect 29561 31433 29595 31467
rect 16957 31365 16991 31399
rect 22385 31365 22419 31399
rect 22477 31365 22511 31399
rect 27261 31365 27295 31399
rect 32505 31365 32539 31399
rect 2237 31297 2271 31331
rect 19073 31297 19107 31331
rect 21005 31297 21039 31331
rect 22109 31297 22143 31331
rect 22202 31297 22236 31331
rect 22574 31297 22608 31331
rect 23397 31297 23431 31331
rect 23673 31297 23707 31331
rect 25513 31297 25547 31331
rect 25881 31297 25915 31331
rect 26157 31297 26191 31331
rect 28089 31297 28123 31331
rect 28181 31297 28215 31331
rect 28457 31297 28491 31331
rect 29377 31297 29411 31331
rect 30297 31297 30331 31331
rect 30389 31297 30423 31331
rect 30573 31297 30607 31331
rect 30665 31297 30699 31331
rect 32321 31297 32355 31331
rect 32597 31297 32631 31331
rect 16681 31229 16715 31263
rect 19349 31229 19383 31263
rect 21281 31229 21315 31263
rect 27445 31229 27479 31263
rect 19257 31161 19291 31195
rect 21097 31161 21131 31195
rect 25421 31161 25455 31195
rect 21189 31093 21223 31127
rect 22753 31093 22787 31127
rect 28365 31093 28399 31127
rect 30113 31093 30147 31127
rect 32137 31093 32171 31127
rect 25513 30889 25547 30923
rect 26341 30889 26375 30923
rect 30205 30889 30239 30923
rect 31217 30889 31251 30923
rect 26525 30821 26559 30855
rect 27997 30821 28031 30855
rect 14565 30753 14599 30787
rect 28825 30753 28859 30787
rect 29009 30753 29043 30787
rect 30849 30753 30883 30787
rect 31769 30753 31803 30787
rect 32045 30753 32079 30787
rect 14105 30685 14139 30719
rect 17693 30685 17727 30719
rect 18061 30685 18095 30719
rect 22098 30685 22132 30719
rect 24409 30685 24443 30719
rect 25421 30685 25455 30719
rect 26065 30685 26099 30719
rect 26249 30685 26283 30719
rect 26341 30685 26375 30719
rect 28733 30685 28767 30719
rect 30021 30685 30055 30719
rect 30297 30685 30331 30719
rect 30941 30685 30975 30719
rect 14289 30617 14323 30651
rect 17877 30617 17911 30651
rect 17969 30617 18003 30651
rect 21281 30617 21315 30651
rect 21465 30617 21499 30651
rect 22385 30617 22419 30651
rect 24501 30617 24535 30651
rect 27813 30617 27847 30651
rect 18245 30549 18279 30583
rect 21649 30549 21683 30583
rect 23857 30549 23891 30583
rect 29009 30549 29043 30583
rect 29837 30549 29871 30583
rect 33517 30549 33551 30583
rect 25697 30345 25731 30379
rect 13737 30277 13771 30311
rect 16129 30277 16163 30311
rect 22017 30277 22051 30311
rect 29561 30277 29595 30311
rect 32505 30277 32539 30311
rect 13645 30209 13679 30243
rect 18245 30209 18279 30243
rect 18429 30209 18463 30243
rect 18521 30209 18555 30243
rect 22201 30209 22235 30243
rect 22661 30209 22695 30243
rect 22845 30209 22879 30243
rect 23029 30209 23063 30243
rect 24593 30209 24627 30243
rect 25513 30209 25547 30243
rect 26985 30209 27019 30243
rect 27169 30209 27203 30243
rect 28365 30209 28399 30243
rect 28549 30209 28583 30243
rect 29193 30209 29227 30243
rect 29377 30209 29411 30243
rect 30021 30209 30055 30243
rect 30205 30209 30239 30243
rect 32413 30209 32447 30243
rect 14289 30141 14323 30175
rect 14473 30141 14507 30175
rect 23121 30141 23155 30175
rect 28733 30073 28767 30107
rect 18061 30005 18095 30039
rect 24685 30005 24719 30039
rect 26985 30005 27019 30039
rect 27353 30005 27387 30039
rect 30205 30005 30239 30039
rect 30389 30005 30423 30039
rect 14657 29801 14691 29835
rect 18429 29801 18463 29835
rect 22477 29801 22511 29835
rect 26157 29801 26191 29835
rect 26801 29801 26835 29835
rect 29561 29801 29595 29835
rect 32229 29801 32263 29835
rect 22661 29733 22695 29767
rect 18245 29665 18279 29699
rect 20821 29665 20855 29699
rect 23397 29665 23431 29699
rect 24409 29665 24443 29699
rect 30481 29665 30515 29699
rect 30757 29665 30791 29699
rect 14565 29597 14599 29631
rect 18153 29597 18187 29631
rect 20637 29597 20671 29631
rect 20913 29597 20947 29631
rect 22109 29597 22143 29631
rect 22477 29597 22511 29631
rect 23121 29597 23155 29631
rect 23305 29597 23339 29631
rect 23489 29597 23523 29631
rect 23673 29597 23707 29631
rect 26709 29597 26743 29631
rect 27629 29597 27663 29631
rect 27813 29597 27847 29631
rect 28273 29597 28307 29631
rect 28457 29597 28491 29631
rect 29837 29597 29871 29631
rect 47317 29597 47351 29631
rect 47593 29597 47627 29631
rect 23857 29529 23891 29563
rect 24685 29529 24719 29563
rect 29561 29529 29595 29563
rect 29745 29529 29779 29563
rect 20453 29461 20487 29495
rect 27721 29461 27755 29495
rect 28641 29461 28675 29495
rect 23489 29257 23523 29291
rect 24593 29257 24627 29291
rect 30481 29257 30515 29291
rect 32229 29257 32263 29291
rect 13093 29121 13127 29155
rect 13737 29121 13771 29155
rect 13921 29121 13955 29155
rect 20177 29119 20211 29153
rect 20349 29119 20383 29153
rect 20453 29121 20487 29155
rect 20729 29121 20763 29155
rect 22293 29121 22327 29155
rect 22477 29121 22511 29155
rect 23121 29121 23155 29155
rect 23305 29121 23339 29155
rect 24501 29121 24535 29155
rect 25789 29121 25823 29155
rect 27077 29121 27111 29155
rect 27905 29121 27939 29155
rect 28181 29121 28215 29155
rect 28273 29121 28307 29155
rect 29193 29121 29227 29155
rect 29377 29121 29411 29155
rect 29561 29121 29595 29155
rect 29745 29121 29779 29155
rect 30389 29121 30423 29155
rect 32137 29121 32171 29155
rect 16681 29053 16715 29087
rect 16865 29053 16899 29087
rect 17141 29053 17175 29087
rect 20545 29053 20579 29087
rect 27169 29053 27203 29087
rect 27997 29053 28031 29087
rect 29469 29053 29503 29087
rect 13185 28985 13219 29019
rect 25973 28985 26007 29019
rect 27445 28985 27479 29019
rect 28089 28985 28123 29019
rect 29929 28985 29963 29019
rect 13829 28917 13863 28951
rect 20913 28917 20947 28951
rect 22293 28917 22327 28951
rect 22661 28917 22695 28951
rect 27261 28917 27295 28951
rect 15853 28713 15887 28747
rect 18705 28713 18739 28747
rect 21005 28713 21039 28747
rect 21557 28713 21591 28747
rect 22017 28713 22051 28747
rect 22477 28713 22511 28747
rect 26893 28713 26927 28747
rect 32321 28713 32355 28747
rect 9781 28577 9815 28611
rect 13277 28577 13311 28611
rect 14105 28577 14139 28611
rect 16957 28577 16991 28611
rect 19533 28577 19567 28611
rect 21741 28577 21775 28611
rect 28273 28577 28307 28611
rect 30849 28577 30883 28611
rect 46489 28577 46523 28611
rect 47685 28577 47719 28611
rect 9321 28509 9355 28543
rect 12081 28509 12115 28543
rect 12265 28509 12299 28543
rect 13185 28509 13219 28543
rect 19257 28509 19291 28543
rect 21465 28509 21499 28543
rect 22477 28509 22511 28543
rect 22661 28509 22695 28543
rect 27905 28509 27939 28543
rect 28089 28509 28123 28543
rect 28181 28509 28215 28543
rect 28457 28509 28491 28543
rect 29653 28509 29687 28543
rect 30573 28509 30607 28543
rect 46305 28509 46339 28543
rect 9505 28441 9539 28475
rect 14381 28441 14415 28475
rect 17233 28441 17267 28475
rect 26801 28441 26835 28475
rect 29837 28441 29871 28475
rect 12173 28373 12207 28407
rect 13553 28373 13587 28407
rect 22845 28373 22879 28407
rect 28641 28373 28675 28407
rect 10057 28169 10091 28203
rect 14749 28169 14783 28203
rect 16037 28169 16071 28203
rect 19073 28169 19107 28203
rect 19993 28169 20027 28203
rect 22845 28169 22879 28203
rect 24057 28169 24091 28203
rect 30205 28169 30239 28203
rect 32229 28169 32263 28203
rect 11805 28101 11839 28135
rect 13921 28101 13955 28135
rect 21005 28101 21039 28135
rect 23857 28101 23891 28135
rect 25513 28101 25547 28135
rect 25881 28101 25915 28135
rect 28733 28101 28767 28135
rect 9965 28033 9999 28067
rect 10885 28033 10919 28067
rect 13829 28033 13863 28067
rect 14657 28033 14691 28067
rect 15945 28033 15979 28067
rect 18981 28033 19015 28067
rect 19901 28033 19935 28067
rect 20821 28033 20855 28067
rect 22661 28033 22695 28067
rect 26985 28033 27019 28067
rect 27261 28033 27295 28067
rect 28457 28033 28491 28067
rect 32137 28033 32171 28067
rect 47593 28033 47627 28067
rect 10977 27965 11011 27999
rect 11529 27965 11563 27999
rect 16681 27965 16715 27999
rect 16865 27965 16899 27999
rect 17141 27965 17175 27999
rect 13277 27829 13311 27863
rect 21189 27829 21223 27863
rect 24041 27829 24075 27863
rect 24225 27829 24259 27863
rect 27077 27829 27111 27863
rect 27537 27829 27571 27863
rect 47041 27829 47075 27863
rect 47685 27829 47719 27863
rect 12173 27625 12207 27659
rect 17049 27625 17083 27659
rect 22293 27625 22327 27659
rect 26525 27625 26559 27659
rect 13277 27557 13311 27591
rect 14105 27557 14139 27591
rect 23121 27557 23155 27591
rect 28917 27557 28951 27591
rect 30849 27557 30883 27591
rect 11989 27489 12023 27523
rect 15577 27489 15611 27523
rect 22201 27489 22235 27523
rect 26893 27489 26927 27523
rect 46305 27489 46339 27523
rect 48145 27489 48179 27523
rect 9413 27421 9447 27455
rect 11805 27421 11839 27455
rect 12173 27421 12207 27455
rect 12725 27421 12759 27455
rect 12909 27421 12943 27455
rect 14289 27421 14323 27455
rect 14381 27421 14415 27455
rect 15761 27421 15795 27455
rect 16957 27421 16991 27455
rect 22293 27421 22327 27455
rect 22937 27421 22971 27455
rect 23673 27421 23707 27455
rect 24501 27421 24535 27455
rect 26709 27421 26743 27455
rect 26985 27421 27019 27455
rect 28733 27421 28767 27455
rect 29561 27421 29595 27455
rect 29749 27415 29783 27449
rect 29840 27421 29874 27455
rect 29929 27421 29963 27455
rect 30067 27421 30101 27455
rect 30757 27421 30791 27455
rect 13093 27353 13127 27387
rect 14473 27353 14507 27387
rect 22017 27353 22051 27387
rect 46489 27353 46523 27387
rect 9413 27285 9447 27319
rect 11897 27285 11931 27319
rect 13001 27285 13035 27319
rect 14657 27285 14691 27319
rect 15945 27285 15979 27319
rect 22477 27285 22511 27319
rect 23765 27285 23799 27319
rect 24685 27285 24719 27319
rect 30297 27285 30331 27319
rect 24593 27081 24627 27115
rect 31585 27081 31619 27115
rect 13645 27013 13679 27047
rect 23673 27013 23707 27047
rect 27997 27013 28031 27047
rect 28181 27013 28215 27047
rect 30113 27013 30147 27047
rect 32229 27013 32263 27047
rect 9137 26945 9171 26979
rect 12817 26945 12851 26979
rect 13001 26945 13035 26979
rect 13553 26945 13587 26979
rect 13737 26945 13771 26979
rect 15393 26945 15427 26979
rect 16681 26945 16715 26979
rect 16865 26945 16899 26979
rect 22201 26945 22235 26979
rect 22293 26945 22327 26979
rect 22477 26945 22511 26979
rect 22661 26945 22695 26979
rect 23489 26945 23523 26979
rect 23765 26945 23799 26979
rect 24685 26945 24719 26979
rect 26065 26945 26099 26979
rect 26985 26945 27019 26979
rect 27261 26945 27295 26979
rect 29837 26945 29871 26979
rect 32137 26945 32171 26979
rect 9413 26877 9447 26911
rect 13093 26877 13127 26911
rect 24777 26877 24811 26911
rect 26157 26877 26191 26911
rect 27169 26877 27203 26911
rect 15577 26809 15611 26843
rect 22385 26809 22419 26843
rect 24225 26809 24259 26843
rect 27445 26809 27479 26843
rect 10885 26741 10919 26775
rect 12633 26741 12667 26775
rect 16681 26741 16715 26775
rect 21925 26741 21959 26775
rect 23305 26741 23339 26775
rect 26341 26741 26375 26775
rect 26985 26741 27019 26775
rect 10241 26537 10275 26571
rect 13553 26537 13587 26571
rect 15393 26537 15427 26571
rect 22109 26537 22143 26571
rect 24961 26537 24995 26571
rect 27629 26537 27663 26571
rect 28641 26537 28675 26571
rect 20545 26469 20579 26503
rect 9965 26401 9999 26435
rect 12081 26401 12115 26435
rect 16405 26401 16439 26435
rect 21189 26401 21223 26435
rect 24777 26401 24811 26435
rect 32321 26401 32355 26435
rect 46305 26401 46339 26435
rect 47777 26401 47811 26435
rect 9873 26333 9907 26367
rect 11805 26333 11839 26367
rect 14105 26333 14139 26367
rect 15393 26333 15427 26367
rect 15669 26333 15703 26367
rect 16129 26333 16163 26367
rect 18337 26333 18371 26367
rect 19901 26333 19935 26367
rect 20913 26333 20947 26367
rect 24409 26333 24443 26367
rect 24567 26333 24601 26367
rect 25697 26333 25731 26367
rect 26065 26333 26099 26367
rect 27261 26333 27295 26367
rect 27537 26333 27571 26367
rect 28273 26333 28307 26367
rect 28457 26333 28491 26367
rect 31309 26333 31343 26367
rect 32045 26333 32079 26367
rect 14197 26265 14231 26299
rect 15577 26265 15611 26299
rect 21741 26265 21775 26299
rect 21925 26265 21959 26299
rect 25881 26265 25915 26299
rect 25973 26265 26007 26299
rect 31401 26265 31435 26299
rect 46489 26265 46523 26299
rect 17877 26197 17911 26231
rect 18429 26197 18463 26231
rect 19717 26197 19751 26231
rect 21005 26197 21039 26231
rect 26249 26197 26283 26231
rect 27813 26197 27847 26231
rect 10333 25993 10367 26027
rect 12725 25993 12759 26027
rect 15761 25993 15795 26027
rect 17049 25993 17083 26027
rect 17233 25993 17267 26027
rect 16681 25925 16715 25959
rect 18521 25925 18555 25959
rect 20177 25925 20211 25959
rect 26985 25925 27019 25959
rect 27353 25925 27387 25959
rect 32321 25925 32355 25959
rect 33977 25925 34011 25959
rect 10241 25857 10275 25891
rect 12633 25857 12667 25891
rect 15577 25857 15611 25891
rect 16865 25857 16899 25891
rect 16957 25857 16991 25891
rect 21005 25857 21039 25891
rect 21833 25857 21867 25891
rect 22293 25857 22327 25891
rect 27169 25857 27203 25891
rect 27997 25857 28031 25891
rect 28181 25857 28215 25891
rect 28549 25857 28583 25891
rect 30941 25857 30975 25891
rect 46581 25857 46615 25891
rect 15393 25789 15427 25823
rect 18337 25789 18371 25823
rect 21281 25789 21315 25823
rect 22201 25789 22235 25823
rect 28273 25789 28307 25823
rect 28365 25789 28399 25823
rect 31309 25789 31343 25823
rect 32137 25789 32171 25823
rect 21097 25721 21131 25755
rect 47777 25721 47811 25755
rect 21189 25653 21223 25687
rect 22293 25653 22327 25687
rect 22477 25653 22511 25687
rect 28733 25653 28767 25687
rect 46673 25653 46707 25687
rect 16681 25449 16715 25483
rect 17601 25449 17635 25483
rect 21465 25449 21499 25483
rect 29009 25449 29043 25483
rect 21741 25381 21775 25415
rect 21833 25381 21867 25415
rect 22477 25381 22511 25415
rect 12725 25313 12759 25347
rect 21005 25313 21039 25347
rect 46489 25313 46523 25347
rect 48145 25313 48179 25347
rect 1409 25245 1443 25279
rect 9873 25245 9907 25279
rect 12633 25245 12667 25279
rect 15761 25245 15795 25279
rect 16037 25245 16071 25279
rect 16589 25245 16623 25279
rect 17509 25245 17543 25279
rect 18521 25245 18555 25279
rect 19257 25245 19291 25279
rect 21649 25245 21683 25279
rect 21914 25245 21948 25279
rect 22753 25245 22787 25279
rect 25329 25245 25363 25279
rect 25605 25245 25639 25279
rect 27261 25245 27295 25279
rect 31493 25245 31527 25279
rect 32137 25245 32171 25279
rect 45661 25245 45695 25279
rect 46305 25245 46339 25279
rect 1685 25177 1719 25211
rect 10149 25177 10183 25211
rect 19533 25177 19567 25211
rect 22477 25177 22511 25211
rect 25513 25177 25547 25211
rect 27537 25177 27571 25211
rect 31309 25177 31343 25211
rect 32781 25177 32815 25211
rect 11621 25109 11655 25143
rect 13001 25109 13035 25143
rect 15577 25109 15611 25143
rect 15945 25109 15979 25143
rect 18613 25109 18647 25143
rect 22661 25109 22695 25143
rect 25145 25109 25179 25143
rect 45753 25109 45787 25143
rect 9873 24905 9907 24939
rect 10517 24905 10551 24939
rect 14565 24905 14599 24939
rect 15761 24905 15795 24939
rect 18429 24905 18463 24939
rect 21281 24905 21315 24939
rect 22753 24905 22787 24939
rect 25237 24905 25271 24939
rect 13093 24837 13127 24871
rect 15485 24837 15519 24871
rect 15669 24837 15703 24871
rect 9781 24769 9815 24803
rect 10425 24769 10459 24803
rect 10609 24769 10643 24803
rect 11529 24769 11563 24803
rect 15853 24769 15887 24803
rect 16037 24769 16071 24803
rect 22569 24769 22603 24803
rect 22845 24769 22879 24803
rect 26157 24769 26191 24803
rect 27997 24769 28031 24803
rect 28089 24769 28123 24803
rect 32137 24769 32171 24803
rect 11621 24701 11655 24735
rect 12817 24701 12851 24735
rect 16681 24701 16715 24735
rect 16957 24701 16991 24735
rect 19533 24701 19567 24735
rect 19809 24701 19843 24735
rect 22385 24701 22419 24735
rect 23489 24701 23523 24735
rect 23765 24701 23799 24735
rect 29377 24701 29411 24735
rect 29561 24701 29595 24735
rect 29837 24701 29871 24735
rect 32321 24701 32355 24735
rect 45201 24701 45235 24735
rect 45385 24701 45419 24735
rect 46857 24701 46891 24735
rect 26249 24565 26283 24599
rect 47777 24565 47811 24599
rect 10333 24361 10367 24395
rect 24593 24361 24627 24395
rect 13461 24293 13495 24327
rect 14105 24293 14139 24327
rect 15301 24293 15335 24327
rect 16497 24293 16531 24327
rect 17785 24293 17819 24327
rect 20453 24293 20487 24327
rect 26893 24293 26927 24327
rect 29653 24293 29687 24327
rect 12541 24225 12575 24259
rect 16313 24225 16347 24259
rect 25145 24225 25179 24259
rect 46029 24225 46063 24259
rect 47317 24225 47351 24259
rect 9137 24157 9171 24191
rect 9689 24157 9723 24191
rect 10609 24157 10643 24191
rect 11069 24157 11103 24191
rect 13369 24157 13403 24191
rect 14105 24157 14139 24191
rect 15669 24157 15703 24191
rect 16773 24157 16807 24191
rect 17693 24157 17727 24191
rect 19441 24157 19475 24191
rect 20361 24157 20395 24191
rect 24501 24157 24535 24191
rect 29561 24157 29595 24191
rect 45845 24157 45879 24191
rect 10333 24089 10367 24123
rect 11253 24089 11287 24123
rect 15577 24089 15611 24123
rect 25421 24089 25455 24123
rect 9137 24021 9171 24055
rect 9781 24021 9815 24055
rect 10517 24021 10551 24055
rect 15485 24021 15519 24055
rect 15853 24021 15887 24055
rect 16681 24021 16715 24055
rect 1961 23817 1995 23851
rect 47685 23817 47719 23851
rect 12173 23749 12207 23783
rect 12389 23749 12423 23783
rect 25973 23749 26007 23783
rect 27169 23749 27203 23783
rect 28825 23749 28859 23783
rect 1869 23681 1903 23715
rect 8217 23681 8251 23715
rect 13277 23681 13311 23715
rect 15301 23681 15335 23715
rect 16681 23681 16715 23715
rect 18705 23681 18739 23715
rect 19349 23681 19383 23715
rect 20085 23681 20119 23715
rect 21833 23681 21867 23715
rect 22937 23681 22971 23715
rect 23581 23681 23615 23715
rect 23765 23681 23799 23715
rect 25881 23681 25915 23715
rect 30389 23681 30423 23715
rect 31217 23681 31251 23715
rect 45845 23681 45879 23715
rect 46213 23681 46247 23715
rect 47593 23681 47627 23715
rect 8493 23613 8527 23647
rect 9965 23613 9999 23647
rect 15577 23613 15611 23647
rect 26985 23613 27019 23647
rect 31125 23613 31159 23647
rect 32229 23613 32263 23647
rect 32413 23613 32447 23647
rect 33149 23613 33183 23647
rect 44465 23613 44499 23647
rect 44741 23613 44775 23647
rect 46765 23613 46799 23647
rect 12541 23545 12575 23579
rect 16681 23545 16715 23579
rect 19533 23545 19567 23579
rect 22017 23545 22051 23579
rect 30481 23545 30515 23579
rect 12357 23477 12391 23511
rect 13461 23477 13495 23511
rect 18797 23477 18831 23511
rect 20177 23477 20211 23511
rect 23029 23477 23063 23511
rect 23581 23477 23615 23511
rect 31585 23477 31619 23511
rect 9045 23273 9079 23307
rect 9597 23273 9631 23307
rect 10333 23273 10367 23307
rect 10517 23273 10551 23307
rect 11621 23273 11655 23307
rect 14565 23273 14599 23307
rect 18245 23273 18279 23307
rect 14749 23205 14783 23239
rect 33517 23205 33551 23239
rect 13369 23137 13403 23171
rect 15485 23137 15519 23171
rect 15761 23137 15795 23171
rect 19257 23137 19291 23171
rect 22293 23137 22327 23171
rect 23765 23137 23799 23171
rect 31309 23137 31343 23171
rect 31769 23137 31803 23171
rect 32045 23137 32079 23171
rect 41797 23137 41831 23171
rect 46305 23137 46339 23171
rect 46765 23137 46799 23171
rect 9226 23069 9260 23103
rect 9689 23069 9723 23103
rect 11529 23069 11563 23103
rect 15393 23069 15427 23103
rect 18061 23069 18095 23103
rect 22017 23069 22051 23103
rect 29561 23069 29595 23103
rect 33977 23069 34011 23103
rect 39957 23069 39991 23103
rect 45845 23069 45879 23103
rect 10149 23001 10183 23035
rect 13093 23001 13127 23035
rect 14381 23001 14415 23035
rect 19441 23001 19475 23035
rect 21097 23001 21131 23035
rect 29837 23001 29871 23035
rect 40141 23001 40175 23035
rect 46489 23001 46523 23035
rect 9229 22933 9263 22967
rect 10349 22933 10383 22967
rect 14591 22933 14625 22967
rect 34069 22933 34103 22967
rect 45661 22933 45695 22967
rect 10609 22729 10643 22763
rect 12725 22729 12759 22763
rect 22477 22729 22511 22763
rect 24133 22729 24167 22763
rect 28549 22729 28583 22763
rect 30757 22729 30791 22763
rect 30941 22729 30975 22763
rect 31493 22729 31527 22763
rect 32229 22729 32263 22763
rect 33057 22729 33091 22763
rect 40141 22729 40175 22763
rect 45201 22729 45235 22763
rect 47685 22729 47719 22763
rect 9321 22661 9355 22695
rect 10241 22661 10275 22695
rect 10457 22661 10491 22695
rect 14381 22661 14415 22695
rect 17693 22661 17727 22695
rect 22293 22661 22327 22695
rect 23029 22661 23063 22695
rect 23245 22661 23279 22695
rect 41521 22661 41555 22695
rect 11897 22593 11931 22627
rect 12541 22593 12575 22627
rect 13369 22593 13403 22627
rect 16773 22593 16807 22627
rect 18429 22593 18463 22627
rect 18797 22593 18831 22627
rect 19625 22593 19659 22627
rect 20177 22593 20211 22627
rect 20913 22593 20947 22627
rect 22569 22593 22603 22627
rect 23857 22593 23891 22627
rect 24041 22593 24075 22627
rect 24225 22593 24259 22627
rect 25053 22593 25087 22627
rect 25881 22593 25915 22627
rect 28549 22593 28583 22627
rect 29285 22593 29319 22627
rect 30389 22593 30423 22627
rect 30573 22593 30607 22627
rect 30665 22593 30699 22627
rect 31401 22593 31435 22627
rect 32137 22593 32171 22627
rect 32965 22593 32999 22627
rect 40049 22593 40083 22627
rect 42441 22593 42475 22627
rect 45017 22593 45051 22627
rect 45201 22593 45235 22627
rect 46397 22593 46431 22627
rect 47593 22593 47627 22627
rect 13553 22525 13587 22559
rect 14105 22525 14139 22559
rect 20821 22525 20855 22559
rect 24409 22525 24443 22559
rect 24869 22525 24903 22559
rect 29377 22525 29411 22559
rect 29653 22525 29687 22559
rect 33701 22525 33735 22559
rect 33885 22525 33919 22559
rect 35541 22525 35575 22559
rect 42717 22525 42751 22559
rect 45661 22525 45695 22559
rect 46765 22525 46799 22559
rect 9597 22457 9631 22491
rect 17877 22457 17911 22491
rect 23397 22457 23431 22491
rect 45937 22457 45971 22491
rect 9781 22389 9815 22423
rect 10425 22389 10459 22423
rect 11989 22389 12023 22423
rect 15853 22389 15887 22423
rect 16865 22389 16899 22423
rect 21281 22389 21315 22423
rect 22293 22389 22327 22423
rect 23213 22389 23247 22423
rect 25237 22389 25271 22423
rect 25697 22389 25731 22423
rect 41613 22389 41647 22423
rect 9505 22185 9539 22219
rect 14105 22185 14139 22219
rect 20256 22185 20290 22219
rect 22293 22185 22327 22219
rect 26433 22185 26467 22219
rect 30205 22185 30239 22219
rect 30389 22185 30423 22219
rect 41429 22185 41463 22219
rect 45845 22185 45879 22219
rect 11897 22049 11931 22083
rect 12173 22049 12207 22083
rect 14933 22049 14967 22083
rect 17969 22049 18003 22083
rect 21741 22049 21775 22083
rect 24685 22049 24719 22083
rect 27169 22049 27203 22083
rect 46489 22049 46523 22083
rect 47777 22049 47811 22083
rect 8401 21981 8435 22015
rect 9689 21981 9723 22015
rect 9975 21959 10009 21993
rect 10609 21981 10643 22015
rect 11713 21981 11747 22015
rect 14105 21981 14139 22015
rect 14841 21981 14875 22015
rect 16773 21981 16807 22015
rect 19257 21981 19291 22015
rect 19993 21981 20027 22015
rect 22477 21981 22511 22015
rect 23581 21981 23615 22015
rect 23857 21981 23891 22015
rect 26893 21981 26927 22015
rect 31125 21981 31159 22015
rect 41245 21981 41279 22015
rect 43913 21981 43947 22015
rect 46305 21981 46339 22015
rect 10793 21913 10827 21947
rect 16957 21913 16991 21947
rect 24961 21913 24995 21947
rect 30021 21913 30055 21947
rect 30849 21913 30883 21947
rect 45477 21913 45511 21947
rect 45661 21913 45695 21947
rect 8217 21845 8251 21879
rect 9873 21845 9907 21879
rect 19441 21845 19475 21879
rect 23679 21845 23713 21879
rect 23765 21845 23799 21879
rect 28641 21845 28675 21879
rect 30221 21845 30255 21879
rect 30947 21845 30981 21879
rect 31033 21845 31067 21879
rect 44005 21845 44039 21879
rect 16037 21641 16071 21675
rect 21005 21641 21039 21675
rect 24869 21641 24903 21675
rect 26249 21641 26283 21675
rect 28273 21641 28307 21675
rect 46213 21641 46247 21675
rect 9413 21573 9447 21607
rect 16865 21573 16899 21607
rect 44005 21573 44039 21607
rect 47961 21573 47995 21607
rect 11897 21505 11931 21539
rect 13185 21505 13219 21539
rect 15301 21505 15335 21539
rect 15945 21505 15979 21539
rect 19993 21505 20027 21539
rect 20821 21505 20855 21539
rect 22201 21505 22235 21539
rect 23213 21505 23247 21539
rect 23765 21505 23799 21539
rect 24777 21505 24811 21539
rect 24961 21505 24995 21539
rect 25421 21505 25455 21539
rect 26157 21505 26191 21539
rect 27353 21505 27387 21539
rect 28181 21505 28215 21539
rect 30113 21505 30147 21539
rect 30297 21505 30331 21539
rect 31217 21505 31251 21539
rect 46121 21505 46155 21539
rect 46305 21505 46339 21539
rect 46857 21505 46891 21539
rect 9137 21437 9171 21471
rect 10885 21437 10919 21471
rect 16681 21437 16715 21471
rect 18337 21437 18371 21471
rect 22293 21437 22327 21471
rect 27261 21437 27295 21471
rect 27721 21437 27755 21471
rect 43821 21437 43855 21471
rect 45385 21437 45419 21471
rect 23029 21369 23063 21403
rect 48145 21369 48179 21403
rect 12081 21301 12115 21335
rect 13369 21301 13403 21335
rect 15393 21301 15427 21335
rect 20269 21301 20303 21335
rect 22569 21301 22603 21335
rect 23857 21301 23891 21335
rect 25605 21301 25639 21335
rect 30113 21301 30147 21335
rect 31309 21301 31343 21335
rect 46949 21301 46983 21335
rect 9229 21097 9263 21131
rect 10241 21097 10275 21131
rect 18153 21097 18187 21131
rect 20269 21097 20303 21131
rect 21097 21097 21131 21131
rect 26065 21029 26099 21063
rect 11989 20961 12023 20995
rect 15853 20961 15887 20995
rect 17509 20961 17543 20995
rect 22109 20961 22143 20995
rect 22385 20961 22419 20995
rect 30481 20961 30515 20995
rect 46489 20961 46523 20995
rect 48145 20961 48179 20995
rect 9413 20893 9447 20927
rect 10149 20893 10183 20927
rect 10885 20893 10919 20927
rect 11529 20893 11563 20927
rect 14565 20893 14599 20927
rect 15669 20893 15703 20927
rect 18061 20893 18095 20927
rect 19257 20893 19291 20927
rect 20453 20893 20487 20927
rect 21005 20893 21039 20927
rect 25973 20893 26007 20927
rect 30205 20893 30239 20927
rect 33333 20893 33367 20927
rect 43729 20893 43763 20927
rect 46305 20893 46339 20927
rect 10977 20825 11011 20859
rect 11713 20825 11747 20859
rect 14657 20757 14691 20791
rect 19349 20757 19383 20791
rect 23857 20757 23891 20791
rect 31953 20757 31987 20791
rect 33425 20757 33459 20791
rect 43821 20757 43855 20791
rect 15393 20553 15427 20587
rect 30205 20553 30239 20587
rect 33333 20485 33367 20519
rect 43821 20485 43855 20519
rect 9321 20417 9355 20451
rect 9965 20417 9999 20451
rect 12357 20417 12391 20451
rect 12909 20417 12943 20451
rect 17049 20417 17083 20451
rect 21833 20417 21867 20451
rect 24869 20417 24903 20451
rect 26249 20417 26283 20451
rect 27445 20417 27479 20451
rect 28089 20417 28123 20451
rect 30021 20417 30055 20451
rect 33149 20417 33183 20451
rect 46397 20417 46431 20451
rect 46857 20417 46891 20451
rect 47777 20417 47811 20451
rect 12449 20349 12483 20383
rect 13645 20349 13679 20383
rect 13921 20349 13955 20383
rect 17693 20349 17727 20383
rect 18337 20349 18371 20383
rect 18613 20349 18647 20383
rect 34989 20349 35023 20383
rect 43637 20349 43671 20383
rect 45477 20349 45511 20383
rect 46029 20349 46063 20383
rect 25053 20281 25087 20315
rect 28273 20281 28307 20315
rect 46765 20281 46799 20315
rect 9137 20213 9171 20247
rect 10057 20213 10091 20247
rect 13093 20213 13127 20247
rect 20085 20213 20119 20247
rect 21925 20213 21959 20247
rect 26341 20213 26375 20247
rect 10701 20009 10735 20043
rect 13553 20009 13587 20043
rect 14657 20009 14691 20043
rect 26985 20009 27019 20043
rect 47777 20009 47811 20043
rect 14105 19941 14139 19975
rect 27721 19941 27755 19975
rect 45477 19941 45511 19975
rect 8953 19873 8987 19907
rect 13277 19873 13311 19907
rect 17969 19873 18003 19907
rect 21925 19873 21959 19907
rect 22201 19873 22235 19907
rect 24501 19873 24535 19907
rect 25513 19873 25547 19907
rect 44373 19873 44407 19907
rect 45201 19873 45235 19907
rect 45661 19873 45695 19907
rect 46305 19873 46339 19907
rect 47133 19873 47167 19907
rect 2053 19805 2087 19839
rect 11437 19805 11471 19839
rect 11713 19805 11747 19839
rect 11897 19805 11931 19839
rect 13185 19805 13219 19839
rect 14289 19805 14323 19839
rect 16405 19805 16439 19839
rect 17233 19805 17267 19839
rect 19441 19805 19475 19839
rect 20821 19805 20855 19839
rect 21741 19805 21775 19839
rect 25973 19805 26007 19839
rect 26157 19805 26191 19839
rect 26617 19805 26651 19839
rect 26801 19805 26835 19839
rect 27445 19805 27479 19839
rect 27629 19805 27663 19839
rect 28825 19805 28859 19839
rect 29561 19805 29595 19839
rect 44281 19805 44315 19839
rect 44465 19805 44499 19839
rect 46397 19805 46431 19839
rect 47685 19805 47719 19839
rect 47869 19805 47903 19839
rect 9229 19737 9263 19771
rect 14473 19737 14507 19771
rect 24593 19737 24627 19771
rect 28917 19737 28951 19771
rect 29745 19737 29779 19771
rect 31401 19737 31435 19771
rect 11253 19669 11287 19703
rect 14381 19669 14415 19703
rect 16589 19669 16623 19703
rect 19441 19669 19475 19703
rect 21005 19669 21039 19703
rect 26157 19669 26191 19703
rect 13277 19465 13311 19499
rect 21925 19465 21959 19499
rect 27261 19465 27295 19499
rect 27353 19465 27387 19499
rect 44833 19465 44867 19499
rect 11805 19397 11839 19431
rect 13921 19397 13955 19431
rect 14289 19397 14323 19431
rect 17417 19397 17451 19431
rect 26341 19397 26375 19431
rect 27537 19397 27571 19431
rect 29561 19397 29595 19431
rect 39313 19397 39347 19431
rect 40233 19397 40267 19431
rect 1777 19329 1811 19363
rect 8861 19329 8895 19363
rect 10885 19329 10919 19363
rect 14105 19329 14139 19363
rect 14197 19329 14231 19363
rect 17141 19329 17175 19363
rect 18429 19329 18463 19363
rect 20729 19329 20763 19363
rect 20913 19329 20947 19363
rect 22109 19329 22143 19363
rect 26249 19329 26283 19363
rect 26433 19329 26467 19363
rect 27169 19329 27203 19363
rect 45201 19329 45235 19363
rect 45293 19329 45327 19363
rect 47593 19329 47627 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 8953 19261 8987 19295
rect 9229 19261 9263 19295
rect 10977 19261 11011 19295
rect 11529 19261 11563 19295
rect 14473 19261 14507 19295
rect 18705 19261 18739 19295
rect 29469 19261 29503 19295
rect 30481 19261 30515 19295
rect 39221 19261 39255 19295
rect 45477 19261 45511 19295
rect 46213 19261 46247 19295
rect 47041 19261 47075 19295
rect 26985 19193 27019 19227
rect 20177 19125 20211 19159
rect 20821 19125 20855 19159
rect 47685 19125 47719 19159
rect 2237 18921 2271 18955
rect 12633 18921 12667 18955
rect 14289 18921 14323 18955
rect 14473 18921 14507 18955
rect 17877 18921 17911 18955
rect 18521 18921 18555 18955
rect 26433 18921 26467 18955
rect 9413 18785 9447 18819
rect 19257 18785 19291 18819
rect 20729 18785 20763 18819
rect 21005 18785 21039 18819
rect 26249 18785 26283 18819
rect 46489 18785 46523 18819
rect 48145 18785 48179 18819
rect 2145 18717 2179 18751
rect 8217 18717 8251 18751
rect 8953 18717 8987 18751
rect 12541 18717 12575 18751
rect 13185 18717 13219 18751
rect 15393 18717 15427 18751
rect 15485 18717 15519 18751
rect 17509 18717 17543 18751
rect 18705 18717 18739 18751
rect 19533 18717 19567 18751
rect 20821 18717 20855 18751
rect 20913 18717 20947 18751
rect 22293 18717 22327 18751
rect 22845 18717 22879 18751
rect 23673 18717 23707 18751
rect 24409 18717 24443 18751
rect 25973 18717 26007 18751
rect 26065 18717 26099 18751
rect 26341 18717 26375 18751
rect 26893 18717 26927 18751
rect 27077 18717 27111 18751
rect 45845 18717 45879 18751
rect 46305 18717 46339 18751
rect 8309 18649 8343 18683
rect 9137 18649 9171 18683
rect 14105 18649 14139 18683
rect 17325 18649 17359 18683
rect 17601 18649 17635 18683
rect 27261 18649 27295 18683
rect 28089 18649 28123 18683
rect 28457 18649 28491 18683
rect 13277 18581 13311 18615
rect 14315 18581 14349 18615
rect 15669 18581 15703 18615
rect 17693 18581 17727 18615
rect 20545 18581 20579 18615
rect 22293 18581 22327 18615
rect 23029 18581 23063 18615
rect 23765 18581 23799 18615
rect 24501 18581 24535 18615
rect 1961 18377 1995 18411
rect 28181 18377 28215 18411
rect 46949 18377 46983 18411
rect 16037 18309 16071 18343
rect 16865 18309 16899 18343
rect 18981 18309 19015 18343
rect 19349 18309 19383 18343
rect 20085 18309 20119 18343
rect 26157 18309 26191 18343
rect 26985 18309 27019 18343
rect 27169 18309 27203 18343
rect 47961 18309 47995 18343
rect 1869 18241 1903 18275
rect 12909 18241 12943 18275
rect 15117 18241 15151 18275
rect 15301 18241 15335 18275
rect 15945 18241 15979 18275
rect 16681 18241 16715 18275
rect 19165 18241 19199 18275
rect 19257 18241 19291 18275
rect 19993 18241 20027 18275
rect 20913 18241 20947 18275
rect 22477 18241 22511 18275
rect 25421 18241 25455 18275
rect 25605 18241 25639 18275
rect 26065 18241 26099 18275
rect 26249 18241 26283 18275
rect 27353 18241 27387 18275
rect 27997 18241 28031 18275
rect 28641 18241 28675 18275
rect 46857 18241 46891 18275
rect 47041 18241 47075 18275
rect 47593 18241 47627 18275
rect 47777 18241 47811 18275
rect 13185 18173 13219 18207
rect 18521 18173 18555 18207
rect 20821 18173 20855 18207
rect 22753 18173 22787 18207
rect 24501 18173 24535 18207
rect 27813 18173 27847 18207
rect 15117 18105 15151 18139
rect 21281 18105 21315 18139
rect 25513 18105 25547 18139
rect 14657 18037 14691 18071
rect 19533 18037 19567 18071
rect 28733 18037 28767 18071
rect 14105 17833 14139 17867
rect 19717 17833 19751 17867
rect 21373 17833 21407 17867
rect 23765 17833 23799 17867
rect 26433 17833 26467 17867
rect 47501 17833 47535 17867
rect 19625 17765 19659 17799
rect 46765 17765 46799 17799
rect 11897 17697 11931 17731
rect 15393 17697 15427 17731
rect 18429 17697 18463 17731
rect 19257 17697 19291 17731
rect 21005 17697 21039 17731
rect 22017 17697 22051 17731
rect 11437 17629 11471 17663
rect 14105 17629 14139 17663
rect 14381 17629 14415 17663
rect 18245 17629 18279 17663
rect 20361 17629 20395 17663
rect 21189 17629 21223 17663
rect 27629 17629 27663 17663
rect 28089 17629 28123 17663
rect 46949 17629 46983 17663
rect 47409 17629 47443 17663
rect 47593 17629 47627 17663
rect 11621 17561 11655 17595
rect 15577 17561 15611 17595
rect 17233 17561 17267 17595
rect 17877 17561 17911 17595
rect 18061 17561 18095 17595
rect 20177 17561 20211 17595
rect 20545 17561 20579 17595
rect 22293 17561 22327 17595
rect 26065 17561 26099 17595
rect 26249 17561 26283 17595
rect 14289 17493 14323 17527
rect 18153 17493 18187 17527
rect 11713 17289 11747 17323
rect 14013 17289 14047 17323
rect 15209 17289 15243 17323
rect 18455 17289 18489 17323
rect 22017 17289 22051 17323
rect 8033 17221 8067 17255
rect 8769 17221 8803 17255
rect 18245 17221 18279 17255
rect 27905 17221 27939 17255
rect 7941 17153 7975 17187
rect 11621 17153 11655 17187
rect 13921 17153 13955 17187
rect 15117 17153 15151 17187
rect 15761 17153 15795 17187
rect 19809 17153 19843 17187
rect 21833 17153 21867 17187
rect 47593 17153 47627 17187
rect 8585 17085 8619 17119
rect 10425 17085 10459 17119
rect 27721 17085 27755 17119
rect 28181 17085 28215 17119
rect 18613 17017 18647 17051
rect 2053 16949 2087 16983
rect 15853 16949 15887 16983
rect 18429 16949 18463 16983
rect 19625 16949 19659 16983
rect 47041 16949 47075 16983
rect 47685 16949 47719 16983
rect 1409 16609 1443 16643
rect 1869 16609 1903 16643
rect 15761 16609 15795 16643
rect 19349 16609 19383 16643
rect 19809 16609 19843 16643
rect 46305 16609 46339 16643
rect 48145 16609 48179 16643
rect 15577 16541 15611 16575
rect 18429 16541 18463 16575
rect 19441 16541 19475 16575
rect 1593 16473 1627 16507
rect 17417 16473 17451 16507
rect 18153 16473 18187 16507
rect 20361 16473 20395 16507
rect 46489 16473 46523 16507
rect 18251 16405 18285 16439
rect 18337 16405 18371 16439
rect 20453 16405 20487 16439
rect 2145 16201 2179 16235
rect 15301 16201 15335 16235
rect 18981 16201 19015 16235
rect 21189 16201 21223 16235
rect 19717 16133 19751 16167
rect 2053 16065 2087 16099
rect 12725 16065 12759 16099
rect 19441 16065 19475 16099
rect 47593 16065 47627 16099
rect 12817 15997 12851 16031
rect 13553 15997 13587 16031
rect 13829 15997 13863 16031
rect 17233 15997 17267 16031
rect 17509 15997 17543 16031
rect 13093 15929 13127 15963
rect 47041 15861 47075 15895
rect 47685 15861 47719 15895
rect 14105 15657 14139 15691
rect 14933 15657 14967 15691
rect 19349 15657 19383 15691
rect 20637 15657 20671 15691
rect 16405 15521 16439 15555
rect 46305 15521 46339 15555
rect 46489 15521 46523 15555
rect 48145 15521 48179 15555
rect 2053 15453 2087 15487
rect 14289 15453 14323 15487
rect 14841 15453 14875 15487
rect 15761 15453 15795 15487
rect 19257 15453 19291 15487
rect 20545 15453 20579 15487
rect 15853 15385 15887 15419
rect 16589 15385 16623 15419
rect 18245 15385 18279 15419
rect 17417 15113 17451 15147
rect 18061 15113 18095 15147
rect 1777 14977 1811 15011
rect 14841 14977 14875 15011
rect 17417 14977 17451 15011
rect 17969 14977 18003 15011
rect 18153 14977 18187 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 14933 14773 14967 14807
rect 2237 14569 2271 14603
rect 17417 14569 17451 14603
rect 17601 14501 17635 14535
rect 2145 14365 2179 14399
rect 14289 14365 14323 14399
rect 15393 14365 15427 14399
rect 15669 14365 15703 14399
rect 15853 14365 15887 14399
rect 16313 14365 16347 14399
rect 18245 14365 18279 14399
rect 19257 14365 19291 14399
rect 17233 14297 17267 14331
rect 17449 14297 17483 14331
rect 14473 14229 14507 14263
rect 15209 14229 15243 14263
rect 16405 14229 16439 14263
rect 18245 14229 18279 14263
rect 19349 14229 19383 14263
rect 16037 14025 16071 14059
rect 17417 14025 17451 14059
rect 20821 14025 20855 14059
rect 17049 13957 17083 13991
rect 17265 13957 17299 13991
rect 19349 13957 19383 13991
rect 14289 13889 14323 13923
rect 18245 13889 18279 13923
rect 47593 13889 47627 13923
rect 18153 13821 18187 13855
rect 18613 13821 18647 13855
rect 19073 13821 19107 13855
rect 14552 13685 14586 13719
rect 17233 13685 17267 13719
rect 47685 13685 47719 13719
rect 19441 13481 19475 13515
rect 20177 13481 20211 13515
rect 15669 13345 15703 13379
rect 15853 13345 15887 13379
rect 16129 13345 16163 13379
rect 18061 13345 18095 13379
rect 46489 13345 46523 13379
rect 18153 13277 18187 13311
rect 19441 13277 19475 13311
rect 20085 13277 20119 13311
rect 46305 13277 46339 13311
rect 48145 13209 48179 13243
rect 18521 13141 18555 13175
rect 1593 12937 1627 12971
rect 17417 12937 17451 12971
rect 19625 12937 19659 12971
rect 18153 12869 18187 12903
rect 1409 12801 1443 12835
rect 17233 12801 17267 12835
rect 17417 12801 17451 12835
rect 17877 12801 17911 12835
rect 47777 12801 47811 12835
rect 46765 12189 46799 12223
rect 46857 12053 46891 12087
rect 18889 11781 18923 11815
rect 19625 11781 19659 11815
rect 17785 11713 17819 11747
rect 18797 11713 18831 11747
rect 19441 11645 19475 11679
rect 21281 11645 21315 11679
rect 17877 11509 17911 11543
rect 47777 11509 47811 11543
rect 16865 11169 16899 11203
rect 17049 11169 17083 11203
rect 17325 11169 17359 11203
rect 46305 11169 46339 11203
rect 46489 11169 46523 11203
rect 48145 11033 48179 11067
rect 46121 10693 46155 10727
rect 17877 10625 17911 10659
rect 18061 10557 18095 10591
rect 18337 10557 18371 10591
rect 46029 10557 46063 10591
rect 46305 10557 46339 10591
rect 47777 10421 47811 10455
rect 18153 10217 18187 10251
rect 46305 10081 46339 10115
rect 48145 10081 48179 10115
rect 18061 10013 18095 10047
rect 46489 9945 46523 9979
rect 46857 9673 46891 9707
rect 47685 9605 47719 9639
rect 47041 9537 47075 9571
rect 47593 9537 47627 9571
rect 47317 8925 47351 8959
rect 47593 8925 47627 8959
rect 47685 8449 47719 8483
rect 47869 8381 47903 8415
rect 46305 7905 46339 7939
rect 46489 7905 46523 7939
rect 47685 7905 47719 7939
rect 48145 7361 48179 7395
rect 47961 7157 47995 7191
rect 47041 6817 47075 6851
rect 48053 6817 48087 6851
rect 47133 6681 47167 6715
rect 46489 6273 46523 6307
rect 48145 6273 48179 6307
rect 46213 6205 46247 6239
rect 47961 6069 47995 6103
rect 47685 5729 47719 5763
rect 46305 5661 46339 5695
rect 46489 5593 46523 5627
rect 46029 5253 46063 5287
rect 46121 5253 46155 5287
rect 47593 5185 47627 5219
rect 46857 5117 46891 5151
rect 47685 4981 47719 5015
rect 46121 4641 46155 4675
rect 46581 4641 46615 4675
rect 7849 4573 7883 4607
rect 18521 4573 18555 4607
rect 19717 4573 19751 4607
rect 20361 4573 20395 4607
rect 21005 4573 21039 4607
rect 21649 4573 21683 4607
rect 21741 4573 21775 4607
rect 22293 4573 22327 4607
rect 22937 4573 22971 4607
rect 42901 4573 42935 4607
rect 45661 4573 45695 4607
rect 19809 4505 19843 4539
rect 46305 4505 46339 4539
rect 18613 4437 18647 4471
rect 20453 4437 20487 4471
rect 21097 4437 21131 4471
rect 22385 4437 22419 4471
rect 23029 4437 23063 4471
rect 20453 4233 20487 4267
rect 47777 4165 47811 4199
rect 2053 4097 2087 4131
rect 6653 4097 6687 4131
rect 7389 4097 7423 4131
rect 8217 4097 8251 4131
rect 18153 4097 18187 4131
rect 19073 4097 19107 4131
rect 19717 4097 19751 4131
rect 19809 4097 19843 4131
rect 20361 4097 20395 4131
rect 21005 4097 21039 4131
rect 22201 4097 22235 4131
rect 22845 4097 22879 4131
rect 23489 4097 23523 4131
rect 23581 4097 23615 4131
rect 24317 4097 24351 4131
rect 39957 4097 39991 4131
rect 42809 4097 42843 4131
rect 46489 4097 46523 4131
rect 21097 4029 21131 4063
rect 29469 4029 29503 4063
rect 29653 4029 29687 4063
rect 31309 4029 31343 4063
rect 43545 4029 43579 4063
rect 43729 4029 43763 4063
rect 44005 4029 44039 4063
rect 46213 4029 46247 4063
rect 22937 3961 22971 3995
rect 47961 3961 47995 3995
rect 2145 3893 2179 3927
rect 2881 3893 2915 3927
rect 6745 3893 6779 3927
rect 7481 3893 7515 3927
rect 8309 3893 8343 3927
rect 9413 3893 9447 3927
rect 11713 3893 11747 3927
rect 18245 3893 18279 3927
rect 19165 3893 19199 3927
rect 22293 3893 22327 3927
rect 24133 3893 24167 3927
rect 40049 3893 40083 3927
rect 42901 3893 42935 3927
rect 19533 3689 19567 3723
rect 20177 3689 20211 3723
rect 20821 3689 20855 3723
rect 22937 3689 22971 3723
rect 3985 3553 4019 3587
rect 6745 3553 6779 3587
rect 7113 3553 7147 3587
rect 9229 3553 9263 3587
rect 9689 3553 9723 3587
rect 29561 3553 29595 3587
rect 29745 3553 29779 3587
rect 37749 3553 37783 3587
rect 42625 3553 42659 3587
rect 42809 3553 42843 3587
rect 43177 3553 43211 3587
rect 45201 3553 45235 3587
rect 46305 3553 46339 3587
rect 46489 3553 46523 3587
rect 2697 3485 2731 3519
rect 6101 3485 6135 3519
rect 6561 3485 6595 3519
rect 12081 3485 12115 3519
rect 13553 3485 13587 3519
rect 14105 3485 14139 3519
rect 15301 3485 15335 3519
rect 17693 3485 17727 3519
rect 18337 3485 18371 3519
rect 19441 3485 19475 3519
rect 20085 3485 20119 3519
rect 20729 3485 20763 3519
rect 21373 3485 21407 3519
rect 22385 3485 22419 3519
rect 22845 3485 22879 3519
rect 23489 3485 23523 3519
rect 24685 3485 24719 3519
rect 25513 3485 25547 3519
rect 33057 3485 33091 3519
rect 33885 3485 33919 3519
rect 35909 3485 35943 3519
rect 39129 3485 39163 3519
rect 40049 3485 40083 3519
rect 40325 3485 40359 3519
rect 41337 3485 41371 3519
rect 41521 3485 41555 3519
rect 45661 3485 45695 3519
rect 1869 3417 1903 3451
rect 2237 3417 2271 3451
rect 9413 3417 9447 3451
rect 15485 3417 15519 3451
rect 17141 3417 17175 3451
rect 31401 3417 31435 3451
rect 36093 3417 36127 3451
rect 48145 3417 48179 3451
rect 2789 3349 2823 3383
rect 12173 3349 12207 3383
rect 14197 3349 14231 3383
rect 17785 3349 17819 3383
rect 18429 3349 18463 3383
rect 21465 3349 21499 3383
rect 23581 3349 23615 3383
rect 24777 3349 24811 3383
rect 33149 3349 33183 3383
rect 39221 3349 39255 3383
rect 41981 3349 42015 3383
rect 45753 3349 45787 3383
rect 17969 3145 18003 3179
rect 18613 3145 18647 3179
rect 19257 3145 19291 3179
rect 20085 3145 20119 3179
rect 20729 3145 20763 3179
rect 36185 3145 36219 3179
rect 1961 3077 1995 3111
rect 7849 3077 7883 3111
rect 10057 3077 10091 3111
rect 11713 3077 11747 3111
rect 14013 3077 14047 3111
rect 22293 3077 22327 3111
rect 24777 3077 24811 3111
rect 27629 3077 27663 3111
rect 33149 3077 33183 3111
rect 42625 3077 42659 3111
rect 44281 3077 44315 3111
rect 45385 3077 45419 3111
rect 1777 3009 1811 3043
rect 7665 3009 7699 3043
rect 9965 3009 9999 3043
rect 11529 3009 11563 3043
rect 13829 3009 13863 3043
rect 17049 3009 17083 3043
rect 17877 3009 17911 3043
rect 18521 3009 18555 3043
rect 19165 3009 19199 3043
rect 19993 3009 20027 3043
rect 20637 3009 20671 3043
rect 24593 3009 24627 3043
rect 27445 3009 27479 3043
rect 32965 3009 32999 3043
rect 36369 3009 36403 3043
rect 37933 3009 37967 3043
rect 38025 3009 38059 3043
rect 39681 3009 39715 3043
rect 42441 3009 42475 3043
rect 47777 3009 47811 3043
rect 2237 2941 2271 2975
rect 8125 2941 8159 2975
rect 11989 2941 12023 2975
rect 14289 2941 14323 2975
rect 16957 2941 16991 2975
rect 17417 2941 17451 2975
rect 22114 2941 22148 2975
rect 22937 2941 22971 2975
rect 25145 2941 25179 2975
rect 33517 2941 33551 2975
rect 38577 2941 38611 2975
rect 38761 2941 38795 2975
rect 39865 2941 39899 2975
rect 41521 2941 41555 2975
rect 45201 2941 45235 2975
rect 47041 2941 47075 2975
rect 39221 2873 39255 2907
rect 6837 2805 6871 2839
rect 47869 2805 47903 2839
rect 15577 2601 15611 2635
rect 17233 2601 17267 2635
rect 17877 2601 17911 2635
rect 23765 2601 23799 2635
rect 28641 2601 28675 2635
rect 38301 2601 38335 2635
rect 39221 2601 39255 2635
rect 40417 2601 40451 2635
rect 43545 2601 43579 2635
rect 44373 2601 44407 2635
rect 20545 2533 20579 2567
rect 22937 2533 22971 2567
rect 45569 2533 45603 2567
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2881 2465 2915 2499
rect 5273 2465 5307 2499
rect 6561 2465 6595 2499
rect 7021 2465 7055 2499
rect 18521 2465 18555 2499
rect 24685 2465 24719 2499
rect 25697 2465 25731 2499
rect 27261 2465 27295 2499
rect 30021 2465 30055 2499
rect 35817 2465 35851 2499
rect 41337 2465 41371 2499
rect 43085 2465 43119 2499
rect 46213 2465 46247 2499
rect 3801 2397 3835 2431
rect 4997 2397 5031 2431
rect 15761 2397 15795 2431
rect 17785 2397 17819 2431
rect 18429 2397 18463 2431
rect 19257 2397 19291 2431
rect 21281 2397 21315 2431
rect 21925 2397 21959 2431
rect 23029 2397 23063 2431
rect 23673 2397 23707 2431
rect 26985 2397 27019 2431
rect 29745 2397 29779 2431
rect 35541 2397 35575 2431
rect 38117 2397 38151 2431
rect 39129 2397 39163 2431
rect 41061 2397 41095 2431
rect 43729 2397 43763 2431
rect 44189 2397 44223 2431
rect 46489 2397 46523 2431
rect 6745 2329 6779 2363
rect 9413 2329 9447 2363
rect 17141 2329 17175 2363
rect 19349 2329 19383 2363
rect 20361 2329 20395 2363
rect 21097 2329 21131 2363
rect 24777 2329 24811 2363
rect 26249 2329 26283 2363
rect 28549 2329 28583 2363
rect 40325 2329 40359 2363
rect 42901 2329 42935 2363
rect 45385 2329 45419 2363
rect 47777 2329 47811 2363
rect 3985 2261 4019 2295
rect 9689 2261 9723 2295
rect 26341 2261 26375 2295
rect 47869 2261 47903 2295
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 29362 47200 29368 47252
rect 29420 47240 29426 47252
rect 29917 47243 29975 47249
rect 29917 47240 29929 47243
rect 29420 47212 29929 47240
rect 29420 47200 29426 47212
rect 29917 47209 29929 47212
rect 29963 47209 29975 47243
rect 29917 47203 29975 47209
rect 13357 47175 13415 47181
rect 13357 47141 13369 47175
rect 13403 47172 13415 47175
rect 17770 47172 17776 47184
rect 13403 47144 17776 47172
rect 13403 47141 13415 47144
rect 13357 47135 13415 47141
rect 17770 47132 17776 47144
rect 17828 47132 17834 47184
rect 19429 47175 19487 47181
rect 19429 47141 19441 47175
rect 19475 47172 19487 47175
rect 20254 47172 20260 47184
rect 19475 47144 20260 47172
rect 19475 47141 19487 47144
rect 19429 47135 19487 47141
rect 20254 47132 20260 47144
rect 20312 47132 20318 47184
rect 47949 47175 48007 47181
rect 47949 47172 47961 47175
rect 26206 47144 47961 47172
rect 11606 47064 11612 47116
rect 11664 47104 11670 47116
rect 11701 47107 11759 47113
rect 11701 47104 11713 47107
rect 11664 47076 11713 47104
rect 11664 47064 11670 47076
rect 11701 47073 11713 47076
rect 11747 47073 11759 47107
rect 20070 47104 20076 47116
rect 20031 47076 20076 47104
rect 11701 47067 11759 47073
rect 20070 47064 20076 47076
rect 20128 47064 20134 47116
rect 26206 47104 26234 47144
rect 47949 47141 47961 47144
rect 47995 47141 48007 47175
rect 47949 47135 48007 47141
rect 30742 47104 30748 47116
rect 20180 47076 26234 47104
rect 30703 47076 30748 47104
rect 1946 47036 1952 47048
rect 1907 47008 1952 47036
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 2590 46996 2596 47048
rect 2648 47036 2654 47048
rect 2685 47039 2743 47045
rect 2685 47036 2697 47039
rect 2648 47008 2697 47036
rect 2648 46996 2654 47008
rect 2685 47005 2697 47008
rect 2731 47005 2743 47039
rect 2685 46999 2743 47005
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4798 47036 4804 47048
rect 4759 47008 4804 47036
rect 3789 46999 3847 47005
rect 4798 46996 4804 47008
rect 4856 46996 4862 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6825 47039 6883 47045
rect 6825 47036 6837 47039
rect 5868 47008 6837 47036
rect 5868 46996 5874 47008
rect 6825 47005 6837 47008
rect 6871 47005 6883 47039
rect 6825 46999 6883 47005
rect 7098 46996 7104 47048
rect 7156 47036 7162 47048
rect 7745 47039 7803 47045
rect 7745 47036 7757 47039
rect 7156 47008 7757 47036
rect 7156 46996 7162 47008
rect 7745 47005 7757 47008
rect 7791 47005 7803 47039
rect 7745 46999 7803 47005
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 9088 47008 9413 47036
rect 9088 46996 9094 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 11974 47036 11980 47048
rect 11935 47008 11980 47036
rect 9401 46999 9459 47005
rect 11974 46996 11980 47008
rect 12032 46996 12038 47048
rect 12894 46996 12900 47048
rect 12952 47036 12958 47048
rect 13081 47039 13139 47045
rect 13081 47036 13093 47039
rect 12952 47008 13093 47036
rect 12952 46996 12958 47008
rect 13081 47005 13093 47008
rect 13127 47005 13139 47039
rect 13081 46999 13139 47005
rect 13814 46996 13820 47048
rect 13872 47036 13878 47048
rect 14553 47039 14611 47045
rect 14553 47036 14565 47039
rect 13872 47008 14565 47036
rect 13872 46996 13878 47008
rect 14553 47005 14565 47008
rect 14599 47005 14611 47039
rect 14553 46999 14611 47005
rect 16482 46996 16488 47048
rect 16540 47036 16546 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16540 47008 16681 47036
rect 16540 46996 16546 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16669 46999 16727 47005
rect 16945 47039 17003 47045
rect 16945 47005 16957 47039
rect 16991 47005 17003 47039
rect 16945 46999 17003 47005
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 7834 46928 7840 46980
rect 7892 46968 7898 46980
rect 7929 46971 7987 46977
rect 7929 46968 7941 46971
rect 7892 46940 7941 46968
rect 7892 46928 7898 46940
rect 7929 46937 7941 46940
rect 7975 46937 7987 46971
rect 7929 46931 7987 46937
rect 9490 46928 9496 46980
rect 9548 46968 9554 46980
rect 9585 46971 9643 46977
rect 9585 46968 9597 46971
rect 9548 46940 9597 46968
rect 9548 46928 9554 46940
rect 9585 46937 9597 46940
rect 9631 46937 9643 46971
rect 9585 46931 9643 46937
rect 14642 46928 14648 46980
rect 14700 46968 14706 46980
rect 14737 46971 14795 46977
rect 14737 46968 14749 46971
rect 14700 46940 14749 46968
rect 14700 46928 14706 46940
rect 14737 46937 14749 46940
rect 14783 46937 14795 46971
rect 16960 46968 16988 46999
rect 18690 46996 18696 47048
rect 18748 47036 18754 47048
rect 19245 47039 19303 47045
rect 19245 47036 19257 47039
rect 18748 47008 19257 47036
rect 18748 46996 18754 47008
rect 19245 47005 19257 47008
rect 19291 47005 19303 47039
rect 19245 46999 19303 47005
rect 19978 46996 19984 47048
rect 20036 47036 20042 47048
rect 20180 47036 20208 47076
rect 30742 47064 30748 47076
rect 30800 47064 30806 47116
rect 44453 47107 44511 47113
rect 44453 47073 44465 47107
rect 44499 47104 44511 47107
rect 45094 47104 45100 47116
rect 44499 47076 45100 47104
rect 44499 47073 44511 47076
rect 44453 47067 44511 47073
rect 45094 47064 45100 47076
rect 45152 47064 45158 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 20036 47008 20208 47036
rect 20349 47039 20407 47045
rect 20036 46996 20042 47008
rect 20349 47005 20361 47039
rect 20395 47036 20407 47039
rect 20438 47036 20444 47048
rect 20395 47008 20444 47036
rect 20395 47005 20407 47008
rect 20349 46999 20407 47005
rect 20438 46996 20444 47008
rect 20496 46996 20502 47048
rect 25682 47036 25688 47048
rect 25643 47008 25688 47036
rect 25682 46996 25688 47008
rect 25740 46996 25746 47048
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28629 47039 28687 47045
rect 28629 47036 28641 47039
rect 28408 47008 28641 47036
rect 28408 46996 28414 47008
rect 28629 47005 28641 47008
rect 28675 47005 28687 47039
rect 28629 46999 28687 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 31021 47039 31079 47045
rect 31021 47005 31033 47039
rect 31067 47036 31079 47039
rect 31110 47036 31116 47048
rect 31067 47008 31116 47036
rect 31067 47005 31079 47008
rect 31021 46999 31079 47005
rect 31110 46996 31116 47008
rect 31168 46996 31174 47048
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38381 47039 38439 47045
rect 38381 47036 38393 47039
rect 38160 47008 38393 47036
rect 38160 46996 38166 47008
rect 38381 47005 38393 47008
rect 38427 47005 38439 47039
rect 38381 46999 38439 47005
rect 42518 46996 42524 47048
rect 42576 47036 42582 47048
rect 42613 47039 42671 47045
rect 42613 47036 42625 47039
rect 42576 47008 42625 47036
rect 42576 46996 42582 47008
rect 42613 47005 42625 47008
rect 42659 47005 42671 47039
rect 45186 47036 45192 47048
rect 45147 47008 45192 47036
rect 42613 46999 42671 47005
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47765 47039 47823 47045
rect 47765 47036 47777 47039
rect 47728 47008 47777 47036
rect 47728 46996 47734 47008
rect 47765 47005 47777 47008
rect 47811 47005 47823 47039
rect 47765 46999 47823 47005
rect 22922 46968 22928 46980
rect 16960 46940 22928 46968
rect 14737 46931 14795 46937
rect 22922 46928 22928 46940
rect 22980 46928 22986 46980
rect 40313 46971 40371 46977
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 40313 46931 40371 46937
rect 2130 46900 2136 46912
rect 2091 46872 2136 46900
rect 2130 46860 2136 46872
rect 2188 46860 2194 46912
rect 2866 46900 2872 46912
rect 2827 46872 2872 46900
rect 2866 46860 2872 46872
rect 2924 46860 2930 46912
rect 4890 46900 4896 46912
rect 4851 46872 4896 46900
rect 4890 46860 4896 46872
rect 4948 46860 4954 46912
rect 6914 46860 6920 46912
rect 6972 46900 6978 46912
rect 6972 46872 7017 46900
rect 6972 46860 6978 46872
rect 27062 46860 27068 46912
rect 27120 46900 27126 46912
rect 27614 46900 27620 46912
rect 27120 46872 27620 46900
rect 27120 46860 27126 46872
rect 27614 46860 27620 46872
rect 27672 46860 27678 46912
rect 28258 46860 28264 46912
rect 28316 46900 28322 46912
rect 28445 46903 28503 46909
rect 28445 46900 28457 46903
rect 28316 46872 28457 46900
rect 28316 46860 28322 46872
rect 28445 46869 28457 46872
rect 28491 46869 28503 46903
rect 28445 46863 28503 46869
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 40402 46928 40408 46980
rect 40460 46968 40466 46980
rect 40497 46971 40555 46977
rect 40497 46968 40509 46971
rect 40460 46940 40509 46968
rect 40460 46928 40466 46940
rect 40497 46937 40509 46940
rect 40543 46937 40555 46971
rect 42794 46968 42800 46980
rect 42755 46940 42800 46968
rect 40497 46931 40555 46937
rect 42794 46928 42800 46940
rect 42852 46928 42858 46980
rect 45370 46968 45376 46980
rect 45331 46940 45376 46968
rect 45370 46928 45376 46940
rect 45428 46928 45434 46980
rect 39356 46872 40356 46900
rect 39356 46860 39362 46872
rect 41230 46860 41236 46912
rect 41288 46900 41294 46912
rect 41782 46900 41788 46912
rect 41288 46872 41788 46900
rect 41288 46860 41294 46872
rect 41782 46860 41788 46872
rect 41840 46860 41846 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 2866 46588 2872 46640
rect 2924 46628 2930 46640
rect 28445 46631 28503 46637
rect 28445 46628 28457 46631
rect 2924 46600 28457 46628
rect 2924 46588 2930 46600
rect 28445 46597 28457 46600
rect 28491 46597 28503 46631
rect 28445 46591 28503 46597
rect 1394 46560 1400 46572
rect 1355 46532 1400 46560
rect 1394 46520 1400 46532
rect 1452 46520 1458 46572
rect 12250 46520 12256 46572
rect 12308 46560 12314 46572
rect 12437 46563 12495 46569
rect 12437 46560 12449 46563
rect 12308 46532 12449 46560
rect 12308 46520 12314 46532
rect 12437 46529 12449 46532
rect 12483 46529 12495 46563
rect 28258 46560 28264 46572
rect 28219 46532 28264 46560
rect 12437 46523 12495 46529
rect 28258 46520 28264 46532
rect 28316 46520 28322 46572
rect 38102 46560 38108 46572
rect 38063 46532 38108 46560
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 47854 46560 47860 46572
rect 47815 46532 47860 46560
rect 47854 46520 47860 46532
rect 47912 46520 47918 46572
rect 13538 46452 13544 46504
rect 13596 46492 13602 46504
rect 13633 46495 13691 46501
rect 13633 46492 13645 46495
rect 13596 46464 13645 46492
rect 13596 46452 13602 46464
rect 13633 46461 13645 46464
rect 13679 46461 13691 46495
rect 13633 46455 13691 46461
rect 13817 46495 13875 46501
rect 13817 46461 13829 46495
rect 13863 46492 13875 46495
rect 14182 46492 14188 46504
rect 13863 46464 14188 46492
rect 13863 46461 13875 46464
rect 13817 46455 13875 46461
rect 14182 46452 14188 46464
rect 14240 46452 14246 46504
rect 14274 46452 14280 46504
rect 14332 46492 14338 46504
rect 18969 46495 19027 46501
rect 14332 46464 14377 46492
rect 14332 46452 14338 46464
rect 18969 46461 18981 46495
rect 19015 46492 19027 46495
rect 19429 46495 19487 46501
rect 19429 46492 19441 46495
rect 19015 46464 19441 46492
rect 19015 46461 19027 46464
rect 18969 46455 19027 46461
rect 19429 46461 19441 46464
rect 19475 46461 19487 46495
rect 19610 46492 19616 46504
rect 19571 46464 19616 46492
rect 19429 46455 19487 46461
rect 19610 46452 19616 46464
rect 19668 46452 19674 46504
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 24581 46495 24639 46501
rect 24581 46461 24593 46495
rect 24627 46461 24639 46495
rect 24581 46455 24639 46461
rect 24765 46495 24823 46501
rect 24765 46461 24777 46495
rect 24811 46492 24823 46495
rect 24946 46492 24952 46504
rect 24811 46464 24952 46492
rect 24811 46461 24823 46464
rect 24765 46455 24823 46461
rect 24596 46424 24624 46455
rect 24946 46452 24952 46464
rect 25004 46452 25010 46504
rect 25774 46492 25780 46504
rect 25735 46464 25780 46492
rect 25774 46452 25780 46464
rect 25832 46452 25838 46504
rect 30101 46495 30159 46501
rect 30101 46461 30113 46495
rect 30147 46492 30159 46495
rect 38286 46492 38292 46504
rect 30147 46464 35894 46492
rect 38247 46464 38292 46492
rect 30147 46461 30159 46464
rect 30101 46455 30159 46461
rect 27157 46427 27215 46433
rect 27157 46424 27169 46427
rect 24596 46396 27169 46424
rect 27157 46393 27169 46396
rect 27203 46393 27215 46427
rect 35866 46424 35894 46464
rect 38286 46452 38292 46464
rect 38344 46452 38350 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 41877 46495 41935 46501
rect 41877 46461 41889 46495
rect 41923 46492 41935 46495
rect 42429 46495 42487 46501
rect 42429 46492 42441 46495
rect 41923 46464 42441 46492
rect 41923 46461 41935 46464
rect 41877 46455 41935 46461
rect 42429 46461 42441 46464
rect 42475 46461 42487 46495
rect 42610 46492 42616 46504
rect 42571 46464 42616 46492
rect 42429 46455 42487 46461
rect 42610 46452 42616 46464
rect 42668 46452 42674 46504
rect 42702 46452 42708 46504
rect 42760 46492 42766 46504
rect 42889 46495 42947 46501
rect 42889 46492 42901 46495
rect 42760 46464 42901 46492
rect 42760 46452 42766 46464
rect 42889 46461 42901 46464
rect 42935 46461 42947 46495
rect 42889 46455 42947 46461
rect 45189 46495 45247 46501
rect 45189 46461 45201 46495
rect 45235 46461 45247 46495
rect 45189 46455 45247 46461
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 46014 46492 46020 46504
rect 45419 46464 46020 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 44266 46424 44272 46436
rect 35866 46396 44272 46424
rect 27157 46387 27215 46393
rect 44266 46384 44272 46396
rect 44324 46384 44330 46436
rect 45204 46424 45232 46455
rect 46014 46452 46020 46464
rect 46072 46452 46078 46504
rect 46842 46492 46848 46504
rect 46803 46464 46848 46492
rect 46842 46452 46848 46464
rect 46900 46452 46906 46504
rect 46934 46424 46940 46436
rect 45204 46396 46940 46424
rect 46934 46384 46940 46396
rect 46992 46384 46998 46436
rect 1581 46359 1639 46365
rect 1581 46325 1593 46359
rect 1627 46356 1639 46359
rect 1670 46356 1676 46368
rect 1627 46328 1676 46356
rect 1627 46325 1639 46328
rect 1581 46319 1639 46325
rect 1670 46316 1676 46328
rect 1728 46316 1734 46368
rect 2314 46356 2320 46368
rect 2275 46328 2320 46356
rect 2314 46316 2320 46328
rect 2372 46316 2378 46368
rect 4433 46359 4491 46365
rect 4433 46325 4445 46359
rect 4479 46356 4491 46359
rect 4614 46356 4620 46368
rect 4479 46328 4620 46356
rect 4479 46325 4491 46328
rect 4433 46319 4491 46325
rect 4614 46316 4620 46328
rect 4672 46316 4678 46368
rect 10410 46316 10416 46368
rect 10468 46356 10474 46368
rect 10689 46359 10747 46365
rect 10689 46356 10701 46359
rect 10468 46328 10701 46356
rect 10468 46316 10474 46328
rect 10689 46325 10701 46328
rect 10735 46325 10747 46359
rect 12526 46356 12532 46368
rect 12487 46328 12532 46356
rect 10689 46319 10747 46325
rect 12526 46316 12532 46328
rect 12584 46316 12590 46368
rect 20070 46316 20076 46368
rect 20128 46356 20134 46368
rect 22005 46359 22063 46365
rect 22005 46356 22017 46359
rect 20128 46328 22017 46356
rect 20128 46316 20134 46328
rect 22005 46325 22017 46328
rect 22051 46325 22063 46359
rect 22005 46319 22063 46325
rect 31662 46316 31668 46368
rect 31720 46356 31726 46368
rect 32309 46359 32367 46365
rect 32309 46356 32321 46359
rect 31720 46328 32321 46356
rect 31720 46316 31726 46328
rect 32309 46325 32321 46328
rect 32355 46325 32367 46359
rect 41230 46356 41236 46368
rect 41191 46328 41236 46356
rect 32309 46319 32367 46325
rect 41230 46316 41236 46328
rect 41288 46316 41294 46368
rect 48038 46356 48044 46368
rect 47999 46328 48044 46356
rect 48038 46316 48044 46328
rect 48096 46316 48102 46368
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 13538 46152 13544 46164
rect 13499 46124 13544 46152
rect 13538 46112 13544 46124
rect 13596 46112 13602 46164
rect 14182 46152 14188 46164
rect 14143 46124 14188 46152
rect 14182 46112 14188 46124
rect 14240 46112 14246 46164
rect 18601 46155 18659 46161
rect 18601 46121 18613 46155
rect 18647 46152 18659 46155
rect 19610 46152 19616 46164
rect 18647 46124 19616 46152
rect 18647 46121 18659 46124
rect 18601 46115 18659 46121
rect 19610 46112 19616 46124
rect 19668 46112 19674 46164
rect 24946 46112 24952 46164
rect 25004 46152 25010 46164
rect 25406 46152 25412 46164
rect 25004 46124 25412 46152
rect 25004 46112 25010 46124
rect 25406 46112 25412 46124
rect 25464 46112 25470 46164
rect 38286 46152 38292 46164
rect 38247 46124 38292 46152
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 3878 46044 3884 46096
rect 3936 46084 3942 46096
rect 3936 46056 4752 46084
rect 3936 46044 3942 46056
rect 1397 46019 1455 46025
rect 1397 45985 1409 46019
rect 1443 46016 1455 46019
rect 2314 46016 2320 46028
rect 1443 45988 2320 46016
rect 1443 45985 1455 45988
rect 1397 45979 1455 45985
rect 2314 45976 2320 45988
rect 2372 45976 2378 46028
rect 2774 46016 2780 46028
rect 2735 45988 2780 46016
rect 2774 45976 2780 45988
rect 2832 45976 2838 46028
rect 4157 46019 4215 46025
rect 4157 45985 4169 46019
rect 4203 46016 4215 46019
rect 4614 46016 4620 46028
rect 4203 45988 4620 46016
rect 4203 45985 4215 45988
rect 4157 45979 4215 45985
rect 4614 45976 4620 45988
rect 4672 45976 4678 46028
rect 4724 46025 4752 46056
rect 25130 46044 25136 46096
rect 25188 46084 25194 46096
rect 45922 46084 45928 46096
rect 25188 46056 25912 46084
rect 25188 46044 25194 46056
rect 4709 46019 4767 46025
rect 4709 45985 4721 46019
rect 4755 45985 4767 46019
rect 10410 46016 10416 46028
rect 10371 45988 10416 46016
rect 4709 45979 4767 45985
rect 10410 45976 10416 45988
rect 10468 45976 10474 46028
rect 10962 45976 10968 46028
rect 11020 46016 11026 46028
rect 11057 46019 11115 46025
rect 11057 46016 11069 46019
rect 11020 45988 11069 46016
rect 11020 45976 11026 45988
rect 11057 45985 11069 45988
rect 11103 45985 11115 46019
rect 20070 46016 20076 46028
rect 20031 45988 20076 46016
rect 11057 45979 11115 45985
rect 20070 45976 20076 45988
rect 20128 45976 20134 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 25409 46019 25467 46025
rect 25409 45985 25421 46019
rect 25455 46016 25467 46019
rect 25682 46016 25688 46028
rect 25455 45988 25688 46016
rect 25455 45985 25467 45988
rect 25409 45979 25467 45985
rect 25682 45976 25688 45988
rect 25740 45976 25746 46028
rect 25884 46025 25912 46056
rect 38212 46056 45928 46084
rect 25869 46019 25927 46025
rect 25869 45985 25881 46019
rect 25915 45985 25927 46019
rect 31662 46016 31668 46028
rect 31623 45988 31668 46016
rect 25869 45979 25927 45985
rect 31662 45976 31668 45988
rect 31720 45976 31726 46028
rect 32214 46016 32220 46028
rect 32175 45988 32220 46016
rect 32214 45976 32220 45988
rect 32272 45976 32278 46028
rect 38212 45960 38240 46056
rect 45922 46044 45928 46056
rect 45980 46044 45986 46096
rect 41230 46016 41236 46028
rect 41191 45988 41236 46016
rect 41230 45976 41236 45988
rect 41288 45976 41294 46028
rect 41874 46016 41880 46028
rect 41835 45988 41880 46016
rect 41874 45976 41880 45988
rect 41932 45976 41938 46028
rect 47026 46016 47032 46028
rect 46987 45988 47032 46016
rect 47026 45976 47032 45988
rect 47084 45976 47090 46028
rect 14090 45948 14096 45960
rect 14003 45920 14096 45948
rect 14090 45908 14096 45920
rect 14148 45948 14154 45960
rect 18509 45951 18567 45957
rect 18509 45948 18521 45951
rect 14148 45920 18521 45948
rect 14148 45908 14154 45920
rect 18509 45917 18521 45920
rect 18555 45948 18567 45951
rect 18782 45948 18788 45960
rect 18555 45920 18788 45948
rect 18555 45917 18567 45920
rect 18509 45911 18567 45917
rect 18782 45908 18788 45920
rect 18840 45908 18846 45960
rect 19429 45951 19487 45957
rect 19429 45917 19441 45951
rect 19475 45917 19487 45951
rect 38194 45948 38200 45960
rect 38107 45920 38200 45948
rect 19429 45911 19487 45917
rect 1581 45883 1639 45889
rect 1581 45849 1593 45883
rect 1627 45880 1639 45883
rect 2314 45880 2320 45892
rect 1627 45852 2320 45880
rect 1627 45849 1639 45852
rect 1581 45843 1639 45849
rect 2314 45840 2320 45852
rect 2372 45840 2378 45892
rect 4341 45883 4399 45889
rect 4341 45849 4353 45883
rect 4387 45880 4399 45883
rect 5074 45880 5080 45892
rect 4387 45852 5080 45880
rect 4387 45849 4399 45852
rect 4341 45843 4399 45849
rect 5074 45840 5080 45852
rect 5132 45840 5138 45892
rect 10594 45880 10600 45892
rect 10555 45852 10600 45880
rect 10594 45840 10600 45852
rect 10652 45840 10658 45892
rect 16666 45840 16672 45892
rect 16724 45880 16730 45892
rect 19444 45880 19472 45911
rect 38194 45908 38200 45920
rect 38252 45908 38258 45960
rect 43806 45908 43812 45960
rect 43864 45948 43870 45960
rect 43901 45951 43959 45957
rect 43901 45948 43913 45951
rect 43864 45920 43913 45948
rect 43864 45908 43870 45920
rect 43901 45917 43913 45920
rect 43947 45917 43959 45951
rect 43901 45911 43959 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45948 45707 45951
rect 45738 45948 45744 45960
rect 45695 45920 45744 45948
rect 45695 45917 45707 45920
rect 45649 45911 45707 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 46290 45948 46296 45960
rect 46251 45920 46296 45948
rect 46290 45908 46296 45920
rect 46348 45908 46354 45960
rect 16724 45852 19472 45880
rect 19521 45883 19579 45889
rect 16724 45840 16730 45852
rect 19521 45849 19533 45883
rect 19567 45880 19579 45883
rect 20257 45883 20315 45889
rect 20257 45880 20269 45883
rect 19567 45852 20269 45880
rect 19567 45849 19579 45852
rect 19521 45843 19579 45849
rect 20257 45849 20269 45852
rect 20303 45849 20315 45883
rect 20257 45843 20315 45849
rect 25593 45883 25651 45889
rect 25593 45849 25605 45883
rect 25639 45880 25651 45883
rect 27062 45880 27068 45892
rect 25639 45852 27068 45880
rect 25639 45849 25651 45852
rect 25593 45843 25651 45849
rect 27062 45840 27068 45852
rect 27120 45840 27126 45892
rect 31849 45883 31907 45889
rect 31849 45849 31861 45883
rect 31895 45880 31907 45883
rect 32214 45880 32220 45892
rect 31895 45852 32220 45880
rect 31895 45849 31907 45852
rect 31849 45843 31907 45849
rect 32214 45840 32220 45852
rect 32272 45840 32278 45892
rect 41414 45880 41420 45892
rect 41375 45852 41420 45880
rect 41414 45840 41420 45852
rect 41472 45840 41478 45892
rect 46474 45880 46480 45892
rect 46435 45852 46480 45880
rect 46474 45840 46480 45852
rect 46532 45840 46538 45892
rect 43990 45772 43996 45824
rect 44048 45812 44054 45824
rect 44085 45815 44143 45821
rect 44085 45812 44097 45815
rect 44048 45784 44097 45812
rect 44048 45772 44054 45784
rect 44085 45781 44097 45784
rect 44131 45781 44143 45815
rect 44085 45775 44143 45781
rect 45741 45815 45799 45821
rect 45741 45781 45753 45815
rect 45787 45812 45799 45815
rect 46566 45812 46572 45824
rect 45787 45784 46572 45812
rect 45787 45781 45799 45784
rect 45741 45775 45799 45781
rect 46566 45772 46572 45784
rect 46624 45772 46630 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 2314 45608 2320 45620
rect 2275 45580 2320 45608
rect 2314 45568 2320 45580
rect 2372 45568 2378 45620
rect 5074 45608 5080 45620
rect 5035 45580 5080 45608
rect 5074 45568 5080 45580
rect 5132 45568 5138 45620
rect 10594 45608 10600 45620
rect 10555 45580 10600 45608
rect 10594 45568 10600 45580
rect 10652 45568 10658 45620
rect 32214 45608 32220 45620
rect 32175 45580 32220 45608
rect 32214 45568 32220 45580
rect 32272 45568 32278 45620
rect 41414 45608 41420 45620
rect 41375 45580 41420 45608
rect 41414 45568 41420 45580
rect 41472 45568 41478 45620
rect 18322 45540 18328 45552
rect 6886 45512 18328 45540
rect 2225 45475 2283 45481
rect 2225 45441 2237 45475
rect 2271 45472 2283 45475
rect 2314 45472 2320 45484
rect 2271 45444 2320 45472
rect 2271 45441 2283 45444
rect 2225 45435 2283 45441
rect 2314 45432 2320 45444
rect 2372 45432 2378 45484
rect 4985 45475 5043 45481
rect 4985 45441 4997 45475
rect 5031 45472 5043 45475
rect 6886 45472 6914 45512
rect 18322 45500 18328 45512
rect 18380 45500 18386 45552
rect 25406 45540 25412 45552
rect 25367 45512 25412 45540
rect 25406 45500 25412 45512
rect 25464 45500 25470 45552
rect 27062 45540 27068 45552
rect 27023 45512 27068 45540
rect 27062 45500 27068 45512
rect 27120 45500 27126 45552
rect 45094 45540 45100 45552
rect 45055 45512 45100 45540
rect 45094 45500 45100 45512
rect 45152 45500 45158 45552
rect 45370 45500 45376 45552
rect 45428 45540 45434 45552
rect 47673 45543 47731 45549
rect 47673 45540 47685 45543
rect 45428 45512 47685 45540
rect 45428 45500 45434 45512
rect 47673 45509 47685 45512
rect 47719 45509 47731 45543
rect 47673 45503 47731 45509
rect 5031 45444 6914 45472
rect 10505 45475 10563 45481
rect 5031 45441 5043 45444
rect 4985 45435 5043 45441
rect 10505 45441 10517 45475
rect 10551 45472 10563 45475
rect 16666 45472 16672 45484
rect 10551 45444 16672 45472
rect 10551 45441 10563 45444
rect 10505 45435 10563 45441
rect 2332 45404 2360 45432
rect 10520 45404 10548 45435
rect 16666 45432 16672 45444
rect 16724 45432 16730 45484
rect 25314 45472 25320 45484
rect 25275 45444 25320 45472
rect 25314 45432 25320 45444
rect 25372 45432 25378 45484
rect 26510 45432 26516 45484
rect 26568 45472 26574 45484
rect 26973 45475 27031 45481
rect 26973 45472 26985 45475
rect 26568 45444 26985 45472
rect 26568 45432 26574 45444
rect 26973 45441 26985 45444
rect 27019 45441 27031 45475
rect 26973 45435 27031 45441
rect 31938 45432 31944 45484
rect 31996 45472 32002 45484
rect 32125 45475 32183 45481
rect 32125 45472 32137 45475
rect 31996 45444 32137 45472
rect 31996 45432 32002 45444
rect 32125 45441 32137 45444
rect 32171 45441 32183 45475
rect 41322 45472 41328 45484
rect 41283 45444 41328 45472
rect 32125 45435 32183 45441
rect 41322 45432 41328 45444
rect 41380 45432 41386 45484
rect 46198 45472 46204 45484
rect 46159 45444 46204 45472
rect 46198 45432 46204 45444
rect 46256 45432 46262 45484
rect 47486 45432 47492 45484
rect 47544 45472 47550 45484
rect 47581 45475 47639 45481
rect 47581 45472 47593 45475
rect 47544 45444 47593 45472
rect 47544 45432 47550 45444
rect 47581 45441 47593 45444
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 42702 45404 42708 45416
rect 2332 45376 10548 45404
rect 42663 45376 42708 45404
rect 42702 45364 42708 45376
rect 42760 45364 42766 45416
rect 42889 45407 42947 45413
rect 42889 45373 42901 45407
rect 42935 45404 42947 45407
rect 43806 45404 43812 45416
rect 42935 45376 43812 45404
rect 42935 45373 42947 45376
rect 42889 45367 42947 45373
rect 43806 45364 43812 45376
rect 43864 45364 43870 45416
rect 44082 45404 44088 45416
rect 44043 45376 44088 45404
rect 44082 45364 44088 45376
rect 44140 45364 44146 45416
rect 45830 45364 45836 45416
rect 45888 45404 45894 45416
rect 46477 45407 46535 45413
rect 46477 45404 46489 45407
rect 45888 45376 46489 45404
rect 45888 45364 45894 45376
rect 46477 45373 46489 45376
rect 46523 45373 46535 45407
rect 46477 45367 46535 45373
rect 25314 45296 25320 45348
rect 25372 45336 25378 45348
rect 45646 45336 45652 45348
rect 25372 45308 45652 45336
rect 25372 45296 25378 45308
rect 45646 45296 45652 45308
rect 45704 45296 45710 45348
rect 45094 45228 45100 45280
rect 45152 45268 45158 45280
rect 45189 45271 45247 45277
rect 45189 45268 45201 45271
rect 45152 45240 45201 45268
rect 45152 45228 45158 45240
rect 45189 45237 45201 45240
rect 45235 45237 45247 45271
rect 45189 45231 45247 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 42061 45067 42119 45073
rect 42061 45033 42073 45067
rect 42107 45064 42119 45067
rect 42610 45064 42616 45076
rect 42107 45036 42616 45064
rect 42107 45033 42119 45036
rect 42061 45027 42119 45033
rect 42610 45024 42616 45036
rect 42668 45024 42674 45076
rect 42794 45024 42800 45076
rect 42852 45064 42858 45076
rect 43165 45067 43223 45073
rect 43165 45064 43177 45067
rect 42852 45036 43177 45064
rect 42852 45024 42858 45036
rect 43165 45033 43177 45036
rect 43211 45033 43223 45067
rect 43806 45064 43812 45076
rect 43767 45036 43812 45064
rect 43165 45027 43223 45033
rect 43806 45024 43812 45036
rect 43864 45024 43870 45076
rect 45741 45067 45799 45073
rect 45741 45033 45753 45067
rect 45787 45064 45799 45067
rect 46474 45064 46480 45076
rect 45787 45036 46480 45064
rect 45787 45033 45799 45036
rect 45741 45027 45799 45033
rect 46474 45024 46480 45036
rect 46532 45024 46538 45076
rect 45189 44999 45247 45005
rect 45189 44965 45201 44999
rect 45235 44996 45247 44999
rect 46290 44996 46296 45008
rect 45235 44968 46296 44996
rect 45235 44965 45247 44968
rect 45189 44959 45247 44965
rect 46290 44956 46296 44968
rect 46348 44956 46354 45008
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 28169 44863 28227 44869
rect 28169 44829 28181 44863
rect 28215 44860 28227 44863
rect 29546 44860 29552 44872
rect 28215 44832 29552 44860
rect 28215 44829 28227 44832
rect 28169 44823 28227 44829
rect 29546 44820 29552 44832
rect 29604 44820 29610 44872
rect 41969 44863 42027 44869
rect 41969 44829 41981 44863
rect 42015 44860 42027 44863
rect 42058 44860 42064 44872
rect 42015 44832 42064 44860
rect 42015 44829 42027 44832
rect 41969 44823 42027 44829
rect 42058 44820 42064 44832
rect 42116 44820 42122 44872
rect 43070 44860 43076 44872
rect 43031 44832 43076 44860
rect 43070 44820 43076 44832
rect 43128 44820 43134 44872
rect 43717 44863 43775 44869
rect 43717 44829 43729 44863
rect 43763 44860 43775 44863
rect 45646 44860 45652 44872
rect 43763 44832 45554 44860
rect 45607 44832 45652 44860
rect 43763 44829 43775 44832
rect 43717 44823 43775 44829
rect 28074 44684 28080 44736
rect 28132 44724 28138 44736
rect 28261 44727 28319 44733
rect 28261 44724 28273 44727
rect 28132 44696 28273 44724
rect 28132 44684 28138 44696
rect 28261 44693 28273 44696
rect 28307 44693 28319 44727
rect 45526 44724 45554 44832
rect 45646 44820 45652 44832
rect 45704 44820 45710 44872
rect 45738 44820 45744 44872
rect 45796 44860 45802 44872
rect 46293 44863 46351 44869
rect 46293 44860 46305 44863
rect 45796 44832 46305 44860
rect 45796 44820 45802 44832
rect 46293 44829 46305 44832
rect 46339 44829 46351 44863
rect 46293 44823 46351 44829
rect 46477 44795 46535 44801
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 46658 44792 46664 44804
rect 46523 44764 46664 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 46658 44752 46664 44764
rect 46716 44752 46722 44804
rect 47578 44724 47584 44736
rect 45526 44696 47584 44724
rect 28261 44687 28319 44693
rect 47578 44684 47584 44696
rect 47636 44684 47642 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 46014 44520 46020 44532
rect 45975 44492 46020 44520
rect 46014 44480 46020 44492
rect 46072 44480 46078 44532
rect 46658 44520 46664 44532
rect 46619 44492 46664 44520
rect 46658 44480 46664 44492
rect 46716 44480 46722 44532
rect 28074 44452 28080 44464
rect 28035 44424 28080 44452
rect 28074 44412 28080 44424
rect 28132 44412 28138 44464
rect 41322 44412 41328 44464
rect 41380 44452 41386 44464
rect 41380 44424 46612 44452
rect 41380 44412 41386 44424
rect 42702 44344 42708 44396
rect 42760 44384 42766 44396
rect 42889 44387 42947 44393
rect 42889 44384 42901 44387
rect 42760 44356 42901 44384
rect 42760 44344 42766 44356
rect 42889 44353 42901 44356
rect 42935 44353 42947 44387
rect 42889 44347 42947 44353
rect 45465 44387 45523 44393
rect 45465 44353 45477 44387
rect 45511 44384 45523 44387
rect 45738 44384 45744 44396
rect 45511 44356 45744 44384
rect 45511 44353 45523 44356
rect 45465 44347 45523 44353
rect 45738 44344 45744 44356
rect 45796 44344 45802 44396
rect 45922 44384 45928 44396
rect 45883 44356 45928 44384
rect 45922 44344 45928 44356
rect 45980 44344 45986 44396
rect 46584 44393 46612 44424
rect 46569 44387 46627 44393
rect 46569 44353 46581 44387
rect 46615 44353 46627 44387
rect 46569 44347 46627 44353
rect 47486 44344 47492 44396
rect 47544 44384 47550 44396
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 47544 44356 47593 44384
rect 47544 44344 47550 44356
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 3510 44276 3516 44328
rect 3568 44316 3574 44328
rect 3568 44288 6914 44316
rect 3568 44276 3574 44288
rect 6886 44248 6914 44288
rect 27706 44276 27712 44328
rect 27764 44316 27770 44328
rect 27893 44319 27951 44325
rect 27893 44316 27905 44319
rect 27764 44288 27905 44316
rect 27764 44276 27770 44288
rect 27893 44285 27905 44288
rect 27939 44285 27951 44319
rect 27893 44279 27951 44285
rect 28353 44319 28411 44325
rect 28353 44285 28365 44319
rect 28399 44285 28411 44319
rect 38654 44316 38660 44328
rect 38615 44288 38660 44316
rect 28353 44279 28411 44285
rect 28368 44248 28396 44279
rect 38654 44276 38660 44288
rect 38712 44276 38718 44328
rect 38838 44316 38844 44328
rect 38799 44288 38844 44316
rect 38838 44276 38844 44288
rect 38896 44276 38902 44328
rect 40034 44316 40040 44328
rect 39995 44288 40040 44316
rect 40034 44276 40040 44288
rect 40092 44276 40098 44328
rect 42518 44276 42524 44328
rect 42576 44316 42582 44328
rect 43993 44319 44051 44325
rect 43993 44316 44005 44319
rect 42576 44288 44005 44316
rect 42576 44276 42582 44288
rect 43993 44285 44005 44288
rect 44039 44285 44051 44319
rect 43993 44279 44051 44285
rect 6886 44220 28396 44248
rect 29546 44140 29552 44192
rect 29604 44180 29610 44192
rect 31938 44180 31944 44192
rect 29604 44152 31944 44180
rect 29604 44140 29610 44152
rect 31938 44140 31944 44152
rect 31996 44140 32002 44192
rect 47670 44180 47676 44192
rect 47631 44152 47676 44180
rect 47670 44140 47676 44152
rect 47728 44140 47734 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 38838 43976 38844 43988
rect 38799 43948 38844 43976
rect 38838 43936 38844 43948
rect 38896 43936 38902 43988
rect 27341 43843 27399 43849
rect 27341 43809 27353 43843
rect 27387 43840 27399 43843
rect 29641 43843 29699 43849
rect 29641 43840 29653 43843
rect 27387 43812 29653 43840
rect 27387 43809 27399 43812
rect 27341 43803 27399 43809
rect 29641 43809 29653 43812
rect 29687 43809 29699 43843
rect 29641 43803 29699 43809
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 47670 43840 47676 43852
rect 46523 43812 47676 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 47670 43800 47676 43812
rect 47728 43800 47734 43852
rect 48130 43840 48136 43852
rect 48091 43812 48136 43840
rect 48130 43800 48136 43812
rect 48188 43800 48194 43852
rect 26970 43732 26976 43784
rect 27028 43772 27034 43784
rect 27157 43775 27215 43781
rect 27157 43772 27169 43775
rect 27028 43744 27169 43772
rect 27028 43732 27034 43744
rect 27157 43741 27169 43744
rect 27203 43741 27215 43775
rect 29546 43772 29552 43784
rect 29507 43744 29552 43772
rect 27157 43735 27215 43741
rect 29546 43732 29552 43744
rect 29604 43732 29610 43784
rect 38746 43772 38752 43784
rect 38707 43744 38752 43772
rect 38746 43732 38752 43744
rect 38804 43732 38810 43784
rect 45833 43775 45891 43781
rect 45833 43741 45845 43775
rect 45879 43772 45891 43775
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 45879 43744 46305 43772
rect 45879 43741 45891 43744
rect 45833 43735 45891 43741
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 27614 43664 27620 43716
rect 27672 43704 27678 43716
rect 28997 43707 29055 43713
rect 28997 43704 29009 43707
rect 27672 43676 29009 43704
rect 27672 43664 27678 43676
rect 28997 43673 29009 43676
rect 29043 43673 29055 43707
rect 28997 43667 29055 43673
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 27157 43367 27215 43373
rect 27157 43364 27169 43367
rect 6886 43336 27169 43364
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 2130 43188 2136 43240
rect 2188 43228 2194 43240
rect 6886 43228 6914 43336
rect 27157 43333 27169 43336
rect 27203 43333 27215 43367
rect 27157 43327 27215 43333
rect 25590 43256 25596 43308
rect 25648 43296 25654 43308
rect 26237 43299 26295 43305
rect 26237 43296 26249 43299
rect 25648 43268 26249 43296
rect 25648 43256 25654 43268
rect 26237 43265 26249 43268
rect 26283 43265 26295 43299
rect 26237 43259 26295 43265
rect 45186 43256 45192 43308
rect 45244 43296 45250 43308
rect 46293 43299 46351 43305
rect 46293 43296 46305 43299
rect 45244 43268 46305 43296
rect 45244 43256 45250 43268
rect 46293 43265 46305 43268
rect 46339 43265 46351 43299
rect 46934 43296 46940 43308
rect 46895 43268 46940 43296
rect 46293 43259 46351 43265
rect 46934 43256 46940 43268
rect 46992 43256 46998 43308
rect 26970 43228 26976 43240
rect 2188 43200 6914 43228
rect 26931 43200 26976 43228
rect 2188 43188 2194 43200
rect 26970 43188 26976 43200
rect 27028 43188 27034 43240
rect 28810 43228 28816 43240
rect 28771 43200 28816 43228
rect 28810 43188 28816 43200
rect 28868 43188 28874 43240
rect 1578 43092 1584 43104
rect 1539 43064 1584 43092
rect 1578 43052 1584 43064
rect 1636 43052 1642 43104
rect 26329 43095 26387 43101
rect 26329 43061 26341 43095
rect 26375 43092 26387 43095
rect 38654 43092 38660 43104
rect 26375 43064 38660 43092
rect 26375 43061 26387 43064
rect 26329 43055 26387 43061
rect 38654 43052 38660 43064
rect 38712 43052 38718 43104
rect 47762 43092 47768 43104
rect 47723 43064 47768 43092
rect 47762 43052 47768 43064
rect 47820 43052 47826 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46293 42755 46351 42761
rect 46293 42721 46305 42755
rect 46339 42752 46351 42755
rect 47762 42752 47768 42764
rect 46339 42724 47768 42752
rect 46339 42721 46351 42724
rect 46293 42715 46351 42721
rect 47762 42712 47768 42724
rect 47820 42712 47826 42764
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 47670 42616 47676 42628
rect 46523 42588 47676 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 47670 42576 47676 42588
rect 47728 42576 47734 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 47670 42344 47676 42356
rect 47631 42316 47676 42344
rect 47670 42304 47676 42316
rect 47728 42304 47734 42356
rect 27157 42279 27215 42285
rect 27157 42276 27169 42279
rect 6886 42248 27169 42276
rect 1578 42100 1584 42152
rect 1636 42140 1642 42152
rect 6886 42140 6914 42248
rect 27157 42245 27169 42248
rect 27203 42245 27215 42279
rect 27157 42239 27215 42245
rect 45646 42168 45652 42220
rect 45704 42208 45710 42220
rect 46845 42211 46903 42217
rect 46845 42208 46857 42211
rect 45704 42180 46857 42208
rect 45704 42168 45710 42180
rect 46845 42177 46857 42180
rect 46891 42177 46903 42211
rect 46845 42171 46903 42177
rect 47302 42168 47308 42220
rect 47360 42208 47366 42220
rect 47578 42208 47584 42220
rect 47360 42180 47584 42208
rect 47360 42168 47366 42180
rect 47578 42168 47584 42180
rect 47636 42168 47642 42220
rect 1636 42112 6914 42140
rect 1636 42100 1642 42112
rect 26694 42100 26700 42152
rect 26752 42140 26758 42152
rect 26973 42143 27031 42149
rect 26973 42140 26985 42143
rect 26752 42112 26985 42140
rect 26752 42100 26758 42112
rect 26973 42109 26985 42112
rect 27019 42109 27031 42143
rect 28810 42140 28816 42152
rect 28771 42112 28816 42140
rect 26973 42103 27031 42109
rect 28810 42100 28816 42112
rect 28868 42100 28874 42152
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 46474 41964 46480 42016
rect 46532 42004 46538 42016
rect 46937 42007 46995 42013
rect 46937 42004 46949 42007
rect 46532 41976 46949 42004
rect 46532 41964 46538 41976
rect 46937 41973 46949 41976
rect 46983 41973 46995 42007
rect 46937 41967 46995 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46474 41664 46480 41676
rect 46435 41636 46480 41664
rect 46474 41624 46480 41636
rect 46532 41624 46538 41676
rect 46293 41599 46351 41605
rect 46293 41565 46305 41599
rect 46339 41565 46351 41599
rect 46293 41559 46351 41565
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46308 41528 46336 41559
rect 47762 41528 47768 41540
rect 46308 41500 47768 41528
rect 47762 41488 47768 41500
rect 47820 41488 47826 41540
rect 48130 41528 48136 41540
rect 48091 41500 48136 41528
rect 48130 41488 48136 41500
rect 48188 41488 48194 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2133 41259 2191 41265
rect 2133 41256 2145 41259
rect 1636 41228 2145 41256
rect 1636 41216 1642 41228
rect 2133 41225 2145 41228
rect 2179 41225 2191 41259
rect 2133 41219 2191 41225
rect 2041 41123 2099 41129
rect 2041 41089 2053 41123
rect 2087 41120 2099 41123
rect 14090 41120 14096 41132
rect 2087 41092 14096 41120
rect 2087 41089 2099 41092
rect 2041 41083 2099 41089
rect 14090 41080 14096 41092
rect 14148 41080 14154 41132
rect 46198 41120 46204 41132
rect 46159 41092 46204 41120
rect 46198 41080 46204 41092
rect 46256 41080 46262 41132
rect 47762 41120 47768 41132
rect 47723 41092 47768 41120
rect 47762 41080 47768 41092
rect 47820 41080 47826 41132
rect 43806 41012 43812 41064
rect 43864 41052 43870 41064
rect 46477 41055 46535 41061
rect 46477 41052 46489 41055
rect 43864 41024 46489 41052
rect 43864 41012 43870 41024
rect 46477 41021 46489 41024
rect 46523 41021 46535 41055
rect 46477 41015 46535 41021
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 46293 40579 46351 40585
rect 46293 40545 46305 40579
rect 46339 40576 46351 40579
rect 47762 40576 47768 40588
rect 46339 40548 47768 40576
rect 46339 40545 46351 40548
rect 46293 40539 46351 40545
rect 47762 40536 47768 40548
rect 47820 40536 47826 40588
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 2038 40440 2044 40452
rect 1999 40412 2044 40440
rect 2038 40400 2044 40412
rect 2096 40400 2102 40452
rect 45554 40400 45560 40452
rect 45612 40440 45618 40452
rect 46477 40443 46535 40449
rect 46477 40440 46489 40443
rect 45612 40412 46489 40440
rect 45612 40400 45618 40412
rect 46477 40409 46489 40412
rect 46523 40409 46535 40443
rect 48130 40440 48136 40452
rect 48091 40412 48136 40440
rect 46477 40403 46535 40409
rect 48130 40400 48136 40412
rect 48188 40400 48194 40452
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 18966 40100 18972 40112
rect 18927 40072 18972 40100
rect 18966 40060 18972 40072
rect 19024 40100 19030 40112
rect 38194 40100 38200 40112
rect 19024 40072 38200 40100
rect 19024 40060 19030 40072
rect 38194 40060 38200 40072
rect 38252 40060 38258 40112
rect 43806 40100 43812 40112
rect 43732 40072 43812 40100
rect 18414 40032 18420 40044
rect 18375 40004 18420 40032
rect 18414 39992 18420 40004
rect 18472 39992 18478 40044
rect 19150 39992 19156 40044
rect 19208 40032 19214 40044
rect 25314 40032 25320 40044
rect 19208 40004 25320 40032
rect 19208 39992 19214 40004
rect 25314 39992 25320 40004
rect 25372 39992 25378 40044
rect 43625 40035 43683 40041
rect 43625 40001 43637 40035
rect 43671 40032 43683 40035
rect 43732 40032 43760 40072
rect 43806 40060 43812 40072
rect 43864 40060 43870 40112
rect 46014 40100 46020 40112
rect 45848 40072 46020 40100
rect 45848 40041 45876 40072
rect 46014 40060 46020 40072
rect 46072 40060 46078 40112
rect 43671 40004 43760 40032
rect 44361 40035 44419 40041
rect 43671 40001 43683 40004
rect 43625 39995 43683 40001
rect 44361 40001 44373 40035
rect 44407 40032 44419 40035
rect 44913 40035 44971 40041
rect 44913 40032 44925 40035
rect 44407 40004 44925 40032
rect 44407 40001 44419 40004
rect 44361 39995 44419 40001
rect 44913 40001 44925 40004
rect 44959 40001 44971 40035
rect 44913 39995 44971 40001
rect 45833 40035 45891 40041
rect 45833 40001 45845 40035
rect 45879 40001 45891 40035
rect 47762 40032 47768 40044
rect 47723 40004 47768 40032
rect 45833 39995 45891 40001
rect 47762 39992 47768 40004
rect 47820 39992 47826 40044
rect 43714 39964 43720 39976
rect 43675 39936 43720 39964
rect 43714 39924 43720 39936
rect 43772 39924 43778 39976
rect 26970 39856 26976 39908
rect 27028 39896 27034 39908
rect 46109 39899 46167 39905
rect 46109 39896 46121 39899
rect 27028 39868 46121 39896
rect 27028 39856 27034 39868
rect 46109 39865 46121 39868
rect 46155 39865 46167 39899
rect 46109 39859 46167 39865
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 18322 39448 18328 39500
rect 18380 39488 18386 39500
rect 18601 39491 18659 39497
rect 18601 39488 18613 39491
rect 18380 39460 18613 39488
rect 18380 39448 18386 39460
rect 18601 39457 18613 39460
rect 18647 39488 18659 39491
rect 22738 39488 22744 39500
rect 18647 39460 22094 39488
rect 22699 39460 22744 39488
rect 18647 39457 18659 39460
rect 18601 39451 18659 39457
rect 17037 39423 17095 39429
rect 17037 39389 17049 39423
rect 17083 39420 17095 39423
rect 18049 39423 18107 39429
rect 18049 39420 18061 39423
rect 17083 39392 18061 39420
rect 17083 39389 17095 39392
rect 17037 39383 17095 39389
rect 18049 39389 18061 39392
rect 18095 39420 18107 39423
rect 18414 39420 18420 39432
rect 18095 39392 18420 39420
rect 18095 39389 18107 39392
rect 18049 39383 18107 39389
rect 18414 39380 18420 39392
rect 18472 39420 18478 39432
rect 19245 39423 19303 39429
rect 19245 39420 19257 39423
rect 18472 39392 19257 39420
rect 18472 39380 18478 39392
rect 19245 39389 19257 39392
rect 19291 39389 19303 39423
rect 22066 39420 22094 39460
rect 22738 39448 22744 39460
rect 22796 39448 22802 39500
rect 46293 39491 46351 39497
rect 46293 39457 46305 39491
rect 46339 39488 46351 39491
rect 47854 39488 47860 39500
rect 46339 39460 47860 39488
rect 46339 39457 46351 39460
rect 46293 39451 46351 39457
rect 47854 39448 47860 39460
rect 47912 39448 47918 39500
rect 38746 39420 38752 39432
rect 22066 39392 38752 39420
rect 19245 39383 19303 39389
rect 38746 39380 38752 39392
rect 38804 39420 38810 39432
rect 39942 39420 39948 39432
rect 38804 39392 39948 39420
rect 38804 39380 38810 39392
rect 39942 39380 39948 39392
rect 40000 39380 40006 39432
rect 16666 39312 16672 39364
rect 16724 39352 16730 39364
rect 17313 39355 17371 39361
rect 17313 39352 17325 39355
rect 16724 39324 17325 39352
rect 16724 39312 16730 39324
rect 17313 39321 17325 39324
rect 17359 39352 17371 39355
rect 17586 39352 17592 39364
rect 17359 39324 17592 39352
rect 17359 39321 17371 39324
rect 17313 39315 17371 39321
rect 17586 39312 17592 39324
rect 17644 39312 17650 39364
rect 20073 39355 20131 39361
rect 20073 39321 20085 39355
rect 20119 39352 20131 39355
rect 20622 39352 20628 39364
rect 20119 39324 20628 39352
rect 20119 39321 20131 39324
rect 20073 39315 20131 39321
rect 20622 39312 20628 39324
rect 20680 39352 20686 39364
rect 42058 39352 42064 39364
rect 20680 39324 42064 39352
rect 20680 39312 20686 39324
rect 42058 39312 42064 39324
rect 42116 39312 42122 39364
rect 46477 39355 46535 39361
rect 46477 39321 46489 39355
rect 46523 39352 46535 39355
rect 47670 39352 47676 39364
rect 46523 39324 47676 39352
rect 46523 39321 46535 39324
rect 46477 39315 46535 39321
rect 47670 39312 47676 39324
rect 47728 39312 47734 39364
rect 48130 39352 48136 39364
rect 48091 39324 48136 39352
rect 48130 39312 48136 39324
rect 48188 39312 48194 39364
rect 22186 39284 22192 39296
rect 22147 39256 22192 39284
rect 22186 39244 22192 39256
rect 22244 39244 22250 39296
rect 22462 39244 22468 39296
rect 22520 39284 22526 39296
rect 22557 39287 22615 39293
rect 22557 39284 22569 39287
rect 22520 39256 22569 39284
rect 22520 39244 22526 39256
rect 22557 39253 22569 39256
rect 22603 39253 22615 39287
rect 22557 39247 22615 39253
rect 22646 39244 22652 39296
rect 22704 39284 22710 39296
rect 22704 39256 22749 39284
rect 22704 39244 22710 39256
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 22462 39040 22468 39092
rect 22520 39080 22526 39092
rect 23569 39083 23627 39089
rect 23569 39080 23581 39083
rect 22520 39052 23581 39080
rect 22520 39040 22526 39052
rect 23569 39049 23581 39052
rect 23615 39049 23627 39083
rect 47670 39080 47676 39092
rect 47631 39052 47676 39080
rect 23569 39043 23627 39049
rect 47670 39040 47676 39052
rect 47728 39040 47734 39092
rect 22554 38972 22560 39024
rect 22612 38972 22618 39024
rect 18414 38944 18420 38956
rect 18375 38916 18420 38944
rect 18414 38904 18420 38916
rect 18472 38904 18478 38956
rect 25777 38947 25835 38953
rect 25777 38913 25789 38947
rect 25823 38944 25835 38947
rect 26970 38944 26976 38956
rect 25823 38916 26976 38944
rect 25823 38913 25835 38916
rect 25777 38907 25835 38913
rect 26970 38904 26976 38916
rect 27028 38904 27034 38956
rect 30190 38904 30196 38956
rect 30248 38944 30254 38956
rect 30285 38947 30343 38953
rect 30285 38944 30297 38947
rect 30248 38916 30297 38944
rect 30248 38904 30254 38916
rect 30285 38913 30297 38916
rect 30331 38913 30343 38947
rect 45646 38944 45652 38956
rect 45607 38916 45652 38944
rect 30285 38907 30343 38913
rect 45646 38904 45652 38916
rect 45704 38904 45710 38956
rect 45830 38944 45836 38956
rect 45791 38916 45836 38944
rect 45830 38904 45836 38916
rect 45888 38904 45894 38956
rect 46382 38944 46388 38956
rect 46343 38916 46388 38944
rect 46382 38904 46388 38916
rect 46440 38904 46446 38956
rect 47581 38947 47639 38953
rect 47581 38913 47593 38947
rect 47627 38944 47639 38947
rect 47670 38944 47676 38956
rect 47627 38916 47676 38944
rect 47627 38913 47639 38916
rect 47581 38907 47639 38913
rect 47670 38904 47676 38916
rect 47728 38904 47734 38956
rect 19150 38876 19156 38888
rect 19111 38848 19156 38876
rect 19150 38836 19156 38848
rect 19208 38836 19214 38888
rect 21818 38876 21824 38888
rect 21779 38848 21824 38876
rect 21818 38836 21824 38848
rect 21876 38836 21882 38888
rect 22094 38836 22100 38888
rect 22152 38876 22158 38888
rect 46842 38876 46848 38888
rect 22152 38848 22197 38876
rect 46803 38848 46848 38876
rect 22152 38836 22158 38848
rect 46842 38836 46848 38848
rect 46900 38836 46906 38888
rect 24854 38700 24860 38752
rect 24912 38740 24918 38752
rect 25593 38743 25651 38749
rect 25593 38740 25605 38743
rect 24912 38712 25605 38740
rect 24912 38700 24918 38712
rect 25593 38709 25605 38712
rect 25639 38709 25651 38743
rect 25593 38703 25651 38709
rect 30469 38743 30527 38749
rect 30469 38709 30481 38743
rect 30515 38740 30527 38743
rect 45554 38740 45560 38752
rect 30515 38712 45560 38740
rect 30515 38709 30527 38712
rect 30469 38703 30527 38709
rect 45554 38700 45560 38712
rect 45612 38700 45618 38752
rect 45649 38743 45707 38749
rect 45649 38709 45661 38743
rect 45695 38740 45707 38743
rect 46106 38740 46112 38752
rect 45695 38712 46112 38740
rect 45695 38709 45707 38712
rect 45649 38703 45707 38709
rect 46106 38700 46112 38712
rect 46164 38700 46170 38752
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 18325 38539 18383 38545
rect 18325 38505 18337 38539
rect 18371 38536 18383 38539
rect 18414 38536 18420 38548
rect 18371 38508 18420 38536
rect 18371 38505 18383 38508
rect 18325 38499 18383 38505
rect 18414 38496 18420 38508
rect 18472 38496 18478 38548
rect 22646 38496 22652 38548
rect 22704 38536 22710 38548
rect 22833 38539 22891 38545
rect 22833 38536 22845 38539
rect 22704 38508 22845 38536
rect 22704 38496 22710 38508
rect 22833 38505 22845 38508
rect 22879 38505 22891 38539
rect 22833 38499 22891 38505
rect 24486 38496 24492 38548
rect 24544 38536 24550 38548
rect 26970 38536 26976 38548
rect 24544 38508 25912 38536
rect 26931 38508 26976 38536
rect 24544 38496 24550 38508
rect 19245 38471 19303 38477
rect 19245 38437 19257 38471
rect 19291 38437 19303 38471
rect 19245 38431 19303 38437
rect 19444 38440 21036 38468
rect 19260 38400 19288 38431
rect 17604 38372 19288 38400
rect 17604 38341 17632 38372
rect 17589 38335 17647 38341
rect 17589 38301 17601 38335
rect 17635 38301 17647 38335
rect 17589 38295 17647 38301
rect 17957 38335 18015 38341
rect 17957 38301 17969 38335
rect 18003 38332 18015 38335
rect 18509 38335 18567 38341
rect 18509 38332 18521 38335
rect 18003 38304 18521 38332
rect 18003 38301 18015 38304
rect 17957 38295 18015 38301
rect 18509 38301 18521 38304
rect 18555 38332 18567 38335
rect 19444 38332 19472 38440
rect 19889 38403 19947 38409
rect 19889 38369 19901 38403
rect 19935 38400 19947 38403
rect 20898 38400 20904 38412
rect 19935 38372 20904 38400
rect 19935 38369 19947 38372
rect 19889 38363 19947 38369
rect 20898 38360 20904 38372
rect 20956 38360 20962 38412
rect 21008 38400 21036 38440
rect 21082 38428 21088 38480
rect 21140 38468 21146 38480
rect 21818 38468 21824 38480
rect 21140 38440 21824 38468
rect 21140 38428 21146 38440
rect 21818 38428 21824 38440
rect 21876 38468 21882 38480
rect 21876 38440 24624 38468
rect 21876 38428 21882 38440
rect 23474 38400 23480 38412
rect 21008 38372 23336 38400
rect 23435 38372 23480 38400
rect 18555 38304 19472 38332
rect 19613 38335 19671 38341
rect 18555 38301 18567 38304
rect 18509 38295 18567 38301
rect 19613 38301 19625 38335
rect 19659 38332 19671 38335
rect 19978 38332 19984 38344
rect 19659 38304 19984 38332
rect 19659 38301 19671 38304
rect 19613 38295 19671 38301
rect 19978 38292 19984 38304
rect 20036 38292 20042 38344
rect 20533 38335 20591 38341
rect 20533 38301 20545 38335
rect 20579 38332 20591 38335
rect 21174 38332 21180 38344
rect 20579 38304 21180 38332
rect 20579 38301 20591 38304
rect 20533 38295 20591 38301
rect 21174 38292 21180 38304
rect 21232 38292 21238 38344
rect 22005 38335 22063 38341
rect 22005 38301 22017 38335
rect 22051 38332 22063 38335
rect 22186 38332 22192 38344
rect 22051 38304 22192 38332
rect 22051 38301 22063 38304
rect 22005 38295 22063 38301
rect 22186 38292 22192 38304
rect 22244 38292 22250 38344
rect 23308 38332 23336 38372
rect 23474 38360 23480 38372
rect 23532 38360 23538 38412
rect 24596 38409 24624 38440
rect 24581 38403 24639 38409
rect 24581 38369 24593 38403
rect 24627 38400 24639 38403
rect 25406 38400 25412 38412
rect 24627 38372 25412 38400
rect 24627 38369 24639 38372
rect 24581 38363 24639 38369
rect 25406 38360 25412 38372
rect 25464 38360 25470 38412
rect 25884 38400 25912 38508
rect 26970 38496 26976 38508
rect 27028 38496 27034 38548
rect 46566 38536 46572 38548
rect 35866 38508 46572 38536
rect 27525 38403 27583 38409
rect 27525 38400 27537 38403
rect 25884 38372 27537 38400
rect 27525 38369 27537 38372
rect 27571 38369 27583 38403
rect 27525 38363 27583 38369
rect 26697 38335 26755 38341
rect 23308 38304 23520 38332
rect 11974 38224 11980 38276
rect 12032 38264 12038 38276
rect 23201 38267 23259 38273
rect 23201 38264 23213 38267
rect 12032 38236 23213 38264
rect 12032 38224 12038 38236
rect 23201 38233 23213 38236
rect 23247 38233 23259 38267
rect 23201 38227 23259 38233
rect 17126 38156 17132 38208
rect 17184 38196 17190 38208
rect 17405 38199 17463 38205
rect 17405 38196 17417 38199
rect 17184 38168 17417 38196
rect 17184 38156 17190 38168
rect 17405 38165 17417 38168
rect 17451 38165 17463 38199
rect 17405 38159 17463 38165
rect 18690 38156 18696 38208
rect 18748 38196 18754 38208
rect 19705 38199 19763 38205
rect 19705 38196 19717 38199
rect 18748 38168 19717 38196
rect 18748 38156 18754 38168
rect 19705 38165 19717 38168
rect 19751 38165 19763 38199
rect 19705 38159 19763 38165
rect 20530 38156 20536 38208
rect 20588 38196 20594 38208
rect 20625 38199 20683 38205
rect 20625 38196 20637 38199
rect 20588 38168 20637 38196
rect 20588 38156 20594 38168
rect 20625 38165 20637 38168
rect 20671 38165 20683 38199
rect 20625 38159 20683 38165
rect 21821 38199 21879 38205
rect 21821 38165 21833 38199
rect 21867 38196 21879 38199
rect 22094 38196 22100 38208
rect 21867 38168 22100 38196
rect 21867 38165 21879 38168
rect 21821 38159 21879 38165
rect 22094 38156 22100 38168
rect 22152 38156 22158 38208
rect 23290 38156 23296 38208
rect 23348 38196 23354 38208
rect 23492 38196 23520 38304
rect 26697 38301 26709 38335
rect 26743 38332 26755 38335
rect 27341 38335 27399 38341
rect 27341 38332 27353 38335
rect 26743 38304 27353 38332
rect 26743 38301 26755 38304
rect 26697 38295 26755 38301
rect 27341 38301 27353 38304
rect 27387 38332 27399 38335
rect 35866 38332 35894 38508
rect 46566 38496 46572 38508
rect 46624 38496 46630 38548
rect 45830 38468 45836 38480
rect 45112 38440 45836 38468
rect 45112 38409 45140 38440
rect 45830 38428 45836 38440
rect 45888 38428 45894 38480
rect 45097 38403 45155 38409
rect 45097 38369 45109 38403
rect 45143 38369 45155 38403
rect 45465 38403 45523 38409
rect 45465 38400 45477 38403
rect 45097 38363 45155 38369
rect 45204 38372 45477 38400
rect 27387 38304 35894 38332
rect 44269 38335 44327 38341
rect 27387 38301 27399 38304
rect 27341 38295 27399 38301
rect 44269 38301 44281 38335
rect 44315 38301 44327 38335
rect 44269 38295 44327 38301
rect 44453 38335 44511 38341
rect 44453 38301 44465 38335
rect 44499 38332 44511 38335
rect 45204 38332 45232 38372
rect 45465 38369 45477 38372
rect 45511 38369 45523 38403
rect 45465 38363 45523 38369
rect 44499 38304 45232 38332
rect 45281 38335 45339 38341
rect 44499 38301 44511 38304
rect 44453 38295 44511 38301
rect 45281 38301 45293 38335
rect 45327 38332 45339 38335
rect 45646 38332 45652 38344
rect 45327 38304 45652 38332
rect 45327 38301 45339 38304
rect 45281 38295 45339 38301
rect 24854 38264 24860 38276
rect 24815 38236 24860 38264
rect 24854 38224 24860 38236
rect 24912 38224 24918 38276
rect 25314 38224 25320 38276
rect 25372 38224 25378 38276
rect 26142 38196 26148 38208
rect 23348 38168 23393 38196
rect 23492 38168 26148 38196
rect 23348 38156 23354 38168
rect 26142 38156 26148 38168
rect 26200 38156 26206 38208
rect 26326 38196 26332 38208
rect 26287 38168 26332 38196
rect 26326 38156 26332 38168
rect 26384 38156 26390 38208
rect 26418 38156 26424 38208
rect 26476 38196 26482 38208
rect 27433 38199 27491 38205
rect 27433 38196 27445 38199
rect 26476 38168 27445 38196
rect 26476 38156 26482 38168
rect 27433 38165 27445 38168
rect 27479 38165 27491 38199
rect 44284 38196 44312 38295
rect 45646 38292 45652 38304
rect 45704 38292 45710 38344
rect 45922 38292 45928 38344
rect 45980 38332 45986 38344
rect 46017 38335 46075 38341
rect 46017 38332 46029 38335
rect 45980 38304 46029 38332
rect 45980 38292 45986 38304
rect 46017 38301 46029 38304
rect 46063 38301 46075 38335
rect 46017 38295 46075 38301
rect 46385 38335 46443 38341
rect 46385 38301 46397 38335
rect 46431 38301 46443 38335
rect 46385 38295 46443 38301
rect 44361 38267 44419 38273
rect 44361 38233 44373 38267
rect 44407 38264 44419 38267
rect 46400 38264 46428 38295
rect 47854 38264 47860 38276
rect 44407 38236 46428 38264
rect 47815 38236 47860 38264
rect 44407 38233 44419 38236
rect 44361 38227 44419 38233
rect 47854 38224 47860 38236
rect 47912 38224 47918 38276
rect 46106 38196 46112 38208
rect 44284 38168 46112 38196
rect 27433 38159 27491 38165
rect 46106 38156 46112 38168
rect 46164 38156 46170 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 22005 37995 22063 38001
rect 22005 37961 22017 37995
rect 22051 37992 22063 37995
rect 22554 37992 22560 38004
rect 22051 37964 22560 37992
rect 22051 37961 22063 37964
rect 22005 37955 22063 37961
rect 22554 37952 22560 37964
rect 22612 37952 22618 38004
rect 23109 37995 23167 38001
rect 23109 37961 23121 37995
rect 23155 37992 23167 37995
rect 23290 37992 23296 38004
rect 23155 37964 23296 37992
rect 23155 37961 23167 37964
rect 23109 37955 23167 37961
rect 23290 37952 23296 37964
rect 23348 37952 23354 38004
rect 24486 37992 24492 38004
rect 24447 37964 24492 37992
rect 24486 37952 24492 37964
rect 24544 37952 24550 38004
rect 25225 37995 25283 38001
rect 25225 37961 25237 37995
rect 25271 37992 25283 37995
rect 25314 37992 25320 38004
rect 25271 37964 25320 37992
rect 25271 37961 25283 37964
rect 25225 37955 25283 37961
rect 25314 37952 25320 37964
rect 25372 37952 25378 38004
rect 26142 37952 26148 38004
rect 26200 37992 26206 38004
rect 46014 37992 46020 38004
rect 26200 37964 35894 37992
rect 45975 37964 46020 37992
rect 26200 37952 26206 37964
rect 17126 37924 17132 37936
rect 17087 37896 17132 37924
rect 17126 37884 17132 37896
rect 17184 37884 17190 37936
rect 18138 37884 18144 37936
rect 18196 37884 18202 37936
rect 20530 37884 20536 37936
rect 20588 37884 20594 37936
rect 21174 37816 21180 37868
rect 21232 37856 21238 37868
rect 21913 37859 21971 37865
rect 21913 37856 21925 37859
rect 21232 37828 21925 37856
rect 21232 37816 21238 37828
rect 21913 37825 21925 37828
rect 21959 37825 21971 37859
rect 21913 37819 21971 37825
rect 22462 37816 22468 37868
rect 22520 37856 22526 37868
rect 22646 37856 22652 37868
rect 22520 37828 22652 37856
rect 22520 37816 22526 37828
rect 22646 37816 22652 37828
rect 22704 37856 22710 37868
rect 22741 37859 22799 37865
rect 22741 37856 22753 37859
rect 22704 37828 22753 37856
rect 22704 37816 22710 37828
rect 22741 37825 22753 37828
rect 22787 37825 22799 37859
rect 22741 37819 22799 37825
rect 23474 37816 23480 37868
rect 23532 37856 23538 37868
rect 24213 37859 24271 37865
rect 24213 37856 24225 37859
rect 23532 37828 24225 37856
rect 23532 37816 23538 37828
rect 24213 37825 24225 37828
rect 24259 37856 24271 37859
rect 24578 37856 24584 37868
rect 24259 37828 24584 37856
rect 24259 37825 24271 37828
rect 24213 37819 24271 37825
rect 24578 37816 24584 37828
rect 24636 37816 24642 37868
rect 24670 37816 24676 37868
rect 24728 37856 24734 37868
rect 25133 37859 25191 37865
rect 25133 37856 25145 37859
rect 24728 37828 25145 37856
rect 24728 37816 24734 37828
rect 25133 37825 25145 37828
rect 25179 37825 25191 37859
rect 25133 37819 25191 37825
rect 26053 37859 26111 37865
rect 26053 37825 26065 37859
rect 26099 37856 26111 37859
rect 26326 37856 26332 37868
rect 26099 37828 26332 37856
rect 26099 37825 26111 37828
rect 26053 37819 26111 37825
rect 26326 37816 26332 37828
rect 26384 37856 26390 37868
rect 26384 37828 26648 37856
rect 26384 37816 26390 37828
rect 16298 37748 16304 37800
rect 16356 37788 16362 37800
rect 16853 37791 16911 37797
rect 16853 37788 16865 37791
rect 16356 37760 16865 37788
rect 16356 37748 16362 37760
rect 16853 37757 16865 37760
rect 16899 37788 16911 37791
rect 19521 37791 19579 37797
rect 19521 37788 19533 37791
rect 16899 37760 19533 37788
rect 16899 37757 16911 37760
rect 16853 37751 16911 37757
rect 19521 37757 19533 37760
rect 19567 37757 19579 37791
rect 19521 37751 19579 37757
rect 19797 37791 19855 37797
rect 19797 37757 19809 37791
rect 19843 37788 19855 37791
rect 20530 37788 20536 37800
rect 19843 37760 20536 37788
rect 19843 37757 19855 37760
rect 19797 37751 19855 37757
rect 18598 37612 18604 37664
rect 18656 37652 18662 37664
rect 19536 37652 19564 37751
rect 20530 37748 20536 37760
rect 20588 37748 20594 37800
rect 22094 37748 22100 37800
rect 22152 37788 22158 37800
rect 22833 37791 22891 37797
rect 22833 37788 22845 37791
rect 22152 37760 22845 37788
rect 22152 37748 22158 37760
rect 22833 37757 22845 37760
rect 22879 37788 22891 37791
rect 26145 37791 26203 37797
rect 22879 37760 25544 37788
rect 22879 37757 22891 37760
rect 22833 37751 22891 37757
rect 20898 37680 20904 37732
rect 20956 37720 20962 37732
rect 24302 37720 24308 37732
rect 20956 37692 24308 37720
rect 20956 37680 20962 37692
rect 24302 37680 24308 37692
rect 24360 37720 24366 37732
rect 24486 37720 24492 37732
rect 24360 37692 24492 37720
rect 24360 37680 24366 37692
rect 24486 37680 24492 37692
rect 24544 37680 24550 37732
rect 20806 37652 20812 37664
rect 18656 37624 18701 37652
rect 19536 37624 20812 37652
rect 18656 37612 18662 37624
rect 20806 37612 20812 37624
rect 20864 37652 20870 37664
rect 21082 37652 21088 37664
rect 20864 37624 21088 37652
rect 20864 37612 20870 37624
rect 21082 37612 21088 37624
rect 21140 37612 21146 37664
rect 21266 37652 21272 37664
rect 21227 37624 21272 37652
rect 21266 37612 21272 37624
rect 21324 37612 21330 37664
rect 25516 37652 25544 37760
rect 26145 37757 26157 37791
rect 26191 37757 26203 37791
rect 26418 37788 26424 37800
rect 26379 37760 26424 37788
rect 26145 37751 26203 37757
rect 26160 37720 26188 37751
rect 26418 37748 26424 37760
rect 26476 37748 26482 37800
rect 26620 37788 26648 37828
rect 26878 37816 26884 37868
rect 26936 37856 26942 37868
rect 26973 37859 27031 37865
rect 26973 37856 26985 37859
rect 26936 37828 26985 37856
rect 26936 37816 26942 37828
rect 26973 37825 26985 37828
rect 27019 37825 27031 37859
rect 26973 37819 27031 37825
rect 29546 37816 29552 37868
rect 29604 37816 29610 37868
rect 27522 37788 27528 37800
rect 26620 37760 27528 37788
rect 27522 37748 27528 37760
rect 27580 37748 27586 37800
rect 28166 37788 28172 37800
rect 28127 37760 28172 37788
rect 28166 37748 28172 37760
rect 28224 37748 28230 37800
rect 28445 37791 28503 37797
rect 28445 37757 28457 37791
rect 28491 37788 28503 37791
rect 28902 37788 28908 37800
rect 28491 37760 28908 37788
rect 28491 37757 28503 37760
rect 28445 37751 28503 37757
rect 28902 37748 28908 37760
rect 28960 37748 28966 37800
rect 26326 37720 26332 37732
rect 26160 37692 26332 37720
rect 26326 37680 26332 37692
rect 26384 37680 26390 37732
rect 35866 37720 35894 37964
rect 46014 37952 46020 37964
rect 46072 37952 46078 38004
rect 39942 37884 39948 37936
rect 40000 37924 40006 37936
rect 45554 37924 45560 37936
rect 40000 37896 45560 37924
rect 40000 37884 40006 37896
rect 45554 37884 45560 37896
rect 45612 37924 45618 37936
rect 45612 37896 46704 37924
rect 45612 37884 45618 37896
rect 45738 37856 45744 37868
rect 45699 37828 45744 37856
rect 45738 37816 45744 37828
rect 45796 37816 45802 37868
rect 46106 37856 46112 37868
rect 46067 37828 46112 37856
rect 46106 37816 46112 37828
rect 46164 37816 46170 37868
rect 46676 37865 46704 37896
rect 46661 37859 46719 37865
rect 46661 37825 46673 37859
rect 46707 37825 46719 37859
rect 46661 37819 46719 37825
rect 45557 37791 45615 37797
rect 45557 37757 45569 37791
rect 45603 37788 45615 37791
rect 45922 37788 45928 37800
rect 45603 37760 45928 37788
rect 45603 37757 45615 37760
rect 45557 37751 45615 37757
rect 45922 37748 45928 37760
rect 45980 37748 45986 37800
rect 46014 37720 46020 37732
rect 35866 37692 46020 37720
rect 46014 37680 46020 37692
rect 46072 37680 46078 37732
rect 26142 37652 26148 37664
rect 25516 37624 26148 37652
rect 26142 37612 26148 37624
rect 26200 37612 26206 37664
rect 27154 37652 27160 37664
rect 27067 37624 27160 37652
rect 27154 37612 27160 37624
rect 27212 37652 27218 37664
rect 28258 37652 28264 37664
rect 27212 37624 28264 37652
rect 27212 37612 27218 37624
rect 28258 37612 28264 37624
rect 28316 37612 28322 37664
rect 29914 37652 29920 37664
rect 29875 37624 29920 37652
rect 29914 37612 29920 37624
rect 29972 37612 29978 37664
rect 46474 37612 46480 37664
rect 46532 37652 46538 37664
rect 46753 37655 46811 37661
rect 46753 37652 46765 37655
rect 46532 37624 46765 37652
rect 46532 37612 46538 37624
rect 46753 37621 46765 37624
rect 46799 37621 46811 37655
rect 47762 37652 47768 37664
rect 47723 37624 47768 37652
rect 46753 37615 46811 37621
rect 47762 37612 47768 37624
rect 47820 37612 47826 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 9490 37408 9496 37460
rect 9548 37448 9554 37460
rect 28902 37448 28908 37460
rect 9548 37420 28580 37448
rect 28863 37420 28908 37448
rect 9548 37408 9554 37420
rect 2038 37340 2044 37392
rect 2096 37380 2102 37392
rect 18690 37380 18696 37392
rect 2096 37352 18368 37380
rect 18651 37352 18696 37380
rect 2096 37340 2102 37352
rect 18230 37312 18236 37324
rect 18191 37284 18236 37312
rect 18230 37272 18236 37284
rect 18288 37272 18294 37324
rect 18340 37312 18368 37352
rect 18690 37340 18696 37352
rect 18748 37340 18754 37392
rect 19978 37380 19984 37392
rect 19306 37352 19984 37380
rect 19306 37312 19334 37352
rect 19978 37340 19984 37352
rect 20036 37340 20042 37392
rect 20530 37380 20536 37392
rect 20491 37352 20536 37380
rect 20530 37340 20536 37352
rect 20588 37340 20594 37392
rect 22094 37380 22100 37392
rect 22055 37352 22100 37380
rect 22094 37340 22100 37352
rect 22152 37340 22158 37392
rect 22646 37380 22652 37392
rect 22204 37352 22652 37380
rect 18340 37284 19334 37312
rect 20073 37315 20131 37321
rect 20073 37281 20085 37315
rect 20119 37312 20131 37315
rect 21266 37312 21272 37324
rect 20119 37284 21272 37312
rect 20119 37281 20131 37284
rect 20073 37275 20131 37281
rect 21266 37272 21272 37284
rect 21324 37312 21330 37324
rect 22204 37321 22232 37352
rect 22646 37340 22652 37352
rect 22704 37340 22710 37392
rect 22189 37315 22247 37321
rect 21324 37284 21956 37312
rect 21324 37272 21330 37284
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 2041 37247 2099 37253
rect 2041 37244 2053 37247
rect 1820 37216 2053 37244
rect 1820 37204 1826 37216
rect 2041 37213 2053 37216
rect 2087 37213 2099 37247
rect 2041 37207 2099 37213
rect 18325 37247 18383 37253
rect 18325 37213 18337 37247
rect 18371 37244 18383 37247
rect 18506 37244 18512 37256
rect 18371 37216 18512 37244
rect 18371 37213 18383 37216
rect 18325 37207 18383 37213
rect 18506 37204 18512 37216
rect 18564 37204 18570 37256
rect 19794 37244 19800 37256
rect 19755 37216 19800 37244
rect 19794 37204 19800 37216
rect 19852 37204 19858 37256
rect 19981 37247 20039 37253
rect 19981 37213 19993 37247
rect 20027 37213 20039 37247
rect 19981 37207 20039 37213
rect 19334 37136 19340 37188
rect 19392 37176 19398 37188
rect 19996 37176 20024 37207
rect 20162 37204 20168 37256
rect 20220 37244 20226 37256
rect 20220 37216 20265 37244
rect 20220 37204 20226 37216
rect 20346 37204 20352 37256
rect 20404 37244 20410 37256
rect 21928 37253 21956 37284
rect 22189 37281 22201 37315
rect 22235 37281 22247 37315
rect 22189 37275 22247 37281
rect 22278 37272 22284 37324
rect 22336 37312 22342 37324
rect 27154 37312 27160 37324
rect 22336 37284 27160 37312
rect 22336 37272 22342 37284
rect 27154 37272 27160 37284
rect 27212 37272 27218 37324
rect 28552 37321 28580 37420
rect 28902 37408 28908 37420
rect 28960 37408 28966 37460
rect 29546 37408 29552 37460
rect 29604 37448 29610 37460
rect 29641 37451 29699 37457
rect 29641 37448 29653 37451
rect 29604 37420 29653 37448
rect 29604 37408 29610 37420
rect 29641 37417 29653 37420
rect 29687 37417 29699 37451
rect 45738 37448 45744 37460
rect 45699 37420 45744 37448
rect 29641 37411 29699 37417
rect 45738 37408 45744 37420
rect 45796 37408 45802 37460
rect 46014 37340 46020 37392
rect 46072 37380 46078 37392
rect 46842 37380 46848 37392
rect 46072 37352 46848 37380
rect 46072 37340 46078 37352
rect 46842 37340 46848 37352
rect 46900 37340 46906 37392
rect 28537 37315 28595 37321
rect 28537 37281 28549 37315
rect 28583 37281 28595 37315
rect 29730 37312 29736 37324
rect 28537 37275 28595 37281
rect 28644 37284 29736 37312
rect 21913 37247 21971 37253
rect 20404 37216 20449 37244
rect 20404 37204 20410 37216
rect 21913 37213 21925 37247
rect 21959 37244 21971 37247
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 21959 37216 22845 37244
rect 21959 37213 21971 37216
rect 21913 37207 21971 37213
rect 22833 37213 22845 37216
rect 22879 37213 22891 37247
rect 22833 37207 22891 37213
rect 28169 37247 28227 37253
rect 28169 37213 28181 37247
rect 28215 37213 28227 37247
rect 28350 37244 28356 37256
rect 28311 37216 28356 37244
rect 28169 37207 28227 37213
rect 22278 37176 22284 37188
rect 19392 37148 22284 37176
rect 19392 37136 19398 37148
rect 22278 37136 22284 37148
rect 22336 37136 22342 37188
rect 22646 37176 22652 37188
rect 22607 37148 22652 37176
rect 22646 37136 22652 37148
rect 22704 37136 22710 37188
rect 22738 37136 22744 37188
rect 22796 37176 22802 37188
rect 26510 37176 26516 37188
rect 22796 37148 26516 37176
rect 22796 37136 22802 37148
rect 26510 37136 26516 37148
rect 26568 37176 26574 37188
rect 26878 37176 26884 37188
rect 26568 37148 26884 37176
rect 26568 37136 26574 37148
rect 26878 37136 26884 37148
rect 26936 37136 26942 37188
rect 28184 37176 28212 37207
rect 28350 37204 28356 37216
rect 28408 37204 28414 37256
rect 28445 37247 28503 37253
rect 28445 37213 28457 37247
rect 28491 37244 28503 37247
rect 28644 37244 28672 37284
rect 29730 37272 29736 37284
rect 29788 37312 29794 37324
rect 29914 37312 29920 37324
rect 29788 37284 29920 37312
rect 29788 37272 29794 37284
rect 29914 37272 29920 37284
rect 29972 37272 29978 37324
rect 45554 37272 45560 37324
rect 45612 37312 45618 37324
rect 45738 37312 45744 37324
rect 45612 37284 45744 37312
rect 45612 37272 45618 37284
rect 45738 37272 45744 37284
rect 45796 37272 45802 37324
rect 46474 37312 46480 37324
rect 46435 37284 46480 37312
rect 46474 37272 46480 37284
rect 46532 37272 46538 37324
rect 48130 37312 48136 37324
rect 48091 37284 48136 37312
rect 48130 37272 48136 37284
rect 48188 37272 48194 37324
rect 28491 37216 28672 37244
rect 28491 37213 28503 37216
rect 28445 37207 28503 37213
rect 28718 37204 28724 37256
rect 28776 37244 28782 37256
rect 29549 37247 29607 37253
rect 29549 37244 29561 37247
rect 28776 37216 28821 37244
rect 29288 37216 29561 37244
rect 28776 37204 28782 37216
rect 29178 37176 29184 37188
rect 28184 37148 29184 37176
rect 29178 37136 29184 37148
rect 29236 37136 29242 37188
rect 21726 37108 21732 37120
rect 21687 37080 21732 37108
rect 21726 37068 21732 37080
rect 21784 37068 21790 37120
rect 23017 37111 23075 37117
rect 23017 37077 23029 37111
rect 23063 37108 23075 37111
rect 23198 37108 23204 37120
rect 23063 37080 23204 37108
rect 23063 37077 23075 37080
rect 23017 37071 23075 37077
rect 23198 37068 23204 37080
rect 23256 37068 23262 37120
rect 26970 37068 26976 37120
rect 27028 37108 27034 37120
rect 29288 37108 29316 37216
rect 29549 37213 29561 37216
rect 29595 37244 29607 37247
rect 30742 37244 30748 37256
rect 29595 37216 30748 37244
rect 29595 37213 29607 37216
rect 29549 37207 29607 37213
rect 30742 37204 30748 37216
rect 30800 37204 30806 37256
rect 45646 37244 45652 37256
rect 45607 37216 45652 37244
rect 45646 37204 45652 37216
rect 45704 37204 45710 37256
rect 45830 37244 45836 37256
rect 45791 37216 45836 37244
rect 45830 37204 45836 37216
rect 45888 37204 45894 37256
rect 46293 37247 46351 37253
rect 46293 37213 46305 37247
rect 46339 37213 46351 37247
rect 46293 37207 46351 37213
rect 46308 37176 46336 37207
rect 47762 37176 47768 37188
rect 46308 37148 47768 37176
rect 47762 37136 47768 37148
rect 47820 37136 47826 37188
rect 27028 37080 29316 37108
rect 27028 37068 27034 37080
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 17773 36907 17831 36913
rect 17773 36873 17785 36907
rect 17819 36904 17831 36907
rect 18138 36904 18144 36916
rect 17819 36876 18144 36904
rect 17819 36873 17831 36876
rect 17773 36867 17831 36873
rect 18138 36864 18144 36876
rect 18196 36864 18202 36916
rect 19978 36864 19984 36916
rect 20036 36904 20042 36916
rect 21269 36907 21327 36913
rect 21269 36904 21281 36907
rect 20036 36876 21281 36904
rect 20036 36864 20042 36876
rect 21269 36873 21281 36876
rect 21315 36873 21327 36907
rect 21269 36867 21327 36873
rect 22465 36907 22523 36913
rect 22465 36873 22477 36907
rect 22511 36904 22523 36907
rect 23842 36904 23848 36916
rect 22511 36876 23848 36904
rect 22511 36873 22523 36876
rect 22465 36867 22523 36873
rect 23842 36864 23848 36876
rect 23900 36904 23906 36916
rect 23900 36876 24348 36904
rect 23900 36864 23906 36876
rect 17788 36808 22094 36836
rect 17788 36780 17816 36808
rect 1762 36768 1768 36780
rect 1723 36740 1768 36768
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 17678 36768 17684 36780
rect 17639 36740 17684 36768
rect 17678 36728 17684 36740
rect 17736 36728 17742 36780
rect 17770 36728 17776 36780
rect 17828 36728 17834 36780
rect 18690 36728 18696 36780
rect 18748 36768 18754 36780
rect 20717 36771 20775 36777
rect 20717 36768 20729 36771
rect 18748 36740 20729 36768
rect 18748 36728 18754 36740
rect 20717 36737 20729 36740
rect 20763 36737 20775 36771
rect 20717 36731 20775 36737
rect 21085 36771 21143 36777
rect 21085 36737 21097 36771
rect 21131 36768 21143 36771
rect 21726 36768 21732 36780
rect 21131 36740 21732 36768
rect 21131 36737 21143 36740
rect 21085 36731 21143 36737
rect 21726 36728 21732 36740
rect 21784 36728 21790 36780
rect 22066 36768 22094 36808
rect 24320 36777 24348 36876
rect 30837 36839 30895 36845
rect 30837 36836 30849 36839
rect 30038 36808 30849 36836
rect 30837 36805 30849 36808
rect 30883 36805 30895 36839
rect 30837 36799 30895 36805
rect 22281 36771 22339 36777
rect 22281 36768 22293 36771
rect 22066 36740 22293 36768
rect 22281 36737 22293 36740
rect 22327 36768 22339 36771
rect 23109 36771 23167 36777
rect 23109 36768 23121 36771
rect 22327 36740 23121 36768
rect 22327 36737 22339 36740
rect 22281 36731 22339 36737
rect 23109 36737 23121 36740
rect 23155 36737 23167 36771
rect 23109 36731 23167 36737
rect 24305 36771 24363 36777
rect 24305 36737 24317 36771
rect 24351 36768 24363 36771
rect 24670 36768 24676 36780
rect 24351 36740 24676 36768
rect 24351 36737 24363 36740
rect 24305 36731 24363 36737
rect 24670 36728 24676 36740
rect 24728 36728 24734 36780
rect 28166 36728 28172 36780
rect 28224 36768 28230 36780
rect 28534 36768 28540 36780
rect 28224 36740 28540 36768
rect 28224 36728 28230 36740
rect 28534 36728 28540 36740
rect 28592 36728 28598 36780
rect 30742 36768 30748 36780
rect 30703 36740 30748 36768
rect 30742 36728 30748 36740
rect 30800 36728 30806 36780
rect 1949 36703 2007 36709
rect 1949 36669 1961 36703
rect 1995 36700 2007 36703
rect 2222 36700 2228 36712
rect 1995 36672 2228 36700
rect 1995 36669 2007 36672
rect 1949 36663 2007 36669
rect 2222 36660 2228 36672
rect 2280 36660 2286 36712
rect 2774 36700 2780 36712
rect 2735 36672 2780 36700
rect 2774 36660 2780 36672
rect 2832 36660 2838 36712
rect 28813 36703 28871 36709
rect 28813 36669 28825 36703
rect 28859 36700 28871 36703
rect 29454 36700 29460 36712
rect 28859 36672 29460 36700
rect 28859 36669 28871 36672
rect 28813 36663 28871 36669
rect 29454 36660 29460 36672
rect 29512 36660 29518 36712
rect 23382 36632 23388 36644
rect 21100 36604 23388 36632
rect 21100 36573 21128 36604
rect 23382 36592 23388 36604
rect 23440 36592 23446 36644
rect 26970 36632 26976 36644
rect 23492 36604 26976 36632
rect 23492 36576 23520 36604
rect 26970 36592 26976 36604
rect 27028 36592 27034 36644
rect 21085 36567 21143 36573
rect 21085 36533 21097 36567
rect 21131 36533 21143 36567
rect 21085 36527 21143 36533
rect 23201 36567 23259 36573
rect 23201 36533 23213 36567
rect 23247 36564 23259 36567
rect 23474 36564 23480 36576
rect 23247 36536 23480 36564
rect 23247 36533 23259 36536
rect 23201 36527 23259 36533
rect 23474 36524 23480 36536
rect 23532 36524 23538 36576
rect 24394 36564 24400 36576
rect 24355 36536 24400 36564
rect 24394 36524 24400 36536
rect 24452 36524 24458 36576
rect 30282 36564 30288 36576
rect 30243 36536 30288 36564
rect 30282 36524 30288 36536
rect 30340 36524 30346 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 2222 36360 2228 36372
rect 2183 36332 2228 36360
rect 2222 36320 2228 36332
rect 2280 36320 2286 36372
rect 23676 36332 28212 36360
rect 20346 36252 20352 36304
rect 20404 36292 20410 36304
rect 23676 36292 23704 36332
rect 20404 36264 23704 36292
rect 20404 36252 20410 36264
rect 16577 36227 16635 36233
rect 16577 36193 16589 36227
rect 16623 36224 16635 36227
rect 19242 36224 19248 36236
rect 16623 36196 19248 36224
rect 16623 36193 16635 36196
rect 16577 36187 16635 36193
rect 19242 36184 19248 36196
rect 19300 36184 19306 36236
rect 22922 36184 22928 36236
rect 22980 36224 22986 36236
rect 23477 36227 23535 36233
rect 23477 36224 23489 36227
rect 22980 36196 23489 36224
rect 22980 36184 22986 36196
rect 23477 36193 23489 36196
rect 23523 36193 23535 36227
rect 23477 36187 23535 36193
rect 23566 36184 23572 36236
rect 23624 36184 23630 36236
rect 2130 36156 2136 36168
rect 2091 36128 2136 36156
rect 2130 36116 2136 36128
rect 2188 36116 2194 36168
rect 15654 36116 15660 36168
rect 15712 36156 15718 36168
rect 16298 36156 16304 36168
rect 15712 36128 16304 36156
rect 15712 36116 15718 36128
rect 16298 36116 16304 36128
rect 16356 36116 16362 36168
rect 22373 36159 22431 36165
rect 22373 36125 22385 36159
rect 22419 36156 22431 36159
rect 22462 36156 22468 36168
rect 22419 36128 22468 36156
rect 22419 36125 22431 36128
rect 22373 36119 22431 36125
rect 22462 36116 22468 36128
rect 22520 36156 22526 36168
rect 22738 36156 22744 36168
rect 22520 36128 22744 36156
rect 22520 36116 22526 36128
rect 22738 36116 22744 36128
rect 22796 36116 22802 36168
rect 23109 36159 23167 36165
rect 23109 36125 23121 36159
rect 23155 36125 23167 36159
rect 23290 36156 23296 36168
rect 23251 36128 23296 36156
rect 23109 36119 23167 36125
rect 17310 36048 17316 36100
rect 17368 36048 17374 36100
rect 23124 36088 23152 36119
rect 23290 36116 23296 36128
rect 23348 36116 23354 36168
rect 23385 36159 23443 36165
rect 23385 36125 23397 36159
rect 23431 36156 23443 36159
rect 23584 36156 23612 36184
rect 23676 36165 23704 36264
rect 25406 36224 25412 36236
rect 25367 36196 25412 36224
rect 25406 36184 25412 36196
rect 25464 36184 25470 36236
rect 25685 36227 25743 36233
rect 25685 36193 25697 36227
rect 25731 36224 25743 36227
rect 26418 36224 26424 36236
rect 25731 36196 26424 36224
rect 25731 36193 25743 36196
rect 25685 36187 25743 36193
rect 26418 36184 26424 36196
rect 26476 36184 26482 36236
rect 23431 36128 23612 36156
rect 23661 36159 23719 36165
rect 23431 36125 23443 36128
rect 23385 36119 23443 36125
rect 23661 36125 23673 36159
rect 23707 36125 23719 36159
rect 23661 36119 23719 36125
rect 23566 36088 23572 36100
rect 23124 36060 23572 36088
rect 23566 36048 23572 36060
rect 23624 36048 23630 36100
rect 27062 36088 27068 36100
rect 26910 36060 27068 36088
rect 27062 36048 27068 36060
rect 27120 36048 27126 36100
rect 27890 36048 27896 36100
rect 27948 36088 27954 36100
rect 28184 36097 28212 36332
rect 29730 36156 29736 36168
rect 29691 36128 29736 36156
rect 29730 36116 29736 36128
rect 29788 36116 29794 36168
rect 29914 36156 29920 36168
rect 29875 36128 29920 36156
rect 29914 36116 29920 36128
rect 29972 36116 29978 36168
rect 30006 36116 30012 36168
rect 30064 36156 30070 36168
rect 30064 36128 30109 36156
rect 30064 36116 30070 36128
rect 27985 36091 28043 36097
rect 27985 36088 27997 36091
rect 27948 36060 27997 36088
rect 27948 36048 27954 36060
rect 27985 36057 27997 36060
rect 28031 36057 28043 36091
rect 27985 36051 28043 36057
rect 28169 36091 28227 36097
rect 28169 36057 28181 36091
rect 28215 36088 28227 36091
rect 28718 36088 28724 36100
rect 28215 36060 28724 36088
rect 28215 36057 28227 36060
rect 28169 36051 28227 36057
rect 28718 36048 28724 36060
rect 28776 36088 28782 36100
rect 29638 36088 29644 36100
rect 28776 36060 29644 36088
rect 28776 36048 28782 36060
rect 29638 36048 29644 36060
rect 29696 36048 29702 36100
rect 18046 36020 18052 36032
rect 18007 35992 18052 36020
rect 18046 35980 18052 35992
rect 18104 36020 18110 36032
rect 19058 36020 19064 36032
rect 18104 35992 19064 36020
rect 18104 35980 18110 35992
rect 19058 35980 19064 35992
rect 19116 35980 19122 36032
rect 22557 36023 22615 36029
rect 22557 35989 22569 36023
rect 22603 36020 22615 36023
rect 22922 36020 22928 36032
rect 22603 35992 22928 36020
rect 22603 35989 22615 35992
rect 22557 35983 22615 35989
rect 22922 35980 22928 35992
rect 22980 36020 22986 36032
rect 23290 36020 23296 36032
rect 22980 35992 23296 36020
rect 22980 35980 22986 35992
rect 23290 35980 23296 35992
rect 23348 35980 23354 36032
rect 23658 35980 23664 36032
rect 23716 36020 23722 36032
rect 23845 36023 23903 36029
rect 23845 36020 23857 36023
rect 23716 35992 23857 36020
rect 23716 35980 23722 35992
rect 23845 35989 23857 35992
rect 23891 35989 23903 36023
rect 27154 36020 27160 36032
rect 27115 35992 27160 36020
rect 23845 35983 23903 35989
rect 27154 35980 27160 35992
rect 27212 35980 27218 36032
rect 28074 35980 28080 36032
rect 28132 36020 28138 36032
rect 28994 36020 29000 36032
rect 28132 35992 29000 36020
rect 28132 35980 28138 35992
rect 28994 35980 29000 35992
rect 29052 35980 29058 36032
rect 29549 36023 29607 36029
rect 29549 35989 29561 36023
rect 29595 36020 29607 36023
rect 29822 36020 29828 36032
rect 29595 35992 29828 36020
rect 29595 35989 29607 35992
rect 29549 35983 29607 35989
rect 29822 35980 29828 35992
rect 29880 35980 29886 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 17310 35816 17316 35828
rect 17271 35788 17316 35816
rect 17310 35776 17316 35788
rect 17368 35776 17374 35828
rect 18892 35788 19196 35816
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 16666 35640 16672 35692
rect 16724 35680 16730 35692
rect 17221 35683 17279 35689
rect 17221 35680 17233 35683
rect 16724 35652 17233 35680
rect 16724 35640 16730 35652
rect 17221 35649 17233 35652
rect 17267 35680 17279 35683
rect 17678 35680 17684 35692
rect 17267 35652 17684 35680
rect 17267 35649 17279 35652
rect 17221 35643 17279 35649
rect 17678 35640 17684 35652
rect 17736 35640 17742 35692
rect 17862 35680 17868 35692
rect 17823 35652 17868 35680
rect 17862 35640 17868 35652
rect 17920 35640 17926 35692
rect 18046 35680 18052 35692
rect 18007 35652 18052 35680
rect 18046 35640 18052 35652
rect 18104 35640 18110 35692
rect 18892 35689 18920 35788
rect 19058 35748 19064 35760
rect 18984 35720 19064 35748
rect 18984 35689 19012 35720
rect 19058 35708 19064 35720
rect 19116 35708 19122 35760
rect 19168 35748 19196 35788
rect 19242 35776 19248 35828
rect 19300 35816 19306 35828
rect 19429 35819 19487 35825
rect 19429 35816 19441 35819
rect 19300 35788 19441 35816
rect 19300 35776 19306 35788
rect 19429 35785 19441 35788
rect 19475 35785 19487 35819
rect 19429 35779 19487 35785
rect 23750 35776 23756 35828
rect 23808 35816 23814 35828
rect 24670 35816 24676 35828
rect 23808 35788 24676 35816
rect 23808 35776 23814 35788
rect 24670 35776 24676 35788
rect 24728 35816 24734 35828
rect 25133 35819 25191 35825
rect 25133 35816 25145 35819
rect 24728 35788 25145 35816
rect 24728 35776 24734 35788
rect 25133 35785 25145 35788
rect 25179 35785 25191 35819
rect 27062 35816 27068 35828
rect 27023 35788 27068 35816
rect 25133 35779 25191 35785
rect 27062 35776 27068 35788
rect 27120 35776 27126 35828
rect 27709 35819 27767 35825
rect 27709 35785 27721 35819
rect 27755 35816 27767 35819
rect 29454 35816 29460 35828
rect 27755 35788 28580 35816
rect 29415 35788 29460 35816
rect 27755 35785 27767 35788
rect 27709 35779 27767 35785
rect 19334 35748 19340 35760
rect 19168 35720 19340 35748
rect 19334 35708 19340 35720
rect 19392 35708 19398 35760
rect 23658 35748 23664 35760
rect 23619 35720 23664 35748
rect 23658 35708 23664 35720
rect 23716 35708 23722 35760
rect 24394 35708 24400 35760
rect 24452 35708 24458 35760
rect 28258 35711 28264 35760
rect 28251 35708 28264 35711
rect 28316 35708 28322 35760
rect 28251 35705 28309 35708
rect 18693 35683 18751 35689
rect 18693 35649 18705 35683
rect 18739 35649 18751 35683
rect 18693 35643 18751 35649
rect 18877 35683 18935 35689
rect 18877 35649 18889 35683
rect 18923 35649 18935 35683
rect 18877 35643 18935 35649
rect 18969 35683 19027 35689
rect 18969 35649 18981 35683
rect 19015 35649 19027 35683
rect 18969 35643 19027 35649
rect 19245 35683 19303 35689
rect 19245 35649 19257 35683
rect 19291 35680 19303 35683
rect 20346 35680 20352 35692
rect 19291 35652 20352 35680
rect 19291 35649 19303 35652
rect 19245 35643 19303 35649
rect 18708 35544 18736 35643
rect 20346 35640 20352 35652
rect 20404 35640 20410 35692
rect 22462 35680 22468 35692
rect 22423 35652 22468 35680
rect 22462 35640 22468 35652
rect 22520 35640 22526 35692
rect 22554 35640 22560 35692
rect 22612 35680 22618 35692
rect 22830 35680 22836 35692
rect 22612 35652 22657 35680
rect 22791 35652 22836 35680
rect 22612 35640 22618 35652
rect 22830 35640 22836 35652
rect 22888 35640 22894 35692
rect 26970 35680 26976 35692
rect 26931 35652 26976 35680
rect 26970 35640 26976 35652
rect 27028 35640 27034 35692
rect 27798 35640 27804 35692
rect 27856 35680 27862 35692
rect 27893 35683 27951 35689
rect 27893 35680 27905 35683
rect 27856 35652 27905 35680
rect 27856 35640 27862 35652
rect 27893 35649 27905 35652
rect 27939 35649 27951 35683
rect 27893 35643 27951 35649
rect 27982 35640 27988 35692
rect 28040 35680 28046 35692
rect 28128 35683 28186 35689
rect 28040 35652 28085 35680
rect 28040 35640 28046 35652
rect 28128 35649 28140 35683
rect 28174 35649 28186 35683
rect 28251 35671 28263 35705
rect 28297 35671 28309 35705
rect 28251 35665 28309 35671
rect 28552 35680 28580 35788
rect 29454 35776 29460 35788
rect 29512 35776 29518 35828
rect 29546 35776 29552 35828
rect 29604 35816 29610 35828
rect 43990 35816 43996 35828
rect 29604 35788 43996 35816
rect 29604 35776 29610 35788
rect 43990 35776 43996 35788
rect 44048 35776 44054 35828
rect 29086 35748 29092 35760
rect 28920 35720 29092 35748
rect 28920 35691 28948 35720
rect 29086 35708 29092 35720
rect 29144 35708 29150 35760
rect 29638 35748 29644 35760
rect 29288 35720 29644 35748
rect 28721 35683 28779 35689
rect 28721 35680 28733 35683
rect 28552 35652 28733 35680
rect 28128 35643 28186 35649
rect 28721 35649 28733 35652
rect 28767 35649 28779 35683
rect 28721 35643 28779 35649
rect 28905 35685 28963 35691
rect 28905 35651 28917 35685
rect 28951 35651 28963 35685
rect 28905 35645 28963 35651
rect 19058 35612 19064 35624
rect 19019 35584 19064 35612
rect 19058 35572 19064 35584
rect 19116 35572 19122 35624
rect 20714 35572 20720 35624
rect 20772 35612 20778 35624
rect 22370 35612 22376 35624
rect 20772 35584 22376 35612
rect 20772 35572 20778 35584
rect 22370 35572 22376 35584
rect 22428 35612 22434 35624
rect 23385 35615 23443 35621
rect 23385 35612 23397 35615
rect 22428 35584 23397 35612
rect 22428 35572 22434 35584
rect 23385 35581 23397 35584
rect 23431 35581 23443 35615
rect 23385 35575 23443 35581
rect 27614 35572 27620 35624
rect 27672 35612 27678 35624
rect 28143 35612 28171 35643
rect 28994 35640 29000 35692
rect 29052 35680 29058 35692
rect 29288 35689 29316 35720
rect 29638 35708 29644 35720
rect 29696 35708 29702 35760
rect 29273 35683 29331 35689
rect 29052 35652 29097 35680
rect 29052 35640 29058 35652
rect 29273 35649 29285 35683
rect 29319 35649 29331 35683
rect 29914 35680 29920 35692
rect 29827 35652 29920 35680
rect 29273 35643 29331 35649
rect 29914 35640 29920 35652
rect 29972 35680 29978 35692
rect 30926 35680 30932 35692
rect 29972 35652 30420 35680
rect 30887 35652 30932 35680
rect 29972 35640 29978 35652
rect 27672 35584 28171 35612
rect 29089 35615 29147 35621
rect 27672 35572 27678 35584
rect 29089 35581 29101 35615
rect 29135 35612 29147 35615
rect 29454 35612 29460 35624
rect 29135 35584 29460 35612
rect 29135 35581 29147 35584
rect 29089 35575 29147 35581
rect 29454 35572 29460 35584
rect 29512 35572 29518 35624
rect 29730 35572 29736 35624
rect 29788 35612 29794 35624
rect 30009 35615 30067 35621
rect 30009 35612 30021 35615
rect 29788 35584 30021 35612
rect 29788 35572 29794 35584
rect 30009 35581 30021 35584
rect 30055 35581 30067 35615
rect 30392 35612 30420 35652
rect 30926 35640 30932 35652
rect 30984 35640 30990 35692
rect 31846 35640 31852 35692
rect 31904 35680 31910 35692
rect 32125 35683 32183 35689
rect 32125 35680 32137 35683
rect 31904 35652 32137 35680
rect 31904 35640 31910 35652
rect 32125 35649 32137 35652
rect 32171 35649 32183 35683
rect 32125 35643 32183 35649
rect 31021 35615 31079 35621
rect 31021 35612 31033 35615
rect 30392 35584 31033 35612
rect 30009 35575 30067 35581
rect 31021 35581 31033 35584
rect 31067 35612 31079 35615
rect 31754 35612 31760 35624
rect 31067 35584 31760 35612
rect 31067 35581 31079 35584
rect 31021 35575 31079 35581
rect 31754 35572 31760 35584
rect 31812 35572 31818 35624
rect 19794 35544 19800 35556
rect 18708 35516 19800 35544
rect 19794 35504 19800 35516
rect 19852 35504 19858 35556
rect 27798 35504 27804 35556
rect 27856 35544 27862 35556
rect 30285 35547 30343 35553
rect 30285 35544 30297 35547
rect 27856 35516 30297 35544
rect 27856 35504 27862 35516
rect 30285 35513 30297 35516
rect 30331 35513 30343 35547
rect 31294 35544 31300 35556
rect 31255 35516 31300 35544
rect 30285 35507 30343 35513
rect 31294 35504 31300 35516
rect 31352 35504 31358 35556
rect 1397 35479 1455 35485
rect 1397 35445 1409 35479
rect 1443 35476 1455 35479
rect 1486 35476 1492 35488
rect 1443 35448 1492 35476
rect 1443 35445 1455 35448
rect 1397 35439 1455 35445
rect 1486 35436 1492 35448
rect 1544 35436 1550 35488
rect 18233 35479 18291 35485
rect 18233 35445 18245 35479
rect 18279 35476 18291 35479
rect 18322 35476 18328 35488
rect 18279 35448 18328 35476
rect 18279 35445 18291 35448
rect 18233 35439 18291 35445
rect 18322 35436 18328 35448
rect 18380 35436 18386 35488
rect 22278 35476 22284 35488
rect 22239 35448 22284 35476
rect 22278 35436 22284 35448
rect 22336 35436 22342 35488
rect 22741 35479 22799 35485
rect 22741 35445 22753 35479
rect 22787 35476 22799 35479
rect 29086 35476 29092 35488
rect 22787 35448 29092 35476
rect 22787 35445 22799 35448
rect 22741 35439 22799 35445
rect 29086 35436 29092 35448
rect 29144 35436 29150 35488
rect 29730 35436 29736 35488
rect 29788 35476 29794 35488
rect 30006 35476 30012 35488
rect 29788 35448 30012 35476
rect 29788 35436 29794 35448
rect 30006 35436 30012 35448
rect 30064 35476 30070 35488
rect 30101 35479 30159 35485
rect 30101 35476 30113 35479
rect 30064 35448 30113 35476
rect 30064 35436 30070 35448
rect 30101 35445 30113 35448
rect 30147 35476 30159 35479
rect 30926 35476 30932 35488
rect 30147 35448 30932 35476
rect 30147 35445 30159 35448
rect 30101 35439 30159 35445
rect 30926 35436 30932 35448
rect 30984 35436 30990 35488
rect 32122 35436 32128 35488
rect 32180 35476 32186 35488
rect 32217 35479 32275 35485
rect 32217 35476 32229 35479
rect 32180 35448 32229 35476
rect 32180 35436 32186 35448
rect 32217 35445 32229 35448
rect 32263 35445 32275 35479
rect 32217 35439 32275 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 18230 35272 18236 35284
rect 18191 35244 18236 35272
rect 18230 35232 18236 35244
rect 18288 35232 18294 35284
rect 19613 35275 19671 35281
rect 19613 35241 19625 35275
rect 19659 35241 19671 35275
rect 19794 35272 19800 35284
rect 19755 35244 19800 35272
rect 19613 35235 19671 35241
rect 17313 35207 17371 35213
rect 17313 35173 17325 35207
rect 17359 35204 17371 35207
rect 19628 35204 19656 35235
rect 19794 35232 19800 35244
rect 19852 35232 19858 35284
rect 22186 35272 22192 35284
rect 19904 35244 22192 35272
rect 19904 35204 19932 35244
rect 22186 35232 22192 35244
rect 22244 35232 22250 35284
rect 22465 35275 22523 35281
rect 22465 35241 22477 35275
rect 22511 35272 22523 35275
rect 22554 35272 22560 35284
rect 22511 35244 22560 35272
rect 22511 35241 22523 35244
rect 22465 35235 22523 35241
rect 22554 35232 22560 35244
rect 22612 35232 22618 35284
rect 23477 35275 23535 35281
rect 23477 35241 23489 35275
rect 23523 35272 23535 35275
rect 24946 35272 24952 35284
rect 23523 35244 24952 35272
rect 23523 35241 23535 35244
rect 23477 35235 23535 35241
rect 24946 35232 24952 35244
rect 25004 35232 25010 35284
rect 25409 35275 25467 35281
rect 25409 35241 25421 35275
rect 25455 35241 25467 35275
rect 25409 35235 25467 35241
rect 17359 35176 19564 35204
rect 19628 35176 19932 35204
rect 17359 35173 17371 35176
rect 17313 35167 17371 35173
rect 18046 35136 18052 35148
rect 17512 35108 18052 35136
rect 17512 35077 17540 35108
rect 18046 35096 18052 35108
rect 18104 35136 18110 35148
rect 18325 35139 18383 35145
rect 18325 35136 18337 35139
rect 18104 35108 18337 35136
rect 18104 35096 18110 35108
rect 18325 35105 18337 35108
rect 18371 35105 18383 35139
rect 18325 35099 18383 35105
rect 18414 35096 18420 35148
rect 18472 35136 18478 35148
rect 19058 35136 19064 35148
rect 18472 35108 19064 35136
rect 18472 35096 18478 35108
rect 19058 35096 19064 35108
rect 19116 35096 19122 35148
rect 19536 35145 19564 35176
rect 23566 35164 23572 35216
rect 23624 35204 23630 35216
rect 23661 35207 23719 35213
rect 23661 35204 23673 35207
rect 23624 35176 23673 35204
rect 23624 35164 23630 35176
rect 23661 35173 23673 35176
rect 23707 35173 23719 35207
rect 25424 35204 25452 35235
rect 26418 35232 26424 35284
rect 26476 35272 26482 35284
rect 26789 35275 26847 35281
rect 26789 35272 26801 35275
rect 26476 35244 26801 35272
rect 26476 35232 26482 35244
rect 26789 35241 26801 35244
rect 26835 35241 26847 35275
rect 26789 35235 26847 35241
rect 27154 35232 27160 35284
rect 27212 35272 27218 35284
rect 27249 35275 27307 35281
rect 27249 35272 27261 35275
rect 27212 35244 27261 35272
rect 27212 35232 27218 35244
rect 27249 35241 27261 35244
rect 27295 35241 27307 35275
rect 27249 35235 27307 35241
rect 28258 35232 28264 35284
rect 28316 35272 28322 35284
rect 28537 35275 28595 35281
rect 28537 35272 28549 35275
rect 28316 35244 28549 35272
rect 28316 35232 28322 35244
rect 28537 35241 28549 35244
rect 28583 35241 28595 35275
rect 28537 35235 28595 35241
rect 28997 35275 29055 35281
rect 28997 35241 29009 35275
rect 29043 35272 29055 35275
rect 29178 35272 29184 35284
rect 29043 35244 29184 35272
rect 29043 35241 29055 35244
rect 28997 35235 29055 35241
rect 29178 35232 29184 35244
rect 29236 35232 29242 35284
rect 29638 35272 29644 35284
rect 29599 35244 29644 35272
rect 29638 35232 29644 35244
rect 29696 35232 29702 35284
rect 27062 35204 27068 35216
rect 25424 35176 27068 35204
rect 23661 35167 23719 35173
rect 27062 35164 27068 35176
rect 27120 35164 27126 35216
rect 27798 35164 27804 35216
rect 27856 35204 27862 35216
rect 27856 35176 28488 35204
rect 27856 35164 27862 35176
rect 19521 35139 19579 35145
rect 19521 35105 19533 35139
rect 19567 35105 19579 35139
rect 20714 35136 20720 35148
rect 20675 35108 20720 35136
rect 19521 35099 19579 35105
rect 20714 35096 20720 35108
rect 20772 35096 20778 35148
rect 21082 35096 21088 35148
rect 21140 35136 21146 35148
rect 25225 35139 25283 35145
rect 25225 35136 25237 35139
rect 21140 35108 25237 35136
rect 21140 35096 21146 35108
rect 25225 35105 25237 35108
rect 25271 35136 25283 35139
rect 25958 35136 25964 35148
rect 25271 35108 25964 35136
rect 25271 35105 25283 35108
rect 25225 35099 25283 35105
rect 25958 35096 25964 35108
rect 26016 35096 26022 35148
rect 26513 35139 26571 35145
rect 26513 35105 26525 35139
rect 26559 35136 26571 35139
rect 27154 35136 27160 35148
rect 26559 35108 27160 35136
rect 26559 35105 26571 35108
rect 26513 35099 26571 35105
rect 27154 35096 27160 35108
rect 27212 35096 27218 35148
rect 27338 35096 27344 35148
rect 27396 35136 27402 35148
rect 27396 35108 28304 35136
rect 27396 35096 27402 35108
rect 17497 35071 17555 35077
rect 17497 35037 17509 35071
rect 17543 35037 17555 35071
rect 17497 35031 17555 35037
rect 17681 35071 17739 35077
rect 17681 35037 17693 35071
rect 17727 35037 17739 35071
rect 17681 35031 17739 35037
rect 17773 35071 17831 35077
rect 17773 35037 17785 35071
rect 17819 35068 17831 35071
rect 17862 35068 17868 35080
rect 17819 35040 17868 35068
rect 17819 35037 17831 35040
rect 17773 35031 17831 35037
rect 17696 35000 17724 35031
rect 17862 35028 17868 35040
rect 17920 35068 17926 35080
rect 18506 35068 18512 35080
rect 17920 35040 18276 35068
rect 18467 35040 18512 35068
rect 17920 35028 17926 35040
rect 18046 35000 18052 35012
rect 17696 34972 18052 35000
rect 18046 34960 18052 34972
rect 18104 34960 18110 35012
rect 18248 35009 18276 35040
rect 18506 35028 18512 35040
rect 18564 35028 18570 35080
rect 18598 35028 18604 35080
rect 18656 35068 18662 35080
rect 19245 35071 19303 35077
rect 19245 35068 19257 35071
rect 18656 35040 19257 35068
rect 18656 35028 18662 35040
rect 19245 35037 19257 35040
rect 19291 35037 19303 35071
rect 23106 35068 23112 35080
rect 23067 35040 23112 35068
rect 19245 35031 19303 35037
rect 23106 35028 23112 35040
rect 23164 35028 23170 35080
rect 23382 35068 23388 35080
rect 23343 35040 23388 35068
rect 23382 35028 23388 35040
rect 23440 35028 23446 35080
rect 24670 35028 24676 35080
rect 24728 35068 24734 35080
rect 25409 35071 25467 35077
rect 25409 35068 25421 35071
rect 24728 35040 25421 35068
rect 24728 35028 24734 35040
rect 25409 35037 25421 35040
rect 25455 35037 25467 35071
rect 25409 35031 25467 35037
rect 26605 35071 26663 35077
rect 26605 35037 26617 35071
rect 26651 35068 26663 35071
rect 27430 35068 27436 35080
rect 26651 35040 27436 35068
rect 26651 35037 26663 35040
rect 26605 35031 26663 35037
rect 27430 35028 27436 35040
rect 27488 35028 27494 35080
rect 27522 35028 27528 35080
rect 27580 35068 27586 35080
rect 27580 35040 27625 35068
rect 27580 35028 27586 35040
rect 18233 35003 18291 35009
rect 18233 34969 18245 35003
rect 18279 35000 18291 35003
rect 20346 35000 20352 35012
rect 18279 34972 20352 35000
rect 18279 34969 18291 34972
rect 18233 34963 18291 34969
rect 20346 34960 20352 34972
rect 20404 34960 20410 35012
rect 20990 35000 20996 35012
rect 20951 34972 20996 35000
rect 20990 34960 20996 34972
rect 21048 34960 21054 35012
rect 21450 34960 21456 35012
rect 21508 34960 21514 35012
rect 23198 35000 23204 35012
rect 22388 34972 23204 35000
rect 18693 34935 18751 34941
rect 18693 34901 18705 34935
rect 18739 34932 18751 34935
rect 19058 34932 19064 34944
rect 18739 34904 19064 34932
rect 18739 34901 18751 34904
rect 18693 34895 18751 34901
rect 19058 34892 19064 34904
rect 19116 34892 19122 34944
rect 19978 34892 19984 34944
rect 20036 34932 20042 34944
rect 22388 34932 22416 34972
rect 23198 34960 23204 34972
rect 23256 34960 23262 35012
rect 25133 35003 25191 35009
rect 25133 34969 25145 35003
rect 25179 35000 25191 35003
rect 25314 35000 25320 35012
rect 25179 34972 25320 35000
rect 25179 34969 25191 34972
rect 25133 34963 25191 34969
rect 25314 34960 25320 34972
rect 25372 35000 25378 35012
rect 27246 35000 27252 35012
rect 25372 34972 26280 35000
rect 27207 34972 27252 35000
rect 25372 34960 25378 34972
rect 20036 34904 22416 34932
rect 20036 34892 20042 34904
rect 22462 34892 22468 34944
rect 22520 34932 22526 34944
rect 25593 34935 25651 34941
rect 25593 34932 25605 34935
rect 22520 34904 25605 34932
rect 22520 34892 22526 34904
rect 25593 34901 25605 34904
rect 25639 34901 25651 34935
rect 25593 34895 25651 34901
rect 25774 34892 25780 34944
rect 25832 34932 25838 34944
rect 26145 34935 26203 34941
rect 26145 34932 26157 34935
rect 25832 34904 26157 34932
rect 25832 34892 25838 34904
rect 26145 34901 26157 34904
rect 26191 34901 26203 34935
rect 26252 34932 26280 34972
rect 27246 34960 27252 34972
rect 27304 34960 27310 35012
rect 28276 35000 28304 35108
rect 28460 35077 28488 35176
rect 28552 35176 31156 35204
rect 28552 35148 28580 35176
rect 28534 35096 28540 35148
rect 28592 35096 28598 35148
rect 29730 35136 29736 35148
rect 29691 35108 29736 35136
rect 29730 35096 29736 35108
rect 29788 35096 29794 35148
rect 31128 35145 31156 35176
rect 31113 35139 31171 35145
rect 31113 35105 31125 35139
rect 31159 35105 31171 35139
rect 31113 35099 31171 35105
rect 28445 35071 28503 35077
rect 28445 35037 28457 35071
rect 28491 35037 28503 35071
rect 28445 35031 28503 35037
rect 28813 35071 28871 35077
rect 28813 35037 28825 35071
rect 28859 35068 28871 35071
rect 29638 35068 29644 35080
rect 28859 35040 29644 35068
rect 28859 35037 28871 35040
rect 28813 35031 28871 35037
rect 29638 35028 29644 35040
rect 29696 35028 29702 35080
rect 29825 35071 29883 35077
rect 29825 35037 29837 35071
rect 29871 35068 29883 35071
rect 30282 35068 30288 35080
rect 29871 35040 30288 35068
rect 29871 35037 29883 35040
rect 29825 35031 29883 35037
rect 30282 35028 30288 35040
rect 30340 35028 30346 35080
rect 48130 35068 48136 35080
rect 48091 35040 48136 35068
rect 48130 35028 48136 35040
rect 48188 35028 48194 35080
rect 29549 35003 29607 35009
rect 28276 34972 28672 35000
rect 28644 34944 28672 34972
rect 29549 34969 29561 35003
rect 29595 35000 29607 35003
rect 30098 35000 30104 35012
rect 29595 34972 30104 35000
rect 29595 34969 29607 34972
rect 29549 34963 29607 34969
rect 30098 34960 30104 34972
rect 30156 34960 30162 35012
rect 31018 34960 31024 35012
rect 31076 35000 31082 35012
rect 31389 35003 31447 35009
rect 31389 35000 31401 35003
rect 31076 34972 31401 35000
rect 31076 34960 31082 34972
rect 31389 34969 31401 34972
rect 31435 34969 31447 35003
rect 31389 34963 31447 34969
rect 32122 34960 32128 35012
rect 32180 34960 32186 35012
rect 27709 34935 27767 34941
rect 27709 34932 27721 34935
rect 26252 34904 27721 34932
rect 26145 34895 26203 34901
rect 27709 34901 27721 34904
rect 27755 34901 27767 34935
rect 27709 34895 27767 34901
rect 28626 34892 28632 34944
rect 28684 34932 28690 34944
rect 30009 34935 30067 34941
rect 30009 34932 30021 34935
rect 28684 34904 30021 34932
rect 28684 34892 28690 34904
rect 30009 34901 30021 34904
rect 30055 34901 30067 34935
rect 32858 34932 32864 34944
rect 32819 34904 32864 34932
rect 30009 34895 30067 34901
rect 32858 34892 32864 34904
rect 32916 34892 32922 34944
rect 47118 34892 47124 34944
rect 47176 34932 47182 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47176 34904 47961 34932
rect 47176 34892 47182 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 18598 34728 18604 34740
rect 18559 34700 18604 34728
rect 18598 34688 18604 34700
rect 18656 34688 18662 34740
rect 19521 34731 19579 34737
rect 19521 34697 19533 34731
rect 19567 34728 19579 34731
rect 21082 34728 21088 34740
rect 19567 34700 21088 34728
rect 19567 34697 19579 34700
rect 19521 34691 19579 34697
rect 21082 34688 21088 34700
rect 21140 34688 21146 34740
rect 21177 34731 21235 34737
rect 21177 34697 21189 34731
rect 21223 34728 21235 34731
rect 21450 34728 21456 34740
rect 21223 34700 21456 34728
rect 21223 34697 21235 34700
rect 21177 34691 21235 34697
rect 21450 34688 21456 34700
rect 21508 34688 21514 34740
rect 24946 34728 24952 34740
rect 24907 34700 24952 34728
rect 24946 34688 24952 34700
rect 25004 34688 25010 34740
rect 27430 34688 27436 34740
rect 27488 34728 27494 34740
rect 28169 34731 28227 34737
rect 28169 34728 28181 34731
rect 27488 34700 28181 34728
rect 27488 34688 27494 34700
rect 28169 34697 28181 34700
rect 28215 34697 28227 34731
rect 28169 34691 28227 34697
rect 28721 34731 28779 34737
rect 28721 34697 28733 34731
rect 28767 34697 28779 34731
rect 28721 34691 28779 34697
rect 30193 34731 30251 34737
rect 30193 34697 30205 34731
rect 30239 34728 30251 34731
rect 31754 34728 31760 34740
rect 30239 34700 31760 34728
rect 30239 34697 30251 34700
rect 30193 34691 30251 34697
rect 17313 34663 17371 34669
rect 17313 34629 17325 34663
rect 17359 34660 17371 34663
rect 17494 34660 17500 34672
rect 17359 34632 17500 34660
rect 17359 34629 17371 34632
rect 17313 34623 17371 34629
rect 17494 34620 17500 34632
rect 17552 34620 17558 34672
rect 18141 34663 18199 34669
rect 18141 34629 18153 34663
rect 18187 34660 18199 34663
rect 18690 34660 18696 34672
rect 18187 34632 18696 34660
rect 18187 34629 18199 34632
rect 18141 34623 18199 34629
rect 18690 34620 18696 34632
rect 18748 34620 18754 34672
rect 19058 34660 19064 34672
rect 19019 34632 19064 34660
rect 19058 34620 19064 34632
rect 19116 34620 19122 34672
rect 19978 34660 19984 34672
rect 19260 34632 19984 34660
rect 17126 34592 17132 34604
rect 17087 34564 17132 34592
rect 17126 34552 17132 34564
rect 17184 34552 17190 34604
rect 17405 34595 17463 34601
rect 17405 34561 17417 34595
rect 17451 34592 17463 34595
rect 17954 34592 17960 34604
rect 17451 34564 17960 34592
rect 17451 34561 17463 34564
rect 17405 34555 17463 34561
rect 17954 34552 17960 34564
rect 18012 34552 18018 34604
rect 18322 34592 18328 34604
rect 18283 34564 18328 34592
rect 18322 34552 18328 34564
rect 18380 34552 18386 34604
rect 18417 34595 18475 34601
rect 18417 34561 18429 34595
rect 18463 34592 18475 34595
rect 18874 34592 18880 34604
rect 18463 34564 18880 34592
rect 18463 34561 18475 34564
rect 18417 34555 18475 34561
rect 18874 34552 18880 34564
rect 18932 34552 18938 34604
rect 19260 34601 19288 34632
rect 19978 34620 19984 34632
rect 20036 34620 20042 34672
rect 22554 34660 22560 34672
rect 20916 34632 22560 34660
rect 19245 34595 19303 34601
rect 19245 34561 19257 34595
rect 19291 34561 19303 34595
rect 19245 34555 19303 34561
rect 19337 34595 19395 34601
rect 19337 34561 19349 34595
rect 19383 34561 19395 34595
rect 19337 34555 19395 34561
rect 20243 34595 20301 34601
rect 20243 34561 20255 34595
rect 20289 34592 20301 34595
rect 20346 34592 20352 34604
rect 20289 34564 20352 34592
rect 20289 34561 20301 34564
rect 20243 34555 20301 34561
rect 18892 34524 18920 34552
rect 19352 34524 19380 34555
rect 20346 34552 20352 34564
rect 20404 34592 20410 34604
rect 20916 34592 20944 34632
rect 22554 34620 22560 34632
rect 22612 34620 22618 34672
rect 25958 34660 25964 34672
rect 25919 34632 25964 34660
rect 25958 34620 25964 34632
rect 26016 34660 26022 34672
rect 26973 34663 27031 34669
rect 26016 34632 26280 34660
rect 26016 34620 26022 34632
rect 21082 34592 21088 34604
rect 20404 34564 20944 34592
rect 21043 34564 21088 34592
rect 20404 34552 20410 34564
rect 21082 34552 21088 34564
rect 21140 34552 21146 34604
rect 22094 34552 22100 34604
rect 22152 34592 22158 34604
rect 22649 34595 22707 34601
rect 22649 34592 22661 34595
rect 22152 34564 22661 34592
rect 22152 34552 22158 34564
rect 22649 34561 22661 34564
rect 22695 34592 22707 34595
rect 23106 34592 23112 34604
rect 22695 34564 23112 34592
rect 22695 34561 22707 34564
rect 22649 34555 22707 34561
rect 23106 34552 23112 34564
rect 23164 34552 23170 34604
rect 24670 34552 24676 34604
rect 24728 34592 24734 34604
rect 25133 34595 25191 34601
rect 25133 34592 25145 34595
rect 24728 34564 25145 34592
rect 24728 34552 24734 34564
rect 25133 34561 25145 34564
rect 25179 34561 25191 34595
rect 25314 34592 25320 34604
rect 25275 34564 25320 34592
rect 25133 34555 25191 34561
rect 25314 34552 25320 34564
rect 25372 34552 25378 34604
rect 26142 34592 26148 34604
rect 26103 34564 26148 34592
rect 26142 34552 26148 34564
rect 26200 34552 26206 34604
rect 26252 34592 26280 34632
rect 26973 34629 26985 34663
rect 27019 34660 27031 34663
rect 27338 34660 27344 34672
rect 27019 34632 27344 34660
rect 27019 34629 27031 34632
rect 26973 34623 27031 34629
rect 27338 34620 27344 34632
rect 27396 34620 27402 34672
rect 27614 34620 27620 34672
rect 27672 34660 27678 34672
rect 28736 34660 28764 34691
rect 31754 34688 31760 34700
rect 31812 34728 31818 34740
rect 32122 34728 32128 34740
rect 31812 34700 32128 34728
rect 31812 34688 31818 34700
rect 32122 34688 32128 34700
rect 32180 34688 32186 34740
rect 27672 34632 28764 34660
rect 27672 34620 27678 34632
rect 26252 34564 27108 34592
rect 20073 34527 20131 34533
rect 20073 34524 20085 34527
rect 18892 34496 19380 34524
rect 19444 34496 20085 34524
rect 18046 34416 18052 34468
rect 18104 34456 18110 34468
rect 19242 34456 19248 34468
rect 18104 34428 19248 34456
rect 18104 34416 18110 34428
rect 19242 34416 19248 34428
rect 19300 34456 19306 34468
rect 19444 34456 19472 34496
rect 20073 34493 20085 34496
rect 20119 34493 20131 34527
rect 20073 34487 20131 34493
rect 22373 34527 22431 34533
rect 22373 34493 22385 34527
rect 22419 34524 22431 34527
rect 22462 34524 22468 34536
rect 22419 34496 22468 34524
rect 22419 34493 22431 34496
rect 22373 34487 22431 34493
rect 22462 34484 22468 34496
rect 22520 34484 22526 34536
rect 27080 34533 27108 34564
rect 27154 34552 27160 34604
rect 27212 34592 27218 34604
rect 27249 34595 27307 34601
rect 27249 34592 27261 34595
rect 27212 34564 27261 34592
rect 27212 34552 27218 34564
rect 27249 34561 27261 34564
rect 27295 34561 27307 34595
rect 27890 34592 27896 34604
rect 27851 34564 27896 34592
rect 27249 34555 27307 34561
rect 27890 34552 27896 34564
rect 27948 34552 27954 34604
rect 28000 34601 28028 34632
rect 30926 34620 30932 34672
rect 30984 34660 30990 34672
rect 32858 34660 32864 34672
rect 30984 34632 32864 34660
rect 30984 34620 30990 34632
rect 27985 34595 28043 34601
rect 27985 34561 27997 34595
rect 28031 34561 28043 34595
rect 28350 34592 28356 34604
rect 27985 34555 28043 34561
rect 28184 34564 28356 34592
rect 28184 34533 28212 34564
rect 28350 34552 28356 34564
rect 28408 34552 28414 34604
rect 28626 34592 28632 34604
rect 28587 34564 28632 34592
rect 28626 34552 28632 34564
rect 28684 34552 28690 34604
rect 28813 34595 28871 34601
rect 28813 34561 28825 34595
rect 28859 34592 28871 34595
rect 29825 34595 29883 34601
rect 29825 34592 29837 34595
rect 28859 34564 29837 34592
rect 28859 34561 28871 34564
rect 28813 34555 28871 34561
rect 29825 34561 29837 34564
rect 29871 34592 29883 34595
rect 29914 34592 29920 34604
rect 29871 34564 29920 34592
rect 29871 34561 29883 34564
rect 29825 34555 29883 34561
rect 25409 34527 25467 34533
rect 25409 34493 25421 34527
rect 25455 34524 25467 34527
rect 26329 34527 26387 34533
rect 26329 34524 26341 34527
rect 25455 34496 26341 34524
rect 25455 34493 25467 34496
rect 25409 34487 25467 34493
rect 26329 34493 26341 34496
rect 26375 34493 26387 34527
rect 26329 34487 26387 34493
rect 27065 34527 27123 34533
rect 27065 34493 27077 34527
rect 27111 34493 27123 34527
rect 27065 34487 27123 34493
rect 28169 34527 28227 34533
rect 28169 34493 28181 34527
rect 28215 34493 28227 34527
rect 28828 34524 28856 34555
rect 29914 34552 29920 34564
rect 29972 34552 29978 34604
rect 30009 34595 30067 34601
rect 30009 34561 30021 34595
rect 30055 34592 30067 34595
rect 30098 34592 30104 34604
rect 30055 34564 30104 34592
rect 30055 34561 30067 34564
rect 30009 34555 30067 34561
rect 30098 34552 30104 34564
rect 30156 34552 30162 34604
rect 31312 34601 31340 34632
rect 32858 34620 32864 34632
rect 32916 34620 32922 34672
rect 31205 34595 31263 34601
rect 31205 34592 31217 34595
rect 30208 34564 31217 34592
rect 30208 34524 30236 34564
rect 31205 34561 31217 34564
rect 31251 34561 31263 34595
rect 31205 34555 31263 34561
rect 31297 34595 31355 34601
rect 31297 34561 31309 34595
rect 31343 34561 31355 34595
rect 31573 34595 31631 34601
rect 31573 34592 31585 34595
rect 31297 34555 31355 34561
rect 31404 34564 31585 34592
rect 28169 34487 28227 34493
rect 28276 34496 28856 34524
rect 28920 34496 30236 34524
rect 19300 34428 19472 34456
rect 26344 34456 26372 34487
rect 28276 34456 28304 34496
rect 26344 34428 28304 34456
rect 19300 34416 19306 34428
rect 28350 34416 28356 34468
rect 28408 34456 28414 34468
rect 28920 34456 28948 34496
rect 30282 34484 30288 34536
rect 30340 34524 30346 34536
rect 31404 34524 31432 34564
rect 31573 34561 31585 34564
rect 31619 34561 31631 34595
rect 48130 34592 48136 34604
rect 48091 34564 48136 34592
rect 31573 34555 31631 34561
rect 48130 34552 48136 34564
rect 48188 34552 48194 34604
rect 30340 34496 31432 34524
rect 31481 34527 31539 34533
rect 30340 34484 30346 34496
rect 31481 34493 31493 34527
rect 31527 34524 31539 34527
rect 46566 34524 46572 34536
rect 31527 34496 46572 34524
rect 31527 34493 31539 34496
rect 31481 34487 31539 34493
rect 46566 34484 46572 34496
rect 46624 34484 46630 34536
rect 28408 34428 28948 34456
rect 28408 34416 28414 34428
rect 16942 34388 16948 34400
rect 16903 34360 16948 34388
rect 16942 34348 16948 34360
rect 17000 34348 17006 34400
rect 18414 34388 18420 34400
rect 18375 34360 18420 34388
rect 18414 34348 18420 34360
rect 18472 34388 18478 34400
rect 19061 34391 19119 34397
rect 19061 34388 19073 34391
rect 18472 34360 19073 34388
rect 18472 34348 18478 34360
rect 19061 34357 19073 34360
rect 19107 34357 19119 34391
rect 19061 34351 19119 34357
rect 20441 34391 20499 34397
rect 20441 34357 20453 34391
rect 20487 34388 20499 34391
rect 21726 34388 21732 34400
rect 20487 34360 21732 34388
rect 20487 34357 20499 34360
rect 20441 34351 20499 34357
rect 21726 34348 21732 34360
rect 21784 34348 21790 34400
rect 26142 34348 26148 34400
rect 26200 34388 26206 34400
rect 27154 34388 27160 34400
rect 26200 34360 27160 34388
rect 26200 34348 26206 34360
rect 27154 34348 27160 34360
rect 27212 34348 27218 34400
rect 27430 34388 27436 34400
rect 27391 34360 27436 34388
rect 27430 34348 27436 34360
rect 27488 34348 27494 34400
rect 27890 34348 27896 34400
rect 27948 34388 27954 34400
rect 28994 34388 29000 34400
rect 27948 34360 29000 34388
rect 27948 34348 27954 34360
rect 28994 34348 29000 34360
rect 29052 34348 29058 34400
rect 31021 34391 31079 34397
rect 31021 34357 31033 34391
rect 31067 34388 31079 34391
rect 31202 34388 31208 34400
rect 31067 34360 31208 34388
rect 31067 34357 31079 34360
rect 31021 34351 31079 34357
rect 31202 34348 31208 34360
rect 31260 34348 31266 34400
rect 47210 34348 47216 34400
rect 47268 34388 47274 34400
rect 47949 34391 48007 34397
rect 47949 34388 47961 34391
rect 47268 34360 47961 34388
rect 47268 34348 47274 34360
rect 47949 34357 47961 34360
rect 47995 34357 48007 34391
rect 47949 34351 48007 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 17954 34184 17960 34196
rect 17915 34156 17960 34184
rect 17954 34144 17960 34156
rect 18012 34144 18018 34196
rect 19429 34187 19487 34193
rect 19429 34153 19441 34187
rect 19475 34184 19487 34187
rect 19475 34156 20760 34184
rect 19475 34153 19487 34156
rect 19429 34147 19487 34153
rect 18138 34076 18144 34128
rect 18196 34116 18202 34128
rect 19613 34119 19671 34125
rect 19613 34116 19625 34119
rect 18196 34088 19625 34116
rect 18196 34076 18202 34088
rect 19613 34085 19625 34088
rect 19659 34085 19671 34119
rect 19613 34079 19671 34085
rect 15933 34051 15991 34057
rect 15933 34017 15945 34051
rect 15979 34048 15991 34051
rect 16942 34048 16948 34060
rect 15979 34020 16948 34048
rect 15979 34017 15991 34020
rect 15933 34011 15991 34017
rect 16942 34008 16948 34020
rect 17000 34008 17006 34060
rect 17405 34051 17463 34057
rect 17405 34017 17417 34051
rect 17451 34048 17463 34051
rect 17451 34020 18276 34048
rect 17451 34017 17463 34020
rect 17405 34011 17463 34017
rect 18248 33992 18276 34020
rect 1302 33940 1308 33992
rect 1360 33980 1366 33992
rect 1581 33983 1639 33989
rect 1581 33980 1593 33983
rect 1360 33952 1593 33980
rect 1360 33940 1366 33952
rect 1581 33949 1593 33952
rect 1627 33949 1639 33983
rect 15654 33980 15660 33992
rect 15615 33952 15660 33980
rect 1581 33943 1639 33949
rect 15654 33940 15660 33952
rect 15712 33940 15718 33992
rect 18138 33980 18144 33992
rect 18099 33952 18144 33980
rect 18138 33940 18144 33952
rect 18196 33940 18202 33992
rect 18230 33940 18236 33992
rect 18288 33980 18294 33992
rect 18325 33983 18383 33989
rect 18325 33980 18337 33983
rect 18288 33952 18337 33980
rect 18288 33940 18294 33952
rect 18325 33949 18337 33952
rect 18371 33949 18383 33983
rect 18325 33943 18383 33949
rect 18417 33983 18475 33989
rect 18417 33949 18429 33983
rect 18463 33980 18475 33983
rect 18598 33980 18604 33992
rect 18463 33952 18604 33980
rect 18463 33949 18475 33952
rect 18417 33943 18475 33949
rect 18598 33940 18604 33952
rect 18656 33940 18662 33992
rect 16022 33872 16028 33924
rect 16080 33912 16086 33924
rect 19245 33915 19303 33921
rect 16080 33884 16422 33912
rect 16080 33872 16086 33884
rect 19245 33881 19257 33915
rect 19291 33912 19303 33915
rect 19334 33912 19340 33924
rect 19291 33884 19340 33912
rect 19291 33881 19303 33884
rect 19245 33875 19303 33881
rect 19334 33872 19340 33884
rect 19392 33872 19398 33924
rect 1397 33847 1455 33853
rect 1397 33813 1409 33847
rect 1443 33844 1455 33847
rect 1578 33844 1584 33856
rect 1443 33816 1584 33844
rect 1443 33813 1455 33816
rect 1397 33807 1455 33813
rect 1578 33804 1584 33816
rect 1636 33804 1642 33856
rect 18598 33804 18604 33856
rect 18656 33844 18662 33856
rect 19445 33847 19503 33853
rect 19445 33844 19457 33847
rect 18656 33816 19457 33844
rect 18656 33804 18662 33816
rect 19445 33813 19457 33816
rect 19491 33813 19503 33847
rect 20732 33844 20760 34156
rect 20990 34144 20996 34196
rect 21048 34184 21054 34196
rect 21361 34187 21419 34193
rect 21361 34184 21373 34187
rect 21048 34156 21373 34184
rect 21048 34144 21054 34156
rect 21361 34153 21373 34156
rect 21407 34153 21419 34187
rect 21726 34184 21732 34196
rect 21687 34156 21732 34184
rect 21361 34147 21419 34153
rect 21726 34144 21732 34156
rect 21784 34144 21790 34196
rect 22370 34144 22376 34196
rect 22428 34184 22434 34196
rect 22465 34187 22523 34193
rect 22465 34184 22477 34187
rect 22428 34156 22477 34184
rect 22428 34144 22434 34156
rect 22465 34153 22477 34156
rect 22511 34153 22523 34187
rect 22465 34147 22523 34153
rect 22830 34144 22836 34196
rect 22888 34184 22894 34196
rect 24949 34187 25007 34193
rect 24949 34184 24961 34187
rect 22888 34156 24961 34184
rect 22888 34144 22894 34156
rect 24949 34153 24961 34156
rect 24995 34184 25007 34187
rect 27798 34184 27804 34196
rect 24995 34156 27804 34184
rect 24995 34153 25007 34156
rect 24949 34147 25007 34153
rect 27798 34144 27804 34156
rect 27856 34184 27862 34196
rect 30282 34184 30288 34196
rect 27856 34156 30288 34184
rect 27856 34144 27862 34156
rect 30282 34144 30288 34156
rect 30340 34144 30346 34196
rect 31018 34184 31024 34196
rect 30979 34156 31024 34184
rect 31018 34144 31024 34156
rect 31076 34144 31082 34196
rect 31294 34144 31300 34196
rect 31352 34184 31358 34196
rect 31389 34187 31447 34193
rect 31389 34184 31401 34187
rect 31352 34156 31401 34184
rect 31352 34144 31358 34156
rect 31389 34153 31401 34156
rect 31435 34153 31447 34187
rect 31389 34147 31447 34153
rect 27525 34119 27583 34125
rect 27525 34085 27537 34119
rect 27571 34116 27583 34119
rect 28074 34116 28080 34128
rect 27571 34088 28080 34116
rect 27571 34085 27583 34088
rect 27525 34079 27583 34085
rect 28074 34076 28080 34088
rect 28132 34116 28138 34128
rect 28350 34116 28356 34128
rect 28132 34088 28356 34116
rect 28132 34076 28138 34088
rect 28350 34076 28356 34088
rect 28408 34076 28414 34128
rect 46106 34076 46112 34128
rect 46164 34116 46170 34128
rect 46164 34088 47440 34116
rect 46164 34076 46170 34088
rect 22278 34048 22284 34060
rect 21560 34020 22284 34048
rect 21560 33989 21588 34020
rect 22278 34008 22284 34020
rect 22336 34008 22342 34060
rect 27430 34048 27436 34060
rect 26068 34020 27436 34048
rect 21545 33983 21603 33989
rect 21545 33949 21557 33983
rect 21591 33949 21603 33983
rect 21545 33943 21603 33949
rect 21821 33983 21879 33989
rect 21821 33949 21833 33983
rect 21867 33949 21879 33983
rect 21821 33943 21879 33949
rect 21082 33872 21088 33924
rect 21140 33912 21146 33924
rect 21836 33912 21864 33943
rect 23474 33940 23480 33992
rect 23532 33980 23538 33992
rect 26068 33989 26096 34020
rect 27430 34008 27436 34020
rect 27488 34008 27494 34060
rect 27890 34008 27896 34060
rect 27948 34048 27954 34060
rect 31481 34051 31539 34057
rect 31481 34048 31493 34051
rect 27948 34020 31493 34048
rect 27948 34008 27954 34020
rect 31481 34017 31493 34020
rect 31527 34017 31539 34051
rect 47118 34048 47124 34060
rect 47079 34020 47124 34048
rect 31481 34011 31539 34017
rect 47118 34008 47124 34020
rect 47176 34008 47182 34060
rect 47412 34057 47440 34088
rect 47397 34051 47455 34057
rect 47397 34017 47409 34051
rect 47443 34017 47455 34051
rect 47397 34011 47455 34017
rect 23661 33983 23719 33989
rect 23661 33980 23673 33983
rect 23532 33952 23673 33980
rect 23532 33940 23538 33952
rect 23661 33949 23673 33952
rect 23707 33949 23719 33983
rect 23661 33943 23719 33949
rect 26053 33983 26111 33989
rect 26053 33949 26065 33983
rect 26099 33949 26111 33983
rect 26053 33943 26111 33949
rect 26237 33983 26295 33989
rect 26237 33949 26249 33983
rect 26283 33980 26295 33983
rect 26786 33980 26792 33992
rect 26283 33952 26792 33980
rect 26283 33949 26295 33952
rect 26237 33943 26295 33949
rect 26786 33940 26792 33952
rect 26844 33980 26850 33992
rect 27246 33980 27252 33992
rect 26844 33952 27252 33980
rect 26844 33940 26850 33952
rect 27246 33940 27252 33952
rect 27304 33940 27310 33992
rect 27614 33940 27620 33992
rect 27672 33980 27678 33992
rect 27985 33983 28043 33989
rect 27985 33980 27997 33983
rect 27672 33952 27997 33980
rect 27672 33940 27678 33952
rect 27985 33949 27997 33952
rect 28031 33949 28043 33983
rect 27985 33943 28043 33949
rect 28169 33983 28227 33989
rect 28169 33949 28181 33983
rect 28215 33949 28227 33983
rect 29914 33980 29920 33992
rect 29875 33952 29920 33980
rect 28169 33943 28227 33949
rect 21140 33884 21864 33912
rect 22373 33915 22431 33921
rect 21140 33872 21146 33884
rect 22373 33881 22385 33915
rect 22419 33912 22431 33915
rect 23290 33912 23296 33924
rect 22419 33884 23296 33912
rect 22419 33881 22431 33884
rect 22373 33875 22431 33881
rect 23290 33872 23296 33884
rect 23348 33872 23354 33924
rect 24578 33872 24584 33924
rect 24636 33912 24642 33924
rect 24857 33915 24915 33921
rect 24857 33912 24869 33915
rect 24636 33884 24869 33912
rect 24636 33872 24642 33884
rect 24857 33881 24869 33884
rect 24903 33881 24915 33915
rect 24857 33875 24915 33881
rect 26510 33872 26516 33924
rect 26568 33912 26574 33924
rect 27341 33915 27399 33921
rect 27341 33912 27353 33915
rect 26568 33884 27353 33912
rect 26568 33872 26574 33884
rect 27341 33881 27353 33884
rect 27387 33881 27399 33915
rect 27341 33875 27399 33881
rect 27522 33872 27528 33924
rect 27580 33912 27586 33924
rect 28184 33912 28212 33943
rect 29914 33940 29920 33952
rect 29972 33940 29978 33992
rect 30098 33980 30104 33992
rect 30059 33952 30104 33980
rect 30098 33940 30104 33952
rect 30156 33940 30162 33992
rect 31202 33980 31208 33992
rect 31163 33952 31208 33980
rect 31202 33940 31208 33952
rect 31260 33940 31266 33992
rect 31941 33983 31999 33989
rect 31941 33949 31953 33983
rect 31987 33949 31999 33983
rect 32122 33980 32128 33992
rect 32083 33952 32128 33980
rect 31941 33943 31999 33949
rect 27580 33884 28212 33912
rect 30009 33915 30067 33921
rect 27580 33872 27586 33884
rect 30009 33881 30021 33915
rect 30055 33912 30067 33915
rect 31956 33912 31984 33943
rect 32122 33940 32128 33952
rect 32180 33940 32186 33992
rect 30055 33884 31984 33912
rect 30055 33881 30067 33884
rect 30009 33875 30067 33881
rect 47210 33872 47216 33924
rect 47268 33912 47274 33924
rect 47268 33884 47313 33912
rect 47268 33872 47274 33884
rect 22462 33844 22468 33856
rect 20732 33816 22468 33844
rect 19445 33807 19503 33813
rect 22462 33804 22468 33816
rect 22520 33804 22526 33856
rect 23750 33844 23756 33856
rect 23711 33816 23756 33844
rect 23750 33804 23756 33816
rect 23808 33804 23814 33856
rect 26142 33844 26148 33856
rect 26103 33816 26148 33844
rect 26142 33804 26148 33816
rect 26200 33804 26206 33856
rect 27982 33804 27988 33856
rect 28040 33844 28046 33856
rect 28077 33847 28135 33853
rect 28077 33844 28089 33847
rect 28040 33816 28089 33844
rect 28040 33804 28046 33816
rect 28077 33813 28089 33816
rect 28123 33813 28135 33847
rect 28077 33807 28135 33813
rect 30834 33804 30840 33856
rect 30892 33844 30898 33856
rect 32033 33847 32091 33853
rect 32033 33844 32045 33847
rect 30892 33816 32045 33844
rect 30892 33804 30898 33816
rect 32033 33813 32045 33816
rect 32079 33813 32091 33847
rect 32033 33807 32091 33813
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 16022 33640 16028 33652
rect 15983 33612 16028 33640
rect 16022 33600 16028 33612
rect 16080 33600 16086 33652
rect 17126 33600 17132 33652
rect 17184 33640 17190 33652
rect 17681 33643 17739 33649
rect 17681 33640 17693 33643
rect 17184 33612 17693 33640
rect 17184 33600 17190 33612
rect 17681 33609 17693 33612
rect 17727 33609 17739 33643
rect 18598 33640 18604 33652
rect 18559 33612 18604 33640
rect 17681 33603 17739 33609
rect 18598 33600 18604 33612
rect 18656 33600 18662 33652
rect 19242 33640 19248 33652
rect 19203 33612 19248 33640
rect 19242 33600 19248 33612
rect 19300 33600 19306 33652
rect 22830 33600 22836 33652
rect 22888 33600 22894 33652
rect 26142 33600 26148 33652
rect 26200 33649 26206 33652
rect 26200 33643 26219 33649
rect 26207 33609 26219 33643
rect 26326 33640 26332 33652
rect 26287 33612 26332 33640
rect 26200 33603 26219 33609
rect 26200 33600 26206 33603
rect 26326 33600 26332 33612
rect 26384 33600 26390 33652
rect 28534 33640 28540 33652
rect 28495 33612 28540 33640
rect 28534 33600 28540 33612
rect 28592 33600 28598 33652
rect 32122 33640 32128 33652
rect 30944 33612 32128 33640
rect 17405 33575 17463 33581
rect 17405 33541 17417 33575
rect 17451 33572 17463 33575
rect 18138 33572 18144 33584
rect 17451 33544 18144 33572
rect 17451 33541 17463 33544
rect 17405 33535 17463 33541
rect 18138 33532 18144 33544
rect 18196 33532 18202 33584
rect 18230 33532 18236 33584
rect 18288 33572 18294 33584
rect 22189 33575 22247 33581
rect 18288 33544 18736 33572
rect 18288 33532 18294 33544
rect 15933 33507 15991 33513
rect 15933 33473 15945 33507
rect 15979 33504 15991 33507
rect 16666 33504 16672 33516
rect 15979 33476 16672 33504
rect 15979 33473 15991 33476
rect 15933 33467 15991 33473
rect 16666 33464 16672 33476
rect 16724 33464 16730 33516
rect 17129 33507 17187 33513
rect 17129 33504 17141 33507
rect 16960 33476 17141 33504
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 1670 33436 1676 33448
rect 1631 33408 1676 33436
rect 1670 33396 1676 33408
rect 1728 33396 1734 33448
rect 16960 33368 16988 33476
rect 17129 33473 17141 33476
rect 17175 33473 17187 33507
rect 17310 33504 17316 33516
rect 17271 33476 17316 33504
rect 17129 33467 17187 33473
rect 17310 33464 17316 33476
rect 17368 33464 17374 33516
rect 17497 33507 17555 33513
rect 17497 33473 17509 33507
rect 17543 33473 17555 33507
rect 18506 33504 18512 33516
rect 18467 33476 18512 33504
rect 17497 33467 17555 33473
rect 17034 33396 17040 33448
rect 17092 33436 17098 33448
rect 17512 33436 17540 33467
rect 18506 33464 18512 33476
rect 18564 33464 18570 33516
rect 18708 33513 18736 33544
rect 22189 33541 22201 33575
rect 22235 33572 22247 33575
rect 22848 33572 22876 33600
rect 22235 33544 22876 33572
rect 22235 33541 22247 33544
rect 22189 33535 22247 33541
rect 23750 33532 23756 33584
rect 23808 33532 23814 33584
rect 25961 33575 26019 33581
rect 25961 33572 25973 33575
rect 25424 33544 25973 33572
rect 18693 33507 18751 33513
rect 18693 33473 18705 33507
rect 18739 33473 18751 33507
rect 18693 33467 18751 33473
rect 18966 33464 18972 33516
rect 19024 33504 19030 33516
rect 19153 33507 19211 33513
rect 19153 33504 19165 33507
rect 19024 33476 19165 33504
rect 19024 33464 19030 33476
rect 19153 33473 19165 33476
rect 19199 33473 19211 33507
rect 19334 33504 19340 33516
rect 19295 33476 19340 33504
rect 19153 33467 19211 33473
rect 19334 33464 19340 33476
rect 19392 33464 19398 33516
rect 22370 33464 22376 33516
rect 22428 33504 22434 33516
rect 22833 33507 22891 33513
rect 22833 33504 22845 33507
rect 22428 33476 22845 33504
rect 22428 33464 22434 33476
rect 22833 33473 22845 33476
rect 22879 33473 22891 33507
rect 22833 33467 22891 33473
rect 24946 33464 24952 33516
rect 25004 33504 25010 33516
rect 25424 33513 25452 33544
rect 25961 33541 25973 33544
rect 26007 33541 26019 33575
rect 26970 33572 26976 33584
rect 26883 33544 26976 33572
rect 25961 33535 26019 33541
rect 26970 33532 26976 33544
rect 27028 33572 27034 33584
rect 27430 33572 27436 33584
rect 27028 33544 27436 33572
rect 27028 33532 27034 33544
rect 27430 33532 27436 33544
rect 27488 33532 27494 33584
rect 30944 33581 30972 33612
rect 32122 33600 32128 33612
rect 32180 33600 32186 33652
rect 30929 33575 30987 33581
rect 30929 33541 30941 33575
rect 30975 33541 30987 33575
rect 30929 33535 30987 33541
rect 31021 33575 31079 33581
rect 31021 33541 31033 33575
rect 31067 33572 31079 33575
rect 32766 33572 32772 33584
rect 31067 33544 32772 33572
rect 31067 33541 31079 33544
rect 31021 33535 31079 33541
rect 25409 33507 25467 33513
rect 25409 33504 25421 33507
rect 25004 33476 25421 33504
rect 25004 33464 25010 33476
rect 25409 33473 25421 33476
rect 25455 33473 25467 33507
rect 25409 33467 25467 33473
rect 25501 33507 25559 33513
rect 25501 33473 25513 33507
rect 25547 33504 25559 33507
rect 25590 33504 25596 33516
rect 25547 33476 25596 33504
rect 25547 33473 25559 33476
rect 25501 33467 25559 33473
rect 25590 33464 25596 33476
rect 25648 33504 25654 33516
rect 25866 33504 25872 33516
rect 25648 33476 25872 33504
rect 25648 33464 25654 33476
rect 25866 33464 25872 33476
rect 25924 33464 25930 33516
rect 27154 33504 27160 33516
rect 27115 33476 27160 33504
rect 27154 33464 27160 33476
rect 27212 33464 27218 33516
rect 28442 33504 28448 33516
rect 28403 33476 28448 33504
rect 28442 33464 28448 33476
rect 28500 33464 28506 33516
rect 29089 33507 29147 33513
rect 29089 33473 29101 33507
rect 29135 33473 29147 33507
rect 30650 33504 30656 33516
rect 30611 33476 30656 33504
rect 29089 33467 29147 33473
rect 23106 33436 23112 33448
rect 17092 33408 17540 33436
rect 23067 33408 23112 33436
rect 17092 33396 17098 33408
rect 23106 33396 23112 33408
rect 23164 33396 23170 33448
rect 24581 33439 24639 33445
rect 24581 33405 24593 33439
rect 24627 33436 24639 33439
rect 25038 33436 25044 33448
rect 24627 33408 25044 33436
rect 24627 33405 24639 33408
rect 24581 33399 24639 33405
rect 25038 33396 25044 33408
rect 25096 33396 25102 33448
rect 26878 33396 26884 33448
rect 26936 33436 26942 33448
rect 29104 33436 29132 33467
rect 30650 33464 30656 33476
rect 30708 33464 30714 33516
rect 30834 33513 30840 33516
rect 30801 33507 30840 33513
rect 30801 33473 30813 33507
rect 30801 33467 30840 33473
rect 30834 33464 30840 33467
rect 30892 33464 30898 33516
rect 26936 33408 29132 33436
rect 26936 33396 26942 33408
rect 30098 33396 30104 33448
rect 30156 33436 30162 33448
rect 31036 33436 31064 33535
rect 32766 33532 32772 33544
rect 32824 33532 32830 33584
rect 31202 33513 31208 33516
rect 31159 33507 31208 33513
rect 31159 33473 31171 33507
rect 31205 33473 31208 33507
rect 31159 33467 31208 33473
rect 31202 33464 31208 33467
rect 31260 33464 31266 33516
rect 31846 33464 31852 33516
rect 31904 33504 31910 33516
rect 32125 33507 32183 33513
rect 32125 33504 32137 33507
rect 31904 33476 32137 33504
rect 31904 33464 31910 33476
rect 32125 33473 32137 33476
rect 32171 33473 32183 33507
rect 47762 33504 47768 33516
rect 47723 33476 47768 33504
rect 32125 33467 32183 33473
rect 47762 33464 47768 33476
rect 47820 33464 47826 33516
rect 48041 33439 48099 33445
rect 48041 33436 48053 33439
rect 30156 33408 31064 33436
rect 31726 33408 48053 33436
rect 30156 33396 30162 33408
rect 18230 33368 18236 33380
rect 16960 33340 18236 33368
rect 18230 33328 18236 33340
rect 18288 33328 18294 33380
rect 19426 33328 19432 33380
rect 19484 33368 19490 33380
rect 31726 33368 31754 33408
rect 48041 33405 48053 33408
rect 48087 33405 48099 33439
rect 48041 33399 48099 33405
rect 19484 33340 22968 33368
rect 19484 33328 19490 33340
rect 18506 33260 18512 33312
rect 18564 33300 18570 33312
rect 18690 33300 18696 33312
rect 18564 33272 18696 33300
rect 18564 33260 18570 33272
rect 18690 33260 18696 33272
rect 18748 33260 18754 33312
rect 22278 33300 22284 33312
rect 22239 33272 22284 33300
rect 22278 33260 22284 33272
rect 22336 33260 22342 33312
rect 22940 33300 22968 33340
rect 24228 33340 31754 33368
rect 23750 33300 23756 33312
rect 22940 33272 23756 33300
rect 23750 33260 23756 33272
rect 23808 33300 23814 33312
rect 24228 33300 24256 33340
rect 25222 33300 25228 33312
rect 23808 33272 24256 33300
rect 25183 33272 25228 33300
rect 23808 33260 23814 33272
rect 25222 33260 25228 33272
rect 25280 33260 25286 33312
rect 26142 33300 26148 33312
rect 26103 33272 26148 33300
rect 26142 33260 26148 33272
rect 26200 33260 26206 33312
rect 26510 33260 26516 33312
rect 26568 33300 26574 33312
rect 27341 33303 27399 33309
rect 27341 33300 27353 33303
rect 26568 33272 27353 33300
rect 26568 33260 26574 33272
rect 27341 33269 27353 33272
rect 27387 33300 27399 33303
rect 27522 33300 27528 33312
rect 27387 33272 27528 33300
rect 27387 33269 27399 33272
rect 27341 33263 27399 33269
rect 27522 33260 27528 33272
rect 27580 33260 27586 33312
rect 29178 33300 29184 33312
rect 29139 33272 29184 33300
rect 29178 33260 29184 33272
rect 29236 33260 29242 33312
rect 31294 33300 31300 33312
rect 31255 33272 31300 33300
rect 31294 33260 31300 33272
rect 31352 33260 31358 33312
rect 32217 33303 32275 33309
rect 32217 33269 32229 33303
rect 32263 33300 32275 33303
rect 32306 33300 32312 33312
rect 32263 33272 32312 33300
rect 32263 33269 32275 33272
rect 32217 33263 32275 33269
rect 32306 33260 32312 33272
rect 32364 33260 32370 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 17494 33056 17500 33108
rect 17552 33096 17558 33108
rect 22278 33096 22284 33108
rect 17552 33068 22284 33096
rect 17552 33056 17558 33068
rect 22278 33056 22284 33068
rect 22336 33056 22342 33108
rect 22741 33099 22799 33105
rect 22741 33065 22753 33099
rect 22787 33096 22799 33099
rect 23014 33096 23020 33108
rect 22787 33068 23020 33096
rect 22787 33065 22799 33068
rect 22741 33059 22799 33065
rect 23014 33056 23020 33068
rect 23072 33056 23078 33108
rect 25222 33056 25228 33108
rect 25280 33096 25286 33108
rect 25593 33099 25651 33105
rect 25593 33096 25605 33099
rect 25280 33068 25605 33096
rect 25280 33056 25286 33068
rect 25593 33065 25605 33068
rect 25639 33065 25651 33099
rect 25593 33059 25651 33065
rect 25685 33099 25743 33105
rect 25685 33065 25697 33099
rect 25731 33096 25743 33099
rect 26326 33096 26332 33108
rect 25731 33068 26332 33096
rect 25731 33065 25743 33068
rect 25685 33059 25743 33065
rect 26326 33056 26332 33068
rect 26384 33056 26390 33108
rect 26786 33096 26792 33108
rect 26747 33068 26792 33096
rect 26786 33056 26792 33068
rect 26844 33056 26850 33108
rect 28166 33056 28172 33108
rect 28224 33096 28230 33108
rect 28997 33099 29055 33105
rect 28997 33096 29009 33099
rect 28224 33068 29009 33096
rect 28224 33056 28230 33068
rect 28997 33065 29009 33068
rect 29043 33065 29055 33099
rect 28997 33059 29055 33065
rect 30098 33056 30104 33108
rect 30156 33096 30162 33108
rect 31846 33096 31852 33108
rect 30156 33068 31852 33096
rect 30156 33056 30162 33068
rect 31846 33056 31852 33068
rect 31904 33056 31910 33108
rect 32766 33096 32772 33108
rect 32727 33068 32772 33096
rect 32766 33056 32772 33068
rect 32824 33056 32830 33108
rect 1486 33028 1492 33040
rect 1412 33000 1492 33028
rect 1412 32969 1440 33000
rect 1486 32988 1492 33000
rect 1544 32988 1550 33040
rect 16666 32988 16672 33040
rect 16724 33028 16730 33040
rect 23109 33031 23167 33037
rect 23109 33028 23121 33031
rect 16724 33000 21404 33028
rect 16724 32988 16730 33000
rect 1397 32963 1455 32969
rect 1397 32929 1409 32963
rect 1443 32929 1455 32963
rect 1578 32960 1584 32972
rect 1539 32932 1584 32960
rect 1397 32923 1455 32929
rect 1578 32920 1584 32932
rect 1636 32920 1642 32972
rect 12526 32920 12532 32972
rect 12584 32960 12590 32972
rect 18414 32960 18420 32972
rect 12584 32932 18420 32960
rect 12584 32920 12590 32932
rect 18414 32920 18420 32932
rect 18472 32920 18478 32972
rect 20806 32960 20812 32972
rect 18524 32932 20812 32960
rect 18524 32904 18552 32932
rect 20806 32920 20812 32932
rect 20864 32920 20870 32972
rect 16761 32895 16819 32901
rect 16761 32861 16773 32895
rect 16807 32892 16819 32895
rect 17405 32895 17463 32901
rect 17405 32892 17417 32895
rect 16807 32864 17417 32892
rect 16807 32861 16819 32864
rect 16761 32855 16819 32861
rect 17405 32861 17417 32864
rect 17451 32892 17463 32895
rect 18230 32892 18236 32904
rect 17451 32864 18236 32892
rect 17451 32861 17463 32864
rect 17405 32855 17463 32861
rect 18230 32852 18236 32864
rect 18288 32852 18294 32904
rect 18506 32892 18512 32904
rect 18467 32864 18512 32892
rect 18506 32852 18512 32864
rect 18564 32852 18570 32904
rect 18598 32852 18604 32904
rect 18656 32892 18662 32904
rect 18693 32895 18751 32901
rect 18693 32892 18705 32895
rect 18656 32864 18705 32892
rect 18656 32852 18662 32864
rect 18693 32861 18705 32864
rect 18739 32861 18751 32895
rect 18693 32855 18751 32861
rect 18874 32852 18880 32904
rect 18932 32892 18938 32904
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18932 32864 19257 32892
rect 18932 32852 18938 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19245 32855 19303 32861
rect 21269 32895 21327 32901
rect 21269 32861 21281 32895
rect 21315 32861 21327 32895
rect 21376 32892 21404 33000
rect 22066 33000 23121 33028
rect 21542 32920 21548 32972
rect 21600 32960 21606 32972
rect 22066 32960 22094 33000
rect 23109 32997 23121 33000
rect 23155 32997 23167 33031
rect 23109 32991 23167 32997
rect 23198 32988 23204 33040
rect 23256 33028 23262 33040
rect 23474 33028 23480 33040
rect 23256 33000 23480 33028
rect 23256 32988 23262 33000
rect 23474 32988 23480 33000
rect 23532 32988 23538 33040
rect 24670 32988 24676 33040
rect 24728 33028 24734 33040
rect 26418 33028 26424 33040
rect 24728 33000 26424 33028
rect 24728 32988 24734 33000
rect 26418 32988 26424 33000
rect 26476 32988 26482 33040
rect 21600 32932 22094 32960
rect 21600 32920 21606 32932
rect 22278 32920 22284 32972
rect 22336 32960 22342 32972
rect 22336 32932 23244 32960
rect 22336 32920 22342 32932
rect 23216 32901 23244 32932
rect 25038 32920 25044 32972
rect 25096 32960 25102 32972
rect 27249 32963 27307 32969
rect 25096 32932 26648 32960
rect 25096 32920 25102 32932
rect 22925 32895 22983 32901
rect 21376 32864 22094 32892
rect 21269 32855 21327 32861
rect 3234 32824 3240 32836
rect 3195 32796 3240 32824
rect 3234 32784 3240 32796
rect 3292 32784 3298 32836
rect 17954 32784 17960 32836
rect 18012 32824 18018 32836
rect 19334 32824 19340 32836
rect 18012 32796 19340 32824
rect 18012 32784 18018 32796
rect 19334 32784 19340 32796
rect 19392 32784 19398 32836
rect 21284 32824 21312 32855
rect 22066 32824 22094 32864
rect 22925 32861 22937 32895
rect 22971 32861 22983 32895
rect 22925 32855 22983 32861
rect 23201 32895 23259 32901
rect 23201 32861 23213 32895
rect 23247 32892 23259 32895
rect 23934 32892 23940 32904
rect 23247 32864 23940 32892
rect 23247 32861 23259 32864
rect 23201 32855 23259 32861
rect 22940 32824 22968 32855
rect 23934 32852 23940 32864
rect 23992 32852 23998 32904
rect 25498 32892 25504 32904
rect 25459 32864 25504 32892
rect 25498 32852 25504 32864
rect 25556 32852 25562 32904
rect 25792 32901 25820 32932
rect 25777 32895 25835 32901
rect 25777 32861 25789 32895
rect 25823 32861 25835 32895
rect 25777 32855 25835 32861
rect 25961 32895 26019 32901
rect 25961 32861 25973 32895
rect 26007 32892 26019 32895
rect 26510 32892 26516 32904
rect 26007 32864 26516 32892
rect 26007 32861 26019 32864
rect 25961 32855 26019 32861
rect 26510 32852 26516 32864
rect 26568 32852 26574 32904
rect 26620 32901 26648 32932
rect 27249 32929 27261 32963
rect 27295 32960 27307 32963
rect 28534 32960 28540 32972
rect 27295 32932 28540 32960
rect 27295 32929 27307 32932
rect 27249 32923 27307 32929
rect 28534 32920 28540 32932
rect 28592 32960 28598 32972
rect 31021 32963 31079 32969
rect 31021 32960 31033 32963
rect 28592 32932 31033 32960
rect 28592 32920 28598 32932
rect 31021 32929 31033 32932
rect 31067 32929 31079 32963
rect 31294 32960 31300 32972
rect 31255 32932 31300 32960
rect 31021 32923 31079 32929
rect 31294 32920 31300 32932
rect 31352 32920 31358 32972
rect 26605 32895 26663 32901
rect 26605 32861 26617 32895
rect 26651 32861 26663 32895
rect 26605 32855 26663 32861
rect 28902 32852 28908 32904
rect 28960 32892 28966 32904
rect 30009 32895 30067 32901
rect 30009 32892 30021 32895
rect 28960 32864 30021 32892
rect 28960 32852 28966 32864
rect 30009 32861 30021 32864
rect 30055 32861 30067 32895
rect 46290 32892 46296 32904
rect 46251 32864 46296 32892
rect 30009 32855 30067 32861
rect 46290 32852 46296 32864
rect 46348 32852 46354 32904
rect 25225 32827 25283 32833
rect 25225 32824 25237 32827
rect 21284 32796 21680 32824
rect 22066 32796 22876 32824
rect 22940 32796 25237 32824
rect 16850 32756 16856 32768
rect 16811 32728 16856 32756
rect 16850 32716 16856 32728
rect 16908 32716 16914 32768
rect 17497 32759 17555 32765
rect 17497 32725 17509 32759
rect 17543 32756 17555 32759
rect 18046 32756 18052 32768
rect 17543 32728 18052 32756
rect 17543 32725 17555 32728
rect 17497 32719 17555 32725
rect 18046 32716 18052 32728
rect 18104 32716 18110 32768
rect 18601 32759 18659 32765
rect 18601 32725 18613 32759
rect 18647 32756 18659 32759
rect 18966 32756 18972 32768
rect 18647 32728 18972 32756
rect 18647 32725 18659 32728
rect 18601 32719 18659 32725
rect 18966 32716 18972 32728
rect 19024 32716 19030 32768
rect 20990 32716 20996 32768
rect 21048 32756 21054 32768
rect 21453 32759 21511 32765
rect 21453 32756 21465 32759
rect 21048 32728 21465 32756
rect 21048 32716 21054 32728
rect 21453 32725 21465 32728
rect 21499 32725 21511 32759
rect 21652 32756 21680 32796
rect 22370 32756 22376 32768
rect 21652 32728 22376 32756
rect 21453 32719 21511 32725
rect 22370 32716 22376 32728
rect 22428 32716 22434 32768
rect 22848 32756 22876 32796
rect 25225 32793 25237 32796
rect 25271 32793 25283 32827
rect 25225 32787 25283 32793
rect 26421 32827 26479 32833
rect 26421 32793 26433 32827
rect 26467 32824 26479 32827
rect 27154 32824 27160 32836
rect 26467 32796 27160 32824
rect 26467 32793 26479 32796
rect 26421 32787 26479 32793
rect 27154 32784 27160 32796
rect 27212 32784 27218 32836
rect 27525 32827 27583 32833
rect 27525 32793 27537 32827
rect 27571 32824 27583 32827
rect 27614 32824 27620 32836
rect 27571 32796 27620 32824
rect 27571 32793 27583 32796
rect 27525 32787 27583 32793
rect 27614 32784 27620 32796
rect 27672 32784 27678 32836
rect 29178 32824 29184 32836
rect 28750 32796 29184 32824
rect 29178 32784 29184 32796
rect 29236 32784 29242 32836
rect 32306 32784 32312 32836
rect 32364 32784 32370 32836
rect 46477 32827 46535 32833
rect 46477 32793 46489 32827
rect 46523 32824 46535 32827
rect 47670 32824 47676 32836
rect 46523 32796 47676 32824
rect 46523 32793 46535 32796
rect 46477 32787 46535 32793
rect 47670 32784 47676 32796
rect 47728 32784 47734 32836
rect 48130 32824 48136 32836
rect 48091 32796 48136 32824
rect 48130 32784 48136 32796
rect 48188 32784 48194 32836
rect 30098 32756 30104 32768
rect 22848 32728 30104 32756
rect 30098 32716 30104 32728
rect 30156 32716 30162 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 18417 32555 18475 32561
rect 18417 32521 18429 32555
rect 18463 32552 18475 32555
rect 18874 32552 18880 32564
rect 18463 32524 18880 32552
rect 18463 32521 18475 32524
rect 18417 32515 18475 32521
rect 18874 32512 18880 32524
rect 18932 32512 18938 32564
rect 19058 32552 19064 32564
rect 19019 32524 19064 32552
rect 19058 32512 19064 32524
rect 19116 32512 19122 32564
rect 20990 32552 20996 32564
rect 19352 32524 20996 32552
rect 1670 32444 1676 32496
rect 1728 32484 1734 32496
rect 2317 32487 2375 32493
rect 2317 32484 2329 32487
rect 1728 32456 2329 32484
rect 1728 32444 1734 32456
rect 2317 32453 2329 32456
rect 2363 32453 2375 32487
rect 2317 32447 2375 32453
rect 16850 32444 16856 32496
rect 16908 32484 16914 32496
rect 16908 32456 17434 32484
rect 16908 32444 16914 32456
rect 18230 32444 18236 32496
rect 18288 32484 18294 32496
rect 19352 32484 19380 32524
rect 20990 32512 20996 32524
rect 21048 32512 21054 32564
rect 22278 32552 22284 32564
rect 21192 32524 22284 32552
rect 18288 32456 19380 32484
rect 18288 32444 18294 32456
rect 19426 32444 19432 32496
rect 19484 32484 19490 32496
rect 20073 32487 20131 32493
rect 20073 32484 20085 32487
rect 19484 32456 20085 32484
rect 19484 32444 19490 32456
rect 20073 32453 20085 32456
rect 20119 32453 20131 32487
rect 21192 32484 21220 32524
rect 22278 32512 22284 32524
rect 22336 32512 22342 32564
rect 25222 32512 25228 32564
rect 25280 32552 25286 32564
rect 25961 32555 26019 32561
rect 25961 32552 25973 32555
rect 25280 32524 25973 32552
rect 25280 32512 25286 32524
rect 25961 32521 25973 32524
rect 26007 32521 26019 32555
rect 27614 32552 27620 32564
rect 27575 32524 27620 32552
rect 25961 32515 26019 32521
rect 27614 32512 27620 32524
rect 27672 32512 27678 32564
rect 30650 32512 30656 32564
rect 30708 32552 30714 32564
rect 30837 32555 30895 32561
rect 30837 32552 30849 32555
rect 30708 32524 30849 32552
rect 30708 32512 30714 32524
rect 30837 32521 30849 32524
rect 30883 32521 30895 32555
rect 47670 32552 47676 32564
rect 47631 32524 47676 32552
rect 30837 32515 30895 32521
rect 47670 32512 47676 32524
rect 47728 32512 47734 32564
rect 23106 32484 23112 32496
rect 20073 32447 20131 32453
rect 21100 32456 21220 32484
rect 22020 32456 23112 32484
rect 15654 32376 15660 32428
rect 15712 32416 15718 32428
rect 21100 32425 21128 32456
rect 22020 32425 22048 32456
rect 23106 32444 23112 32456
rect 23164 32444 23170 32496
rect 25133 32487 25191 32493
rect 25133 32453 25145 32487
rect 25179 32484 25191 32487
rect 25590 32484 25596 32496
rect 25179 32456 25596 32484
rect 25179 32453 25191 32456
rect 25133 32447 25191 32453
rect 25590 32444 25596 32456
rect 25648 32484 25654 32496
rect 26142 32484 26148 32496
rect 25648 32456 26148 32484
rect 25648 32444 25654 32456
rect 26142 32444 26148 32456
rect 26200 32444 26206 32496
rect 27065 32487 27123 32493
rect 27065 32453 27077 32487
rect 27111 32484 27123 32487
rect 27522 32484 27528 32496
rect 27111 32456 27528 32484
rect 27111 32453 27123 32456
rect 27065 32447 27123 32453
rect 27522 32444 27528 32456
rect 27580 32444 27586 32496
rect 27890 32444 27896 32496
rect 27948 32484 27954 32496
rect 27948 32456 28120 32484
rect 27948 32444 27954 32456
rect 16669 32419 16727 32425
rect 16669 32416 16681 32419
rect 15712 32388 16681 32416
rect 15712 32376 15718 32388
rect 16669 32385 16681 32388
rect 16715 32385 16727 32419
rect 16669 32379 16727 32385
rect 19058 32419 19116 32425
rect 19058 32385 19070 32419
rect 19104 32416 19116 32419
rect 21085 32419 21143 32425
rect 19104 32388 19288 32416
rect 19104 32385 19116 32388
rect 19058 32379 19116 32385
rect 2133 32351 2191 32357
rect 2133 32317 2145 32351
rect 2179 32348 2191 32351
rect 2406 32348 2412 32360
rect 2179 32320 2412 32348
rect 2179 32317 2191 32320
rect 2133 32311 2191 32317
rect 2406 32308 2412 32320
rect 2464 32308 2470 32360
rect 3234 32348 3240 32360
rect 3195 32320 3240 32348
rect 3234 32308 3240 32320
rect 3292 32308 3298 32360
rect 16942 32348 16948 32360
rect 16903 32320 16948 32348
rect 16942 32308 16948 32320
rect 17000 32308 17006 32360
rect 19260 32280 19288 32388
rect 21085 32385 21097 32419
rect 21131 32385 21143 32419
rect 21085 32379 21143 32385
rect 21177 32419 21235 32425
rect 21177 32385 21189 32419
rect 21223 32416 21235 32419
rect 22005 32419 22063 32425
rect 22005 32416 22017 32419
rect 21223 32388 22017 32416
rect 21223 32385 21235 32388
rect 21177 32379 21235 32385
rect 22005 32385 22017 32388
rect 22051 32385 22063 32419
rect 22005 32379 22063 32385
rect 22465 32419 22523 32425
rect 22465 32385 22477 32419
rect 22511 32416 22523 32419
rect 22830 32416 22836 32428
rect 22511 32388 22836 32416
rect 22511 32385 22523 32388
rect 22465 32379 22523 32385
rect 22830 32376 22836 32388
rect 22888 32376 22894 32428
rect 23198 32416 23204 32428
rect 23159 32388 23204 32416
rect 23198 32376 23204 32388
rect 23256 32376 23262 32428
rect 23842 32416 23848 32428
rect 23803 32388 23848 32416
rect 23842 32376 23848 32388
rect 23900 32376 23906 32428
rect 24670 32416 24676 32428
rect 24631 32388 24676 32416
rect 24670 32376 24676 32388
rect 24728 32376 24734 32428
rect 24854 32416 24860 32428
rect 24815 32388 24860 32416
rect 24854 32376 24860 32388
rect 24912 32376 24918 32428
rect 24946 32376 24952 32428
rect 25004 32416 25010 32428
rect 25041 32419 25099 32425
rect 25041 32416 25053 32419
rect 25004 32388 25053 32416
rect 25004 32376 25010 32388
rect 25041 32385 25053 32388
rect 25087 32385 25099 32419
rect 25041 32379 25099 32385
rect 25498 32376 25504 32428
rect 25556 32416 25562 32428
rect 25902 32419 25960 32425
rect 25902 32416 25914 32419
rect 25556 32388 25914 32416
rect 25556 32376 25562 32388
rect 25884 32385 25914 32388
rect 25948 32385 25960 32419
rect 25884 32379 25960 32385
rect 26329 32419 26387 32425
rect 26329 32385 26341 32419
rect 26375 32416 26387 32419
rect 26970 32416 26976 32428
rect 26375 32388 26976 32416
rect 26375 32385 26387 32388
rect 26329 32379 26387 32385
rect 19518 32348 19524 32360
rect 19479 32320 19524 32348
rect 19518 32308 19524 32320
rect 19576 32308 19582 32360
rect 22186 32348 22192 32360
rect 22147 32320 22192 32348
rect 22186 32308 22192 32320
rect 22244 32308 22250 32360
rect 22281 32351 22339 32357
rect 22281 32317 22293 32351
rect 22327 32348 22339 32351
rect 22554 32348 22560 32360
rect 22327 32320 22560 32348
rect 22327 32317 22339 32320
rect 22281 32311 22339 32317
rect 22554 32308 22560 32320
rect 22612 32308 22618 32360
rect 23290 32308 23296 32360
rect 23348 32348 23354 32360
rect 23385 32351 23443 32357
rect 23385 32348 23397 32351
rect 23348 32320 23397 32348
rect 23348 32308 23354 32320
rect 23385 32317 23397 32320
rect 23431 32317 23443 32351
rect 23385 32311 23443 32317
rect 19260 32252 19564 32280
rect 1394 32172 1400 32224
rect 1452 32212 1458 32224
rect 1673 32215 1731 32221
rect 1673 32212 1685 32215
rect 1452 32184 1685 32212
rect 1452 32172 1458 32184
rect 1673 32181 1685 32184
rect 1719 32181 1731 32215
rect 18874 32212 18880 32224
rect 18835 32184 18880 32212
rect 1673 32175 1731 32181
rect 18874 32172 18880 32184
rect 18932 32172 18938 32224
rect 19242 32172 19248 32224
rect 19300 32212 19306 32224
rect 19429 32215 19487 32221
rect 19429 32212 19441 32215
rect 19300 32184 19441 32212
rect 19300 32172 19306 32184
rect 19429 32181 19441 32184
rect 19475 32181 19487 32215
rect 19536 32212 19564 32252
rect 22094 32240 22100 32292
rect 22152 32280 22158 32292
rect 22152 32252 22197 32280
rect 22152 32240 22158 32252
rect 22370 32240 22376 32292
rect 22428 32280 22434 32292
rect 25774 32280 25780 32292
rect 22428 32252 25636 32280
rect 25735 32252 25780 32280
rect 22428 32240 22434 32252
rect 19702 32212 19708 32224
rect 19536 32184 19708 32212
rect 19429 32175 19487 32181
rect 19702 32172 19708 32184
rect 19760 32172 19766 32224
rect 20162 32212 20168 32224
rect 20123 32184 20168 32212
rect 20162 32172 20168 32184
rect 20220 32172 20226 32224
rect 21821 32215 21879 32221
rect 21821 32181 21833 32215
rect 21867 32212 21879 32215
rect 22738 32212 22744 32224
rect 21867 32184 22744 32212
rect 21867 32181 21879 32184
rect 21821 32175 21879 32181
rect 22738 32172 22744 32184
rect 22796 32172 22802 32224
rect 23014 32172 23020 32224
rect 23072 32212 23078 32224
rect 23937 32215 23995 32221
rect 23937 32212 23949 32215
rect 23072 32184 23949 32212
rect 23072 32172 23078 32184
rect 23937 32181 23949 32184
rect 23983 32181 23995 32215
rect 25608 32212 25636 32252
rect 25774 32240 25780 32252
rect 25832 32240 25838 32292
rect 25884 32280 25912 32379
rect 26970 32376 26976 32388
rect 27028 32376 27034 32428
rect 27154 32416 27160 32428
rect 27115 32388 27160 32416
rect 27154 32376 27160 32388
rect 27212 32376 27218 32428
rect 27798 32376 27804 32428
rect 27856 32416 27862 32428
rect 27982 32416 27988 32428
rect 27856 32388 27901 32416
rect 27943 32388 27988 32416
rect 27856 32376 27862 32388
rect 27982 32376 27988 32388
rect 28040 32376 28046 32428
rect 28092 32425 28120 32456
rect 28077 32419 28135 32425
rect 28077 32385 28089 32419
rect 28123 32385 28135 32419
rect 28077 32379 28135 32385
rect 30653 32419 30711 32425
rect 30653 32385 30665 32419
rect 30699 32416 30711 32419
rect 31570 32416 31576 32428
rect 30699 32388 31576 32416
rect 30699 32385 30711 32388
rect 30653 32379 30711 32385
rect 31570 32376 31576 32388
rect 31628 32376 31634 32428
rect 46290 32376 46296 32428
rect 46348 32416 46354 32428
rect 47029 32419 47087 32425
rect 47029 32416 47041 32419
rect 46348 32388 47041 32416
rect 46348 32376 46354 32388
rect 47029 32385 47041 32388
rect 47075 32385 47087 32419
rect 47029 32379 47087 32385
rect 47486 32376 47492 32428
rect 47544 32416 47550 32428
rect 47581 32419 47639 32425
rect 47581 32416 47593 32419
rect 47544 32388 47593 32416
rect 47544 32376 47550 32388
rect 47581 32385 47593 32388
rect 47627 32385 47639 32419
rect 47581 32379 47639 32385
rect 26418 32348 26424 32360
rect 26331 32320 26424 32348
rect 26418 32308 26424 32320
rect 26476 32348 26482 32360
rect 28258 32348 28264 32360
rect 26476 32320 28264 32348
rect 26476 32308 26482 32320
rect 28258 32308 28264 32320
rect 28316 32308 28322 32360
rect 30466 32348 30472 32360
rect 30427 32320 30472 32348
rect 30466 32308 30472 32320
rect 30524 32308 30530 32360
rect 26786 32280 26792 32292
rect 25884 32252 26792 32280
rect 26786 32240 26792 32252
rect 26844 32240 26850 32292
rect 27154 32240 27160 32292
rect 27212 32280 27218 32292
rect 28166 32280 28172 32292
rect 27212 32252 28172 32280
rect 27212 32240 27218 32252
rect 28166 32240 28172 32252
rect 28224 32240 28230 32292
rect 29086 32240 29092 32292
rect 29144 32280 29150 32292
rect 29454 32280 29460 32292
rect 29144 32252 29460 32280
rect 29144 32240 29150 32252
rect 29454 32240 29460 32252
rect 29512 32240 29518 32292
rect 28902 32212 28908 32224
rect 25608 32184 28908 32212
rect 23937 32175 23995 32181
rect 28902 32172 28908 32184
rect 28960 32172 28966 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 16942 31968 16948 32020
rect 17000 32008 17006 32020
rect 18049 32011 18107 32017
rect 18049 32008 18061 32011
rect 17000 31980 18061 32008
rect 17000 31968 17006 31980
rect 18049 31977 18061 31980
rect 18095 31977 18107 32011
rect 20990 32008 20996 32020
rect 18049 31971 18107 31977
rect 19536 31980 20996 32008
rect 17957 31943 18015 31949
rect 17957 31940 17969 31943
rect 17052 31912 17969 31940
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 1854 31872 1860 31884
rect 1815 31844 1860 31872
rect 1854 31832 1860 31844
rect 1912 31832 1918 31884
rect 17052 31813 17080 31912
rect 17957 31909 17969 31912
rect 18003 31940 18015 31943
rect 19245 31943 19303 31949
rect 19245 31940 19257 31943
rect 18003 31912 19257 31940
rect 18003 31909 18015 31912
rect 17957 31903 18015 31909
rect 19245 31909 19257 31912
rect 19291 31909 19303 31943
rect 19245 31903 19303 31909
rect 17310 31872 17316 31884
rect 17271 31844 17316 31872
rect 17310 31832 17316 31844
rect 17368 31832 17374 31884
rect 18141 31875 18199 31881
rect 17788 31844 18092 31872
rect 17037 31807 17095 31813
rect 17037 31773 17049 31807
rect 17083 31773 17095 31807
rect 17037 31767 17095 31773
rect 17129 31807 17187 31813
rect 17129 31773 17141 31807
rect 17175 31804 17187 31807
rect 17405 31807 17463 31813
rect 17175 31776 17356 31804
rect 17175 31773 17187 31776
rect 17129 31767 17187 31773
rect 1578 31736 1584 31748
rect 1539 31708 1584 31736
rect 1578 31696 1584 31708
rect 1636 31696 1642 31748
rect 17328 31736 17356 31776
rect 17405 31773 17417 31807
rect 17451 31804 17463 31807
rect 17494 31804 17500 31816
rect 17451 31776 17500 31804
rect 17451 31773 17463 31776
rect 17405 31767 17463 31773
rect 17494 31764 17500 31776
rect 17552 31764 17558 31816
rect 17788 31736 17816 31844
rect 17865 31807 17923 31813
rect 17865 31773 17877 31807
rect 17911 31804 17923 31807
rect 17954 31804 17960 31816
rect 17911 31776 17960 31804
rect 17911 31773 17923 31776
rect 17865 31767 17923 31773
rect 17954 31764 17960 31776
rect 18012 31764 18018 31816
rect 18064 31804 18092 31844
rect 18141 31841 18153 31875
rect 18187 31872 18199 31875
rect 18874 31872 18880 31884
rect 18187 31844 18880 31872
rect 18187 31841 18199 31844
rect 18141 31835 18199 31841
rect 18874 31832 18880 31844
rect 18932 31832 18938 31884
rect 18966 31832 18972 31884
rect 19024 31872 19030 31884
rect 19536 31881 19564 31980
rect 20990 31968 20996 31980
rect 21048 31968 21054 32020
rect 21174 31968 21180 32020
rect 21232 32008 21238 32020
rect 21232 31980 23152 32008
rect 21232 31968 21238 31980
rect 22925 31943 22983 31949
rect 22925 31940 22937 31943
rect 22204 31912 22937 31940
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 19024 31844 19441 31872
rect 19024 31832 19030 31844
rect 19429 31841 19441 31844
rect 19475 31841 19487 31875
rect 19429 31835 19487 31841
rect 19521 31875 19579 31881
rect 19521 31841 19533 31875
rect 19567 31841 19579 31875
rect 19521 31835 19579 31841
rect 19613 31875 19671 31881
rect 19613 31841 19625 31875
rect 19659 31872 19671 31875
rect 20162 31872 20168 31884
rect 19659 31844 20168 31872
rect 19659 31841 19671 31844
rect 19613 31835 19671 31841
rect 20162 31832 20168 31844
rect 20220 31832 20226 31884
rect 20533 31875 20591 31881
rect 20533 31872 20545 31875
rect 20456 31844 20545 31872
rect 18690 31804 18696 31816
rect 18064 31776 18696 31804
rect 18690 31764 18696 31776
rect 18748 31764 18754 31816
rect 19702 31804 19708 31816
rect 19663 31776 19708 31804
rect 19702 31764 19708 31776
rect 19760 31764 19766 31816
rect 20456 31736 20484 31844
rect 20533 31841 20545 31844
rect 20579 31841 20591 31875
rect 20533 31835 20591 31841
rect 20809 31875 20867 31881
rect 20809 31841 20821 31875
rect 20855 31872 20867 31875
rect 22204 31872 22232 31912
rect 22925 31909 22937 31912
rect 22971 31909 22983 31943
rect 23124 31940 23152 31980
rect 23198 31968 23204 32020
rect 23256 32008 23262 32020
rect 26510 32008 26516 32020
rect 23256 31980 26516 32008
rect 23256 31968 23262 31980
rect 26510 31968 26516 31980
rect 26568 31968 26574 32020
rect 26786 31968 26792 32020
rect 26844 32008 26850 32020
rect 30101 32011 30159 32017
rect 30101 32008 30113 32011
rect 26844 31980 30113 32008
rect 26844 31968 26850 31980
rect 30101 31977 30113 31980
rect 30147 32008 30159 32011
rect 30466 32008 30472 32020
rect 30147 31980 30472 32008
rect 30147 31977 30159 31980
rect 30101 31971 30159 31977
rect 30466 31968 30472 31980
rect 30524 31968 30530 32020
rect 27709 31943 27767 31949
rect 27709 31940 27721 31943
rect 23124 31912 27721 31940
rect 22925 31903 22983 31909
rect 27709 31909 27721 31912
rect 27755 31940 27767 31943
rect 27890 31940 27896 31952
rect 27755 31912 27896 31940
rect 27755 31909 27767 31912
rect 27709 31903 27767 31909
rect 27890 31900 27896 31912
rect 27948 31900 27954 31952
rect 28442 31940 28448 31952
rect 28403 31912 28448 31940
rect 28442 31900 28448 31912
rect 28500 31900 28506 31952
rect 31205 31943 31263 31949
rect 31205 31909 31217 31943
rect 31251 31940 31263 31943
rect 32306 31940 32312 31952
rect 31251 31912 32312 31940
rect 31251 31909 31263 31912
rect 31205 31903 31263 31909
rect 32306 31900 32312 31912
rect 32364 31900 32370 31952
rect 20855 31844 22232 31872
rect 20855 31841 20867 31844
rect 20809 31835 20867 31841
rect 22278 31832 22284 31884
rect 22336 31872 22342 31884
rect 22738 31872 22744 31884
rect 22336 31844 22381 31872
rect 22699 31844 22744 31872
rect 22336 31832 22342 31844
rect 22738 31832 22744 31844
rect 22796 31832 22802 31884
rect 30098 31832 30104 31884
rect 30156 31872 30162 31884
rect 47302 31872 47308 31884
rect 30156 31844 30972 31872
rect 47263 31844 47308 31872
rect 30156 31832 30162 31844
rect 23014 31804 23020 31816
rect 22940 31782 23020 31804
rect 22848 31776 23020 31782
rect 22848 31754 22968 31776
rect 23014 31764 23020 31776
rect 23072 31764 23078 31816
rect 23198 31764 23204 31816
rect 23256 31804 23262 31816
rect 25222 31804 25228 31816
rect 23256 31776 23301 31804
rect 25183 31776 25228 31804
rect 23256 31764 23262 31776
rect 25222 31764 25228 31776
rect 25280 31764 25286 31816
rect 26510 31764 26516 31816
rect 26568 31804 26574 31816
rect 28261 31807 28319 31813
rect 28261 31804 28273 31807
rect 26568 31776 28273 31804
rect 26568 31764 26574 31776
rect 28261 31773 28273 31776
rect 28307 31773 28319 31807
rect 30650 31804 30656 31816
rect 30611 31776 30656 31804
rect 28261 31767 28319 31773
rect 30650 31764 30656 31776
rect 30708 31764 30714 31816
rect 30944 31813 30972 31844
rect 47302 31832 47308 31844
rect 47360 31832 47366 31884
rect 30929 31807 30987 31813
rect 30929 31773 30941 31807
rect 30975 31773 30987 31807
rect 30929 31767 30987 31773
rect 31021 31807 31079 31813
rect 31021 31773 31033 31807
rect 31067 31804 31079 31807
rect 31110 31804 31116 31816
rect 31067 31776 31116 31804
rect 31067 31773 31079 31776
rect 31021 31767 31079 31773
rect 31110 31764 31116 31776
rect 31168 31764 31174 31816
rect 46566 31764 46572 31816
rect 46624 31804 46630 31816
rect 47581 31807 47639 31813
rect 47581 31804 47593 31807
rect 46624 31776 47593 31804
rect 46624 31764 46630 31776
rect 47581 31773 47593 31776
rect 47627 31773 47639 31807
rect 47581 31767 47639 31773
rect 20714 31736 20720 31748
rect 17328 31708 17816 31736
rect 19306 31708 20720 31736
rect 16850 31668 16856 31680
rect 16811 31640 16856 31668
rect 16850 31628 16856 31640
rect 16908 31628 16914 31680
rect 17954 31628 17960 31680
rect 18012 31668 18018 31680
rect 19306 31668 19334 31708
rect 20714 31696 20720 31708
rect 20772 31696 20778 31748
rect 22848 31736 22876 31754
rect 23106 31736 23112 31748
rect 22034 31708 22876 31736
rect 23067 31708 23112 31736
rect 23106 31696 23112 31708
rect 23164 31696 23170 31748
rect 25590 31696 25596 31748
rect 25648 31736 25654 31748
rect 26142 31736 26148 31748
rect 25648 31708 26148 31736
rect 25648 31696 25654 31708
rect 26142 31696 26148 31708
rect 26200 31696 26206 31748
rect 27522 31736 27528 31748
rect 27483 31708 27528 31736
rect 27522 31696 27528 31708
rect 27580 31696 27586 31748
rect 27632 31708 28994 31736
rect 18012 31640 19334 31668
rect 18012 31628 18018 31640
rect 20530 31628 20536 31680
rect 20588 31668 20594 31680
rect 27632 31668 27660 31708
rect 28966 31680 28994 31708
rect 29546 31696 29552 31748
rect 29604 31736 29610 31748
rect 30009 31739 30067 31745
rect 30009 31736 30021 31739
rect 29604 31708 30021 31736
rect 29604 31696 29610 31708
rect 30009 31705 30021 31708
rect 30055 31705 30067 31739
rect 30009 31699 30067 31705
rect 30558 31696 30564 31748
rect 30616 31736 30622 31748
rect 30837 31739 30895 31745
rect 30837 31736 30849 31739
rect 30616 31708 30849 31736
rect 30616 31696 30622 31708
rect 30837 31705 30849 31708
rect 30883 31736 30895 31739
rect 31202 31736 31208 31748
rect 30883 31708 31208 31736
rect 30883 31705 30895 31708
rect 30837 31699 30895 31705
rect 31202 31696 31208 31708
rect 31260 31696 31266 31748
rect 28966 31668 29000 31680
rect 20588 31640 27660 31668
rect 28907 31640 29000 31668
rect 20588 31628 20594 31640
rect 28994 31628 29000 31640
rect 29052 31668 29058 31680
rect 29454 31668 29460 31680
rect 29052 31640 29460 31668
rect 29052 31628 29058 31640
rect 29454 31628 29460 31640
rect 29512 31668 29518 31680
rect 30098 31668 30104 31680
rect 29512 31640 30104 31668
rect 29512 31628 29518 31640
rect 30098 31628 30104 31640
rect 30156 31628 30162 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1578 31424 1584 31476
rect 1636 31464 1642 31476
rect 2317 31467 2375 31473
rect 2317 31464 2329 31467
rect 1636 31436 2329 31464
rect 1636 31424 1642 31436
rect 2317 31433 2329 31436
rect 2363 31433 2375 31467
rect 2317 31427 2375 31433
rect 18417 31467 18475 31473
rect 18417 31433 18429 31467
rect 18463 31464 18475 31467
rect 18598 31464 18604 31476
rect 18463 31436 18604 31464
rect 18463 31433 18475 31436
rect 18417 31427 18475 31433
rect 18598 31424 18604 31436
rect 18656 31424 18662 31476
rect 18690 31424 18696 31476
rect 18748 31464 18754 31476
rect 18877 31467 18935 31473
rect 18877 31464 18889 31467
rect 18748 31436 18889 31464
rect 18748 31424 18754 31436
rect 18877 31433 18889 31436
rect 18923 31433 18935 31467
rect 23198 31464 23204 31476
rect 18877 31427 18935 31433
rect 22388 31436 23204 31464
rect 16850 31356 16856 31408
rect 16908 31396 16914 31408
rect 16945 31399 17003 31405
rect 16945 31396 16957 31399
rect 16908 31368 16957 31396
rect 16908 31356 16914 31368
rect 16945 31365 16957 31368
rect 16991 31365 17003 31399
rect 16945 31359 17003 31365
rect 2225 31331 2283 31337
rect 2225 31297 2237 31331
rect 2271 31328 2283 31331
rect 2314 31328 2320 31340
rect 2271 31300 2320 31328
rect 2271 31297 2283 31300
rect 2225 31291 2283 31297
rect 2314 31288 2320 31300
rect 2372 31288 2378 31340
rect 18046 31288 18052 31340
rect 18104 31288 18110 31340
rect 18616 31328 18644 31424
rect 20438 31356 20444 31408
rect 20496 31396 20502 31408
rect 22388 31405 22416 31436
rect 23198 31424 23204 31436
rect 23256 31424 23262 31476
rect 23569 31467 23627 31473
rect 23569 31433 23581 31467
rect 23615 31464 23627 31467
rect 23658 31464 23664 31476
rect 23615 31436 23664 31464
rect 23615 31433 23627 31436
rect 23569 31427 23627 31433
rect 23658 31424 23664 31436
rect 23716 31464 23722 31476
rect 24302 31464 24308 31476
rect 23716 31436 24308 31464
rect 23716 31424 23722 31436
rect 24302 31424 24308 31436
rect 24360 31424 24366 31476
rect 24762 31424 24768 31476
rect 24820 31464 24826 31476
rect 24820 31436 27292 31464
rect 24820 31424 24826 31436
rect 22373 31399 22431 31405
rect 20496 31368 22324 31396
rect 20496 31356 20502 31368
rect 19061 31331 19119 31337
rect 19061 31328 19073 31331
rect 18616 31300 19073 31328
rect 19061 31297 19073 31300
rect 19107 31297 19119 31331
rect 20990 31328 20996 31340
rect 20951 31300 20996 31328
rect 19061 31291 19119 31297
rect 20990 31288 20996 31300
rect 21048 31288 21054 31340
rect 22002 31288 22008 31340
rect 22060 31328 22066 31340
rect 22097 31331 22155 31337
rect 22097 31328 22109 31331
rect 22060 31300 22109 31328
rect 22060 31288 22066 31300
rect 22097 31297 22109 31300
rect 22143 31297 22155 31331
rect 22097 31291 22155 31297
rect 22190 31331 22248 31337
rect 22190 31297 22202 31331
rect 22236 31297 22248 31331
rect 22296 31328 22324 31368
rect 22373 31365 22385 31399
rect 22419 31365 22431 31399
rect 22373 31359 22431 31365
rect 22465 31399 22523 31405
rect 22465 31365 22477 31399
rect 22511 31396 22523 31399
rect 24854 31396 24860 31408
rect 22511 31368 24860 31396
rect 22511 31365 22523 31368
rect 22465 31359 22523 31365
rect 24854 31356 24860 31368
rect 24912 31356 24918 31408
rect 24946 31356 24952 31408
rect 25004 31396 25010 31408
rect 27264 31405 27292 31436
rect 27798 31424 27804 31476
rect 27856 31464 27862 31476
rect 27893 31467 27951 31473
rect 27893 31464 27905 31467
rect 27856 31436 27905 31464
rect 27856 31424 27862 31436
rect 27893 31433 27905 31436
rect 27939 31433 27951 31467
rect 27893 31427 27951 31433
rect 29454 31424 29460 31476
rect 29512 31464 29518 31476
rect 29549 31467 29607 31473
rect 29549 31464 29561 31467
rect 29512 31436 29561 31464
rect 29512 31424 29518 31436
rect 29549 31433 29561 31436
rect 29595 31433 29607 31467
rect 45094 31464 45100 31476
rect 29549 31427 29607 31433
rect 30300 31436 45100 31464
rect 27249 31399 27307 31405
rect 25004 31368 25912 31396
rect 25004 31356 25010 31368
rect 22562 31331 22620 31337
rect 22562 31328 22574 31331
rect 22296 31300 22574 31328
rect 22190 31291 22248 31297
rect 22562 31297 22574 31300
rect 22608 31297 22620 31331
rect 22562 31291 22620 31297
rect 16669 31263 16727 31269
rect 16669 31229 16681 31263
rect 16715 31260 16727 31263
rect 16715 31232 16804 31260
rect 16715 31229 16727 31232
rect 16669 31223 16727 31229
rect 16776 31124 16804 31232
rect 19334 31220 19340 31272
rect 19392 31260 19398 31272
rect 21269 31263 21327 31269
rect 19392 31232 19437 31260
rect 19392 31220 19398 31232
rect 21269 31229 21281 31263
rect 21315 31260 21327 31263
rect 22204 31260 22232 31291
rect 23106 31288 23112 31340
rect 23164 31328 23170 31340
rect 23385 31331 23443 31337
rect 23385 31328 23397 31331
rect 23164 31300 23397 31328
rect 23164 31288 23170 31300
rect 23385 31297 23397 31300
rect 23431 31297 23443 31331
rect 23385 31291 23443 31297
rect 22462 31260 22468 31272
rect 21315 31232 21404 31260
rect 21315 31229 21327 31232
rect 21269 31223 21327 31229
rect 19245 31195 19303 31201
rect 19245 31161 19257 31195
rect 19291 31192 19303 31195
rect 20806 31192 20812 31204
rect 19291 31164 20812 31192
rect 19291 31161 19303 31164
rect 19245 31155 19303 31161
rect 20806 31152 20812 31164
rect 20864 31152 20870 31204
rect 21082 31192 21088 31204
rect 21043 31164 21088 31192
rect 21082 31152 21088 31164
rect 21140 31152 21146 31204
rect 21376 31192 21404 31232
rect 21652 31232 22468 31260
rect 21652 31192 21680 31232
rect 22462 31220 22468 31232
rect 22520 31220 22526 31272
rect 21376 31164 21680 31192
rect 23400 31192 23428 31291
rect 23566 31288 23572 31340
rect 23624 31328 23630 31340
rect 23661 31331 23719 31337
rect 23661 31328 23673 31331
rect 23624 31300 23673 31328
rect 23624 31288 23630 31300
rect 23661 31297 23673 31300
rect 23707 31297 23719 31331
rect 23661 31291 23719 31297
rect 25406 31288 25412 31340
rect 25464 31328 25470 31340
rect 25884 31337 25912 31368
rect 27249 31365 27261 31399
rect 27295 31365 27307 31399
rect 27249 31359 27307 31365
rect 25501 31331 25559 31337
rect 25501 31328 25513 31331
rect 25464 31300 25513 31328
rect 25464 31288 25470 31300
rect 25501 31297 25513 31300
rect 25547 31328 25559 31331
rect 25869 31331 25927 31337
rect 25547 31300 25820 31328
rect 25547 31297 25559 31300
rect 25501 31291 25559 31297
rect 24762 31220 24768 31272
rect 24820 31260 24826 31272
rect 24946 31260 24952 31272
rect 24820 31232 24952 31260
rect 24820 31220 24826 31232
rect 24946 31220 24952 31232
rect 25004 31220 25010 31272
rect 25409 31195 25467 31201
rect 25409 31192 25421 31195
rect 23400 31164 25421 31192
rect 25409 31161 25421 31164
rect 25455 31192 25467 31195
rect 25498 31192 25504 31204
rect 25455 31164 25504 31192
rect 25455 31161 25467 31164
rect 25409 31155 25467 31161
rect 25498 31152 25504 31164
rect 25556 31152 25562 31204
rect 25792 31192 25820 31300
rect 25869 31297 25881 31331
rect 25915 31297 25927 31331
rect 26142 31328 26148 31340
rect 26103 31300 26148 31328
rect 25869 31291 25927 31297
rect 26142 31288 26148 31300
rect 26200 31288 26206 31340
rect 27982 31288 27988 31340
rect 28040 31328 28046 31340
rect 28077 31331 28135 31337
rect 28077 31328 28089 31331
rect 28040 31300 28089 31328
rect 28040 31288 28046 31300
rect 28077 31297 28089 31300
rect 28123 31297 28135 31331
rect 28077 31291 28135 31297
rect 28166 31288 28172 31340
rect 28224 31328 28230 31340
rect 28224 31300 28269 31328
rect 28224 31288 28230 31300
rect 28350 31288 28356 31340
rect 28408 31328 28414 31340
rect 28445 31331 28503 31337
rect 28445 31328 28457 31331
rect 28408 31300 28457 31328
rect 28408 31288 28414 31300
rect 28445 31297 28457 31300
rect 28491 31297 28503 31331
rect 28445 31291 28503 31297
rect 29365 31331 29423 31337
rect 29365 31297 29377 31331
rect 29411 31328 29423 31331
rect 29546 31328 29552 31340
rect 29411 31300 29552 31328
rect 29411 31297 29423 31300
rect 29365 31291 29423 31297
rect 27433 31263 27491 31269
rect 27433 31229 27445 31263
rect 27479 31260 27491 31263
rect 29380 31260 29408 31291
rect 29546 31288 29552 31300
rect 29604 31288 29610 31340
rect 30300 31337 30328 31436
rect 45094 31424 45100 31436
rect 45152 31424 45158 31476
rect 32122 31356 32128 31408
rect 32180 31396 32186 31408
rect 32493 31399 32551 31405
rect 32493 31396 32505 31399
rect 32180 31368 32505 31396
rect 32180 31356 32186 31368
rect 32493 31365 32505 31368
rect 32539 31365 32551 31399
rect 32493 31359 32551 31365
rect 30285 31331 30343 31337
rect 30285 31297 30297 31331
rect 30331 31297 30343 31331
rect 30285 31291 30343 31297
rect 30377 31331 30435 31337
rect 30377 31297 30389 31331
rect 30423 31297 30435 31331
rect 30558 31328 30564 31340
rect 30519 31300 30564 31328
rect 30377 31291 30435 31297
rect 27479 31232 29408 31260
rect 27479 31229 27491 31232
rect 27433 31223 27491 31229
rect 27448 31192 27476 31223
rect 30098 31220 30104 31272
rect 30156 31260 30162 31272
rect 30392 31260 30420 31291
rect 30558 31288 30564 31300
rect 30616 31288 30622 31340
rect 30653 31331 30711 31337
rect 30653 31297 30665 31331
rect 30699 31297 30711 31331
rect 32306 31328 32312 31340
rect 32267 31300 32312 31328
rect 30653 31291 30711 31297
rect 30156 31232 30420 31260
rect 30156 31220 30162 31232
rect 25792 31164 27476 31192
rect 29914 31152 29920 31204
rect 29972 31192 29978 31204
rect 30668 31192 30696 31291
rect 32306 31288 32312 31300
rect 32364 31288 32370 31340
rect 32582 31288 32588 31340
rect 32640 31328 32646 31340
rect 32640 31300 32685 31328
rect 32640 31288 32646 31300
rect 29972 31164 30696 31192
rect 29972 31152 29978 31164
rect 45554 31152 45560 31204
rect 45612 31192 45618 31204
rect 46014 31192 46020 31204
rect 45612 31164 46020 31192
rect 45612 31152 45618 31164
rect 46014 31152 46020 31164
rect 46072 31152 46078 31204
rect 17954 31124 17960 31136
rect 16776 31096 17960 31124
rect 17954 31084 17960 31096
rect 18012 31084 18018 31136
rect 21177 31127 21235 31133
rect 21177 31093 21189 31127
rect 21223 31124 21235 31127
rect 22002 31124 22008 31136
rect 21223 31096 22008 31124
rect 21223 31093 21235 31096
rect 21177 31087 21235 31093
rect 22002 31084 22008 31096
rect 22060 31084 22066 31136
rect 22646 31084 22652 31136
rect 22704 31124 22710 31136
rect 22741 31127 22799 31133
rect 22741 31124 22753 31127
rect 22704 31096 22753 31124
rect 22704 31084 22710 31096
rect 22741 31093 22753 31096
rect 22787 31093 22799 31127
rect 22741 31087 22799 31093
rect 28353 31127 28411 31133
rect 28353 31093 28365 31127
rect 28399 31124 28411 31127
rect 28626 31124 28632 31136
rect 28399 31096 28632 31124
rect 28399 31093 28411 31096
rect 28353 31087 28411 31093
rect 28626 31084 28632 31096
rect 28684 31084 28690 31136
rect 30006 31084 30012 31136
rect 30064 31124 30070 31136
rect 30101 31127 30159 31133
rect 30101 31124 30113 31127
rect 30064 31096 30113 31124
rect 30064 31084 30070 31096
rect 30101 31093 30113 31096
rect 30147 31093 30159 31127
rect 30101 31087 30159 31093
rect 32030 31084 32036 31136
rect 32088 31124 32094 31136
rect 32125 31127 32183 31133
rect 32125 31124 32137 31127
rect 32088 31096 32137 31124
rect 32088 31084 32094 31096
rect 32125 31093 32137 31096
rect 32171 31093 32183 31127
rect 32125 31087 32183 31093
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 22370 30880 22376 30932
rect 22428 30920 22434 30932
rect 22428 30892 23428 30920
rect 22428 30880 22434 30892
rect 23400 30852 23428 30892
rect 24854 30880 24860 30932
rect 24912 30920 24918 30932
rect 25501 30923 25559 30929
rect 25501 30920 25513 30923
rect 24912 30892 25513 30920
rect 24912 30880 24918 30892
rect 25501 30889 25513 30892
rect 25547 30889 25559 30923
rect 25501 30883 25559 30889
rect 26329 30923 26387 30929
rect 26329 30889 26341 30923
rect 26375 30920 26387 30923
rect 26970 30920 26976 30932
rect 26375 30892 26976 30920
rect 26375 30889 26387 30892
rect 26329 30883 26387 30889
rect 26970 30880 26976 30892
rect 27028 30880 27034 30932
rect 29270 30880 29276 30932
rect 29328 30920 29334 30932
rect 30193 30923 30251 30929
rect 30193 30920 30205 30923
rect 29328 30892 30205 30920
rect 29328 30880 29334 30892
rect 30193 30889 30205 30892
rect 30239 30889 30251 30923
rect 30193 30883 30251 30889
rect 31205 30923 31263 30929
rect 31205 30889 31217 30923
rect 31251 30920 31263 30923
rect 32582 30920 32588 30932
rect 31251 30892 32588 30920
rect 31251 30889 31263 30892
rect 31205 30883 31263 30889
rect 32582 30880 32588 30892
rect 32640 30880 32646 30932
rect 26513 30855 26571 30861
rect 26513 30852 26525 30855
rect 23400 30824 26525 30852
rect 26513 30821 26525 30824
rect 26559 30821 26571 30855
rect 26513 30815 26571 30821
rect 27985 30855 28043 30861
rect 27985 30821 27997 30855
rect 28031 30852 28043 30855
rect 28258 30852 28264 30864
rect 28031 30824 28264 30852
rect 28031 30821 28043 30824
rect 27985 30815 28043 30821
rect 28258 30812 28264 30824
rect 28316 30812 28322 30864
rect 29822 30812 29828 30864
rect 29880 30852 29886 30864
rect 29880 30824 30880 30852
rect 29880 30812 29886 30824
rect 8294 30744 8300 30796
rect 8352 30784 8358 30796
rect 14553 30787 14611 30793
rect 14553 30784 14565 30787
rect 8352 30756 14565 30784
rect 8352 30744 8358 30756
rect 14553 30753 14565 30756
rect 14599 30753 14611 30787
rect 14553 30747 14611 30753
rect 14642 30744 14648 30796
rect 14700 30784 14706 30796
rect 14700 30756 18092 30784
rect 14700 30744 14706 30756
rect 13998 30676 14004 30728
rect 14056 30716 14062 30728
rect 18064 30725 18092 30756
rect 23382 30744 23388 30796
rect 23440 30784 23446 30796
rect 28813 30787 28871 30793
rect 28813 30784 28825 30787
rect 23440 30756 26096 30784
rect 23440 30744 23446 30756
rect 14093 30719 14151 30725
rect 14093 30716 14105 30719
rect 14056 30688 14105 30716
rect 14056 30676 14062 30688
rect 14093 30685 14105 30688
rect 14139 30685 14151 30719
rect 14093 30679 14151 30685
rect 17681 30719 17739 30725
rect 17681 30685 17693 30719
rect 17727 30685 17739 30719
rect 17681 30679 17739 30685
rect 18049 30719 18107 30725
rect 18049 30685 18061 30719
rect 18095 30685 18107 30719
rect 18049 30679 18107 30685
rect 14274 30648 14280 30660
rect 14235 30620 14280 30648
rect 14274 30608 14280 30620
rect 14332 30608 14338 30660
rect 17696 30580 17724 30679
rect 20714 30676 20720 30728
rect 20772 30716 20778 30728
rect 21910 30716 21916 30728
rect 20772 30688 21916 30716
rect 20772 30676 20778 30688
rect 21910 30676 21916 30688
rect 21968 30716 21974 30728
rect 22086 30719 22144 30725
rect 22086 30716 22098 30719
rect 21968 30688 22098 30716
rect 21968 30676 21974 30688
rect 22086 30685 22098 30688
rect 22132 30685 22144 30719
rect 22086 30679 22144 30685
rect 23842 30676 23848 30728
rect 23900 30716 23906 30728
rect 24397 30719 24455 30725
rect 24397 30716 24409 30719
rect 23900 30688 24409 30716
rect 23900 30676 23906 30688
rect 24397 30685 24409 30688
rect 24443 30716 24455 30719
rect 24578 30716 24584 30728
rect 24443 30688 24584 30716
rect 24443 30685 24455 30688
rect 24397 30679 24455 30685
rect 24578 30676 24584 30688
rect 24636 30676 24642 30728
rect 25406 30716 25412 30728
rect 25367 30688 25412 30716
rect 25406 30676 25412 30688
rect 25464 30676 25470 30728
rect 26068 30725 26096 30756
rect 26804 30756 28825 30784
rect 26804 30728 26832 30756
rect 28813 30753 28825 30756
rect 28859 30784 28871 30787
rect 28997 30787 29055 30793
rect 28859 30756 28948 30784
rect 28859 30753 28871 30756
rect 28813 30747 28871 30753
rect 26053 30719 26111 30725
rect 26053 30685 26065 30719
rect 26099 30685 26111 30719
rect 26234 30716 26240 30728
rect 26195 30688 26240 30716
rect 26053 30679 26111 30685
rect 26234 30676 26240 30688
rect 26292 30676 26298 30728
rect 26329 30719 26387 30725
rect 26329 30685 26341 30719
rect 26375 30716 26387 30719
rect 26786 30716 26792 30728
rect 26375 30688 26792 30716
rect 26375 30685 26387 30688
rect 26329 30679 26387 30685
rect 26786 30676 26792 30688
rect 26844 30676 26850 30728
rect 28721 30719 28779 30725
rect 28721 30685 28733 30719
rect 28767 30685 28779 30719
rect 28920 30716 28948 30756
rect 28997 30753 29009 30787
rect 29043 30784 29055 30787
rect 29270 30784 29276 30796
rect 29043 30756 29276 30784
rect 29043 30753 29055 30756
rect 28997 30747 29055 30753
rect 29270 30744 29276 30756
rect 29328 30784 29334 30796
rect 30852 30793 30880 30824
rect 30837 30787 30895 30793
rect 29328 30756 30328 30784
rect 29328 30744 29334 30756
rect 30300 30728 30328 30756
rect 30837 30753 30849 30787
rect 30883 30753 30895 30787
rect 30837 30747 30895 30753
rect 31757 30787 31815 30793
rect 31757 30753 31769 30787
rect 31803 30753 31815 30787
rect 32030 30784 32036 30796
rect 31991 30756 32036 30784
rect 31757 30747 31815 30753
rect 29822 30716 29828 30728
rect 28920 30688 29828 30716
rect 28721 30679 28779 30685
rect 17862 30648 17868 30660
rect 17823 30620 17868 30648
rect 17862 30608 17868 30620
rect 17920 30608 17926 30660
rect 17957 30651 18015 30657
rect 17957 30617 17969 30651
rect 18003 30648 18015 30651
rect 18138 30648 18144 30660
rect 18003 30620 18144 30648
rect 18003 30617 18015 30620
rect 17957 30611 18015 30617
rect 18138 30608 18144 30620
rect 18196 30648 18202 30660
rect 20530 30648 20536 30660
rect 18196 30620 20536 30648
rect 18196 30608 18202 30620
rect 20530 30608 20536 30620
rect 20588 30608 20594 30660
rect 21266 30648 21272 30660
rect 21227 30620 21272 30648
rect 21266 30608 21272 30620
rect 21324 30608 21330 30660
rect 21453 30651 21511 30657
rect 21453 30617 21465 30651
rect 21499 30648 21511 30651
rect 22278 30648 22284 30660
rect 21499 30620 22284 30648
rect 21499 30617 21511 30620
rect 21453 30611 21511 30617
rect 22278 30608 22284 30620
rect 22336 30608 22342 30660
rect 22373 30651 22431 30657
rect 22373 30617 22385 30651
rect 22419 30648 22431 30651
rect 22646 30648 22652 30660
rect 22419 30620 22652 30648
rect 22419 30617 22431 30620
rect 22373 30611 22431 30617
rect 22646 30608 22652 30620
rect 22704 30608 22710 30660
rect 24489 30651 24547 30657
rect 24489 30648 24501 30651
rect 23598 30620 24501 30648
rect 24489 30617 24501 30620
rect 24535 30617 24547 30651
rect 24489 30611 24547 30617
rect 27154 30608 27160 30660
rect 27212 30648 27218 30660
rect 27522 30648 27528 30660
rect 27212 30620 27528 30648
rect 27212 30608 27218 30620
rect 27522 30608 27528 30620
rect 27580 30648 27586 30660
rect 27801 30651 27859 30657
rect 27801 30648 27813 30651
rect 27580 30620 27813 30648
rect 27580 30608 27586 30620
rect 27801 30617 27813 30620
rect 27847 30617 27859 30651
rect 28736 30648 28764 30679
rect 29822 30676 29828 30688
rect 29880 30676 29886 30728
rect 30006 30716 30012 30728
rect 29967 30688 30012 30716
rect 30006 30676 30012 30688
rect 30064 30676 30070 30728
rect 30282 30676 30288 30728
rect 30340 30716 30346 30728
rect 30340 30688 30385 30716
rect 30340 30676 30346 30688
rect 30650 30676 30656 30728
rect 30708 30716 30714 30728
rect 30926 30716 30932 30728
rect 30708 30688 30932 30716
rect 30708 30676 30714 30688
rect 30926 30676 30932 30688
rect 30984 30676 30990 30728
rect 29178 30648 29184 30660
rect 28736 30620 29184 30648
rect 27801 30611 27859 30617
rect 29178 30608 29184 30620
rect 29236 30608 29242 30660
rect 30466 30608 30472 30660
rect 30524 30648 30530 30660
rect 31772 30648 31800 30747
rect 32030 30744 32036 30756
rect 32088 30744 32094 30796
rect 30524 30620 31800 30648
rect 30524 30608 30530 30620
rect 32490 30608 32496 30660
rect 32548 30608 32554 30660
rect 18046 30580 18052 30592
rect 17696 30552 18052 30580
rect 18046 30540 18052 30552
rect 18104 30540 18110 30592
rect 18230 30580 18236 30592
rect 18191 30552 18236 30580
rect 18230 30540 18236 30552
rect 18288 30540 18294 30592
rect 21174 30540 21180 30592
rect 21232 30580 21238 30592
rect 21637 30583 21695 30589
rect 21637 30580 21649 30583
rect 21232 30552 21649 30580
rect 21232 30540 21238 30552
rect 21637 30549 21649 30552
rect 21683 30580 21695 30583
rect 23014 30580 23020 30592
rect 21683 30552 23020 30580
rect 21683 30549 21695 30552
rect 21637 30543 21695 30549
rect 23014 30540 23020 30552
rect 23072 30540 23078 30592
rect 23106 30540 23112 30592
rect 23164 30580 23170 30592
rect 23845 30583 23903 30589
rect 23845 30580 23857 30583
rect 23164 30552 23857 30580
rect 23164 30540 23170 30552
rect 23845 30549 23857 30552
rect 23891 30549 23903 30583
rect 28994 30580 29000 30592
rect 28955 30552 29000 30580
rect 23845 30543 23903 30549
rect 28994 30540 29000 30552
rect 29052 30540 29058 30592
rect 29825 30583 29883 30589
rect 29825 30549 29837 30583
rect 29871 30580 29883 30583
rect 30742 30580 30748 30592
rect 29871 30552 30748 30580
rect 29871 30549 29883 30552
rect 29825 30543 29883 30549
rect 30742 30540 30748 30552
rect 30800 30540 30806 30592
rect 30926 30540 30932 30592
rect 30984 30580 30990 30592
rect 33505 30583 33563 30589
rect 33505 30580 33517 30583
rect 30984 30552 33517 30580
rect 30984 30540 30990 30552
rect 33505 30549 33517 30552
rect 33551 30549 33563 30583
rect 33505 30543 33563 30549
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 17402 30336 17408 30388
rect 17460 30376 17466 30388
rect 17862 30376 17868 30388
rect 17460 30348 17868 30376
rect 17460 30336 17466 30348
rect 17862 30336 17868 30348
rect 17920 30376 17926 30388
rect 25685 30379 25743 30385
rect 25685 30376 25697 30379
rect 17920 30348 25697 30376
rect 17920 30336 17926 30348
rect 25685 30345 25697 30348
rect 25731 30376 25743 30379
rect 30558 30376 30564 30388
rect 25731 30348 30564 30376
rect 25731 30345 25743 30348
rect 25685 30339 25743 30345
rect 30558 30336 30564 30348
rect 30616 30336 30622 30388
rect 13725 30311 13783 30317
rect 13725 30277 13737 30311
rect 13771 30308 13783 30311
rect 14274 30308 14280 30320
rect 13771 30280 14280 30308
rect 13771 30277 13783 30280
rect 13725 30271 13783 30277
rect 14274 30268 14280 30280
rect 14332 30268 14338 30320
rect 16114 30308 16120 30320
rect 16075 30280 16120 30308
rect 16114 30268 16120 30280
rect 16172 30268 16178 30320
rect 22005 30311 22063 30317
rect 22005 30277 22017 30311
rect 22051 30308 22063 30311
rect 23290 30308 23296 30320
rect 22051 30280 23296 30308
rect 22051 30277 22063 30280
rect 22005 30271 22063 30277
rect 23290 30268 23296 30280
rect 23348 30268 23354 30320
rect 26234 30268 26240 30320
rect 26292 30308 26298 30320
rect 29549 30311 29607 30317
rect 29549 30308 29561 30311
rect 26292 30280 29561 30308
rect 26292 30268 26298 30280
rect 13630 30240 13636 30252
rect 13591 30212 13636 30240
rect 13630 30200 13636 30212
rect 13688 30200 13694 30252
rect 18230 30240 18236 30252
rect 18191 30212 18236 30240
rect 18230 30200 18236 30212
rect 18288 30200 18294 30252
rect 18417 30243 18475 30249
rect 18417 30209 18429 30243
rect 18463 30209 18475 30243
rect 18417 30203 18475 30209
rect 13906 30132 13912 30184
rect 13964 30172 13970 30184
rect 14277 30175 14335 30181
rect 14277 30172 14289 30175
rect 13964 30144 14289 30172
rect 13964 30132 13970 30144
rect 14277 30141 14289 30144
rect 14323 30141 14335 30175
rect 14277 30135 14335 30141
rect 14461 30175 14519 30181
rect 14461 30141 14473 30175
rect 14507 30172 14519 30175
rect 14642 30172 14648 30184
rect 14507 30144 14648 30172
rect 14507 30141 14519 30144
rect 14461 30135 14519 30141
rect 14642 30132 14648 30144
rect 14700 30132 14706 30184
rect 18432 30172 18460 30203
rect 18506 30200 18512 30252
rect 18564 30240 18570 30252
rect 18564 30212 18609 30240
rect 18564 30200 18570 30212
rect 21910 30200 21916 30252
rect 21968 30240 21974 30252
rect 22189 30243 22247 30249
rect 22189 30240 22201 30243
rect 21968 30212 22201 30240
rect 21968 30200 21974 30212
rect 22189 30209 22201 30212
rect 22235 30209 22247 30243
rect 22189 30203 22247 30209
rect 22462 30200 22468 30252
rect 22520 30240 22526 30252
rect 22649 30243 22707 30249
rect 22649 30240 22661 30243
rect 22520 30212 22661 30240
rect 22520 30200 22526 30212
rect 22649 30209 22661 30212
rect 22695 30209 22707 30243
rect 22830 30240 22836 30252
rect 22791 30212 22836 30240
rect 22649 30203 22707 30209
rect 22830 30200 22836 30212
rect 22888 30200 22894 30252
rect 23014 30200 23020 30252
rect 23072 30240 23078 30252
rect 23566 30240 23572 30252
rect 23072 30212 23572 30240
rect 23072 30200 23078 30212
rect 23566 30200 23572 30212
rect 23624 30200 23630 30252
rect 24578 30240 24584 30252
rect 24539 30212 24584 30240
rect 24578 30200 24584 30212
rect 24636 30200 24642 30252
rect 25498 30240 25504 30252
rect 25459 30212 25504 30240
rect 25498 30200 25504 30212
rect 25556 30240 25562 30252
rect 25774 30240 25780 30252
rect 25556 30212 25780 30240
rect 25556 30200 25562 30212
rect 25774 30200 25780 30212
rect 25832 30200 25838 30252
rect 26988 30249 27016 30280
rect 29549 30277 29561 30280
rect 29595 30277 29607 30311
rect 32122 30308 32128 30320
rect 29549 30271 29607 30277
rect 31726 30280 32128 30308
rect 26973 30243 27031 30249
rect 26973 30209 26985 30243
rect 27019 30209 27031 30243
rect 26973 30203 27031 30209
rect 27157 30243 27215 30249
rect 27157 30209 27169 30243
rect 27203 30240 27215 30243
rect 27430 30240 27436 30252
rect 27203 30212 27436 30240
rect 27203 30209 27215 30212
rect 27157 30203 27215 30209
rect 27430 30200 27436 30212
rect 27488 30200 27494 30252
rect 28353 30243 28411 30249
rect 28353 30209 28365 30243
rect 28399 30209 28411 30243
rect 28353 30203 28411 30209
rect 18432 30144 19334 30172
rect 19306 30104 19334 30144
rect 22370 30132 22376 30184
rect 22428 30172 22434 30184
rect 23106 30172 23112 30184
rect 22428 30144 23112 30172
rect 22428 30132 22434 30144
rect 23106 30132 23112 30144
rect 23164 30132 23170 30184
rect 28368 30172 28396 30203
rect 28442 30200 28448 30252
rect 28500 30240 28506 30252
rect 28537 30243 28595 30249
rect 28537 30240 28549 30243
rect 28500 30212 28549 30240
rect 28500 30200 28506 30212
rect 28537 30209 28549 30212
rect 28583 30209 28595 30243
rect 29178 30240 29184 30252
rect 29091 30212 29184 30240
rect 28537 30203 28595 30209
rect 29178 30200 29184 30212
rect 29236 30200 29242 30252
rect 29365 30243 29423 30249
rect 29365 30209 29377 30243
rect 29411 30240 29423 30243
rect 29730 30240 29736 30252
rect 29411 30212 29736 30240
rect 29411 30209 29423 30212
rect 29365 30203 29423 30209
rect 29730 30200 29736 30212
rect 29788 30200 29794 30252
rect 29822 30200 29828 30252
rect 29880 30240 29886 30252
rect 30009 30243 30067 30249
rect 30009 30240 30021 30243
rect 29880 30212 30021 30240
rect 29880 30200 29886 30212
rect 30009 30209 30021 30212
rect 30055 30209 30067 30243
rect 30009 30203 30067 30209
rect 30193 30243 30251 30249
rect 30193 30209 30205 30243
rect 30239 30240 30251 30243
rect 30282 30240 30288 30252
rect 30239 30212 30288 30240
rect 30239 30209 30251 30212
rect 30193 30203 30251 30209
rect 30282 30200 30288 30212
rect 30340 30240 30346 30252
rect 30558 30240 30564 30252
rect 30340 30212 30564 30240
rect 30340 30200 30346 30212
rect 30558 30200 30564 30212
rect 30616 30200 30622 30252
rect 28368 30144 28994 30172
rect 25682 30104 25688 30116
rect 19306 30076 25688 30104
rect 25682 30064 25688 30076
rect 25740 30064 25746 30116
rect 28721 30107 28779 30113
rect 28721 30104 28733 30107
rect 26988 30076 28733 30104
rect 26988 30048 27016 30076
rect 28721 30073 28733 30076
rect 28767 30073 28779 30107
rect 28721 30067 28779 30073
rect 18046 30036 18052 30048
rect 18007 30008 18052 30036
rect 18046 29996 18052 30008
rect 18104 29996 18110 30048
rect 21266 29996 21272 30048
rect 21324 30036 21330 30048
rect 22094 30036 22100 30048
rect 21324 30008 22100 30036
rect 21324 29996 21330 30008
rect 22094 29996 22100 30008
rect 22152 30036 22158 30048
rect 22646 30036 22652 30048
rect 22152 30008 22652 30036
rect 22152 29996 22158 30008
rect 22646 29996 22652 30008
rect 22704 29996 22710 30048
rect 24673 30039 24731 30045
rect 24673 30005 24685 30039
rect 24719 30036 24731 30039
rect 25130 30036 25136 30048
rect 24719 30008 25136 30036
rect 24719 30005 24731 30008
rect 24673 29999 24731 30005
rect 25130 29996 25136 30008
rect 25188 29996 25194 30048
rect 26970 30036 26976 30048
rect 26931 30008 26976 30036
rect 26970 29996 26976 30008
rect 27028 29996 27034 30048
rect 27062 29996 27068 30048
rect 27120 30036 27126 30048
rect 27341 30039 27399 30045
rect 27341 30036 27353 30039
rect 27120 30008 27353 30036
rect 27120 29996 27126 30008
rect 27341 30005 27353 30008
rect 27387 30005 27399 30039
rect 28966 30036 28994 30144
rect 29196 30104 29224 30200
rect 29638 30132 29644 30184
rect 29696 30172 29702 30184
rect 31726 30172 31754 30280
rect 32122 30268 32128 30280
rect 32180 30268 32186 30320
rect 32490 30308 32496 30320
rect 32451 30280 32496 30308
rect 32490 30268 32496 30280
rect 32548 30268 32554 30320
rect 32214 30200 32220 30252
rect 32272 30240 32278 30252
rect 32401 30243 32459 30249
rect 32401 30240 32413 30243
rect 32272 30212 32413 30240
rect 32272 30200 32278 30212
rect 32401 30209 32413 30212
rect 32447 30209 32459 30243
rect 32401 30203 32459 30209
rect 29696 30144 31754 30172
rect 29696 30132 29702 30144
rect 30650 30104 30656 30116
rect 29196 30076 30656 30104
rect 29270 30036 29276 30048
rect 28966 30008 29276 30036
rect 27341 29999 27399 30005
rect 29270 29996 29276 30008
rect 29328 29996 29334 30048
rect 30208 30045 30236 30076
rect 30650 30064 30656 30076
rect 30708 30064 30714 30116
rect 30193 30039 30251 30045
rect 30193 30005 30205 30039
rect 30239 30005 30251 30039
rect 30374 30036 30380 30048
rect 30335 30008 30380 30036
rect 30193 29999 30251 30005
rect 30374 29996 30380 30008
rect 30432 29996 30438 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 14642 29832 14648 29844
rect 14603 29804 14648 29832
rect 14642 29792 14648 29804
rect 14700 29792 14706 29844
rect 18417 29835 18475 29841
rect 18417 29801 18429 29835
rect 18463 29832 18475 29835
rect 18506 29832 18512 29844
rect 18463 29804 18512 29832
rect 18463 29801 18475 29804
rect 18417 29795 18475 29801
rect 18506 29792 18512 29804
rect 18564 29792 18570 29844
rect 22462 29832 22468 29844
rect 22423 29804 22468 29832
rect 22462 29792 22468 29804
rect 22520 29792 22526 29844
rect 26145 29835 26203 29841
rect 26145 29832 26157 29835
rect 23682 29804 26157 29832
rect 22649 29767 22707 29773
rect 22649 29733 22661 29767
rect 22695 29733 22707 29767
rect 22649 29727 22707 29733
rect 18233 29699 18291 29705
rect 18233 29665 18245 29699
rect 18279 29696 18291 29699
rect 20809 29699 20867 29705
rect 20809 29696 20821 29699
rect 18279 29668 20821 29696
rect 18279 29665 18291 29668
rect 18233 29659 18291 29665
rect 20809 29665 20821 29668
rect 20855 29696 20867 29699
rect 20855 29668 22094 29696
rect 20855 29665 20867 29668
rect 20809 29659 20867 29665
rect 22066 29640 22094 29668
rect 22186 29656 22192 29708
rect 22244 29696 22250 29708
rect 22244 29668 22508 29696
rect 22244 29656 22250 29668
rect 22480 29640 22508 29668
rect 13630 29588 13636 29640
rect 13688 29628 13694 29640
rect 14553 29631 14611 29637
rect 14553 29628 14565 29631
rect 13688 29600 14565 29628
rect 13688 29588 13694 29600
rect 14553 29597 14565 29600
rect 14599 29597 14611 29631
rect 18138 29628 18144 29640
rect 18099 29600 18144 29628
rect 14553 29591 14611 29597
rect 14568 29560 14596 29591
rect 18138 29588 18144 29600
rect 18196 29588 18202 29640
rect 20625 29631 20683 29637
rect 20625 29597 20637 29631
rect 20671 29628 20683 29631
rect 20714 29628 20720 29640
rect 20671 29600 20720 29628
rect 20671 29597 20683 29600
rect 20625 29591 20683 29597
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 20898 29628 20904 29640
rect 20859 29600 20904 29628
rect 20898 29588 20904 29600
rect 20956 29588 20962 29640
rect 22066 29600 22100 29640
rect 22094 29588 22100 29600
rect 22152 29628 22158 29640
rect 22462 29628 22468 29640
rect 22152 29600 22197 29628
rect 22423 29600 22468 29628
rect 22152 29588 22158 29600
rect 22462 29588 22468 29600
rect 22520 29588 22526 29640
rect 22664 29628 22692 29727
rect 22830 29656 22836 29708
rect 22888 29696 22894 29708
rect 23385 29699 23443 29705
rect 23385 29696 23397 29699
rect 22888 29668 23397 29696
rect 22888 29656 22894 29668
rect 23385 29665 23397 29668
rect 23431 29696 23443 29699
rect 23682 29696 23710 29804
rect 26145 29801 26157 29804
rect 26191 29801 26203 29835
rect 26145 29795 26203 29801
rect 26789 29835 26847 29841
rect 26789 29801 26801 29835
rect 26835 29832 26847 29835
rect 27246 29832 27252 29844
rect 26835 29804 27252 29832
rect 26835 29801 26847 29804
rect 26789 29795 26847 29801
rect 27246 29792 27252 29804
rect 27304 29832 27310 29844
rect 28442 29832 28448 29844
rect 27304 29804 28448 29832
rect 27304 29792 27310 29804
rect 28442 29792 28448 29804
rect 28500 29792 28506 29844
rect 29549 29835 29607 29841
rect 29549 29801 29561 29835
rect 29595 29832 29607 29835
rect 29914 29832 29920 29844
rect 29595 29804 29920 29832
rect 29595 29801 29607 29804
rect 29549 29795 29607 29801
rect 29914 29792 29920 29804
rect 29972 29792 29978 29844
rect 30558 29792 30564 29844
rect 30616 29832 30622 29844
rect 32217 29835 32275 29841
rect 32217 29832 32229 29835
rect 30616 29804 32229 29832
rect 30616 29792 30622 29804
rect 32217 29801 32229 29804
rect 32263 29801 32275 29835
rect 32217 29795 32275 29801
rect 25682 29724 25688 29776
rect 25740 29764 25746 29776
rect 28074 29764 28080 29776
rect 25740 29736 28080 29764
rect 25740 29724 25746 29736
rect 28074 29724 28080 29736
rect 28132 29764 28138 29776
rect 29638 29764 29644 29776
rect 28132 29736 29644 29764
rect 28132 29724 28138 29736
rect 29638 29724 29644 29736
rect 29696 29724 29702 29776
rect 23431 29668 23710 29696
rect 24397 29699 24455 29705
rect 23431 29665 23443 29668
rect 23385 29659 23443 29665
rect 24397 29665 24409 29699
rect 24443 29696 24455 29699
rect 30466 29696 30472 29708
rect 24443 29668 30472 29696
rect 24443 29665 24455 29668
rect 24397 29659 24455 29665
rect 30466 29656 30472 29668
rect 30524 29656 30530 29708
rect 30742 29696 30748 29708
rect 30703 29668 30748 29696
rect 30742 29656 30748 29668
rect 30800 29656 30806 29708
rect 23109 29631 23167 29637
rect 23109 29628 23121 29631
rect 22664 29600 23121 29628
rect 23109 29597 23121 29600
rect 23155 29597 23167 29631
rect 23290 29628 23296 29640
rect 23251 29600 23296 29628
rect 23109 29591 23167 29597
rect 23290 29588 23296 29600
rect 23348 29588 23354 29640
rect 23477 29631 23535 29637
rect 23477 29597 23489 29631
rect 23523 29628 23535 29631
rect 23566 29628 23572 29640
rect 23523 29600 23572 29628
rect 23523 29597 23535 29600
rect 23477 29591 23535 29597
rect 23566 29588 23572 29600
rect 23624 29588 23630 29640
rect 23661 29631 23719 29637
rect 23661 29597 23673 29631
rect 23707 29628 23719 29631
rect 23934 29628 23940 29640
rect 23707 29600 23940 29628
rect 23707 29597 23719 29600
rect 23661 29591 23719 29597
rect 18322 29560 18328 29572
rect 14568 29532 18328 29560
rect 18322 29520 18328 29532
rect 18380 29520 18386 29572
rect 19978 29520 19984 29572
rect 20036 29560 20042 29572
rect 20036 29532 22140 29560
rect 20036 29520 20042 29532
rect 20441 29495 20499 29501
rect 20441 29461 20453 29495
rect 20487 29492 20499 29495
rect 21542 29492 21548 29504
rect 20487 29464 21548 29492
rect 20487 29461 20499 29464
rect 20441 29455 20499 29461
rect 21542 29452 21548 29464
rect 21600 29452 21606 29504
rect 22112 29492 22140 29532
rect 22186 29520 22192 29572
rect 22244 29560 22250 29572
rect 23676 29560 23704 29591
rect 23934 29588 23940 29600
rect 23992 29588 23998 29640
rect 26697 29631 26755 29637
rect 26697 29597 26709 29631
rect 26743 29628 26755 29631
rect 27062 29628 27068 29640
rect 26743 29600 27068 29628
rect 26743 29597 26755 29600
rect 26697 29591 26755 29597
rect 27062 29588 27068 29600
rect 27120 29588 27126 29640
rect 27617 29631 27675 29637
rect 27617 29597 27629 29631
rect 27663 29597 27675 29631
rect 27617 29591 27675 29597
rect 27801 29631 27859 29637
rect 27801 29597 27813 29631
rect 27847 29628 27859 29631
rect 28166 29628 28172 29640
rect 27847 29600 28172 29628
rect 27847 29597 27859 29600
rect 27801 29591 27859 29597
rect 22244 29532 23704 29560
rect 23845 29563 23903 29569
rect 22244 29520 22250 29532
rect 23845 29529 23857 29563
rect 23891 29560 23903 29563
rect 24673 29563 24731 29569
rect 24673 29560 24685 29563
rect 23891 29532 24685 29560
rect 23891 29529 23903 29532
rect 23845 29523 23903 29529
rect 24673 29529 24685 29532
rect 24719 29529 24731 29563
rect 24673 29523 24731 29529
rect 25130 29520 25136 29572
rect 25188 29520 25194 29572
rect 27632 29560 27660 29591
rect 28166 29588 28172 29600
rect 28224 29628 28230 29640
rect 28261 29631 28319 29637
rect 28261 29628 28273 29631
rect 28224 29600 28273 29628
rect 28224 29588 28230 29600
rect 28261 29597 28273 29600
rect 28307 29628 28319 29631
rect 28350 29628 28356 29640
rect 28307 29600 28356 29628
rect 28307 29597 28319 29600
rect 28261 29591 28319 29597
rect 28350 29588 28356 29600
rect 28408 29588 28414 29640
rect 28445 29631 28503 29637
rect 28445 29597 28457 29631
rect 28491 29628 28503 29631
rect 28491 29600 28948 29628
rect 28491 29597 28503 29600
rect 28445 29591 28503 29597
rect 28460 29560 28488 29591
rect 27632 29532 28488 29560
rect 22922 29492 22928 29504
rect 22112 29464 22928 29492
rect 22922 29452 22928 29464
rect 22980 29492 22986 29504
rect 23290 29492 23296 29504
rect 22980 29464 23296 29492
rect 22980 29452 22986 29464
rect 23290 29452 23296 29464
rect 23348 29452 23354 29504
rect 27706 29492 27712 29504
rect 27667 29464 27712 29492
rect 27706 29452 27712 29464
rect 27764 29452 27770 29504
rect 27798 29452 27804 29504
rect 27856 29492 27862 29504
rect 28629 29495 28687 29501
rect 28629 29492 28641 29495
rect 27856 29464 28641 29492
rect 27856 29452 27862 29464
rect 28629 29461 28641 29464
rect 28675 29461 28687 29495
rect 28920 29492 28948 29600
rect 28994 29588 29000 29640
rect 29052 29628 29058 29640
rect 29825 29631 29883 29637
rect 29825 29628 29837 29631
rect 29052 29600 29837 29628
rect 29052 29588 29058 29600
rect 29825 29597 29837 29600
rect 29871 29597 29883 29631
rect 47302 29628 47308 29640
rect 47263 29600 47308 29628
rect 29825 29591 29883 29597
rect 47302 29588 47308 29600
rect 47360 29588 47366 29640
rect 47394 29588 47400 29640
rect 47452 29628 47458 29640
rect 47581 29631 47639 29637
rect 47581 29628 47593 29631
rect 47452 29600 47593 29628
rect 47452 29588 47458 29600
rect 47581 29597 47593 29600
rect 47627 29597 47639 29631
rect 47581 29591 47639 29597
rect 29546 29560 29552 29572
rect 29507 29532 29552 29560
rect 29546 29520 29552 29532
rect 29604 29520 29610 29572
rect 29733 29563 29791 29569
rect 29733 29529 29745 29563
rect 29779 29560 29791 29563
rect 30374 29560 30380 29572
rect 29779 29532 30380 29560
rect 29779 29529 29791 29532
rect 29733 29523 29791 29529
rect 29748 29492 29776 29523
rect 30374 29520 30380 29532
rect 30432 29520 30438 29572
rect 32122 29560 32128 29572
rect 31970 29532 32128 29560
rect 32122 29520 32128 29532
rect 32180 29520 32186 29572
rect 28920 29464 29776 29492
rect 28629 29455 28687 29461
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 20530 29288 20536 29300
rect 19306 29260 20536 29288
rect 7834 29180 7840 29232
rect 7892 29220 7898 29232
rect 19306 29220 19334 29260
rect 20530 29248 20536 29260
rect 20588 29248 20594 29300
rect 20714 29248 20720 29300
rect 20772 29248 20778 29300
rect 22094 29248 22100 29300
rect 22152 29288 22158 29300
rect 23477 29291 23535 29297
rect 23477 29288 23489 29291
rect 22152 29260 23489 29288
rect 22152 29248 22158 29260
rect 23477 29257 23489 29260
rect 23523 29257 23535 29291
rect 23477 29251 23535 29257
rect 24486 29248 24492 29300
rect 24544 29288 24550 29300
rect 24581 29291 24639 29297
rect 24581 29288 24593 29291
rect 24544 29260 24593 29288
rect 24544 29248 24550 29260
rect 24581 29257 24593 29260
rect 24627 29257 24639 29291
rect 30469 29291 30527 29297
rect 30469 29288 30481 29291
rect 24581 29251 24639 29257
rect 27908 29260 28304 29288
rect 20732 29220 20760 29248
rect 22186 29220 22192 29232
rect 7892 29192 19334 29220
rect 20456 29192 20760 29220
rect 21836 29192 22192 29220
rect 7892 29180 7898 29192
rect 10870 29112 10876 29164
rect 10928 29152 10934 29164
rect 13081 29155 13139 29161
rect 13081 29152 13093 29155
rect 10928 29124 13093 29152
rect 10928 29112 10934 29124
rect 13081 29121 13093 29124
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 13538 29112 13544 29164
rect 13596 29152 13602 29164
rect 13725 29155 13783 29161
rect 13725 29152 13737 29155
rect 13596 29124 13737 29152
rect 13596 29112 13602 29124
rect 13725 29121 13737 29124
rect 13771 29121 13783 29155
rect 13906 29152 13912 29164
rect 13867 29124 13912 29152
rect 13725 29115 13783 29121
rect 13906 29112 13912 29124
rect 13964 29112 13970 29164
rect 20162 29112 20168 29164
rect 20220 29150 20226 29164
rect 20456 29161 20484 29192
rect 20337 29153 20395 29159
rect 20220 29122 20263 29150
rect 20220 29112 20226 29122
rect 20337 29119 20349 29153
rect 20383 29119 20395 29153
rect 20337 29113 20395 29119
rect 20441 29155 20499 29161
rect 20441 29121 20453 29155
rect 20487 29121 20499 29155
rect 20441 29115 20499 29121
rect 20717 29155 20775 29161
rect 20717 29121 20729 29155
rect 20763 29152 20775 29155
rect 21836 29152 21864 29192
rect 22186 29180 22192 29192
rect 22244 29180 22250 29232
rect 22830 29220 22836 29232
rect 22480 29192 22836 29220
rect 22278 29152 22284 29164
rect 20763 29124 21864 29152
rect 22239 29124 22284 29152
rect 20763 29121 20775 29124
rect 20717 29115 20775 29121
rect 15838 29044 15844 29096
rect 15896 29084 15902 29096
rect 16669 29087 16727 29093
rect 16669 29084 16681 29087
rect 15896 29056 16681 29084
rect 15896 29044 15902 29056
rect 16669 29053 16681 29056
rect 16715 29053 16727 29087
rect 16850 29084 16856 29096
rect 16811 29056 16856 29084
rect 16669 29047 16727 29053
rect 16850 29044 16856 29056
rect 16908 29044 16914 29096
rect 17129 29087 17187 29093
rect 17129 29053 17141 29087
rect 17175 29053 17187 29087
rect 17129 29047 17187 29053
rect 13173 29019 13231 29025
rect 13173 28985 13185 29019
rect 13219 29016 13231 29019
rect 14090 29016 14096 29028
rect 13219 28988 14096 29016
rect 13219 28985 13231 28988
rect 13173 28979 13231 28985
rect 14090 28976 14096 28988
rect 14148 28976 14154 29028
rect 16574 28976 16580 29028
rect 16632 29016 16638 29028
rect 17144 29016 17172 29047
rect 19978 29044 19984 29096
rect 20036 29084 20042 29096
rect 20364 29084 20392 29113
rect 22278 29112 22284 29124
rect 22336 29112 22342 29164
rect 22480 29161 22508 29192
rect 22830 29180 22836 29192
rect 22888 29180 22894 29232
rect 22465 29155 22523 29161
rect 22465 29121 22477 29155
rect 22511 29121 22523 29155
rect 23109 29155 23167 29161
rect 23109 29152 23121 29155
rect 22465 29115 22523 29121
rect 22664 29124 23121 29152
rect 20036 29056 20392 29084
rect 20036 29044 20042 29056
rect 20530 29044 20536 29096
rect 20588 29084 20594 29096
rect 20588 29056 20633 29084
rect 20588 29044 20594 29056
rect 16632 28988 17172 29016
rect 16632 28976 16638 28988
rect 20162 28976 20168 29028
rect 20220 29016 20226 29028
rect 22002 29016 22008 29028
rect 20220 28988 22008 29016
rect 20220 28976 20226 28988
rect 22002 28976 22008 28988
rect 22060 28976 22066 29028
rect 22094 28976 22100 29028
rect 22152 29016 22158 29028
rect 22462 29016 22468 29028
rect 22152 28988 22468 29016
rect 22152 28976 22158 28988
rect 22462 28976 22468 28988
rect 22520 28976 22526 29028
rect 13814 28948 13820 28960
rect 13775 28920 13820 28948
rect 13814 28908 13820 28920
rect 13872 28908 13878 28960
rect 20898 28948 20904 28960
rect 20859 28920 20904 28948
rect 20898 28908 20904 28920
rect 20956 28908 20962 28960
rect 22278 28948 22284 28960
rect 22239 28920 22284 28948
rect 22278 28908 22284 28920
rect 22336 28908 22342 28960
rect 22370 28908 22376 28960
rect 22428 28948 22434 28960
rect 22664 28957 22692 29124
rect 23109 29121 23121 29124
rect 23155 29121 23167 29155
rect 23290 29152 23296 29164
rect 23251 29124 23296 29152
rect 23109 29115 23167 29121
rect 23290 29112 23296 29124
rect 23348 29112 23354 29164
rect 24489 29155 24547 29161
rect 24489 29121 24501 29155
rect 24535 29152 24547 29155
rect 24946 29152 24952 29164
rect 24535 29124 24952 29152
rect 24535 29121 24547 29124
rect 24489 29115 24547 29121
rect 24946 29112 24952 29124
rect 25004 29112 25010 29164
rect 25777 29155 25835 29161
rect 25777 29121 25789 29155
rect 25823 29121 25835 29155
rect 25777 29115 25835 29121
rect 27065 29155 27123 29161
rect 27065 29121 27077 29155
rect 27111 29152 27123 29155
rect 27798 29152 27804 29164
rect 27111 29124 27804 29152
rect 27111 29121 27123 29124
rect 27065 29115 27123 29121
rect 25792 29084 25820 29115
rect 27798 29112 27804 29124
rect 27856 29112 27862 29164
rect 27908 29161 27936 29260
rect 28276 29220 28304 29260
rect 28644 29260 30481 29288
rect 28644 29220 28672 29260
rect 30469 29257 30481 29260
rect 30515 29257 30527 29291
rect 30469 29251 30527 29257
rect 32122 29248 32128 29300
rect 32180 29288 32186 29300
rect 32217 29291 32275 29297
rect 32217 29288 32229 29291
rect 32180 29260 32229 29288
rect 32180 29248 32186 29260
rect 32217 29257 32229 29260
rect 32263 29257 32275 29291
rect 32217 29251 32275 29257
rect 28276 29192 28672 29220
rect 28718 29180 28724 29232
rect 28776 29220 28782 29232
rect 38286 29220 38292 29232
rect 28776 29192 29408 29220
rect 28776 29180 28782 29192
rect 27893 29155 27951 29161
rect 27893 29121 27905 29155
rect 27939 29121 27951 29155
rect 27893 29115 27951 29121
rect 28074 29112 28080 29164
rect 28132 29152 28138 29164
rect 28169 29155 28227 29161
rect 28169 29152 28181 29155
rect 28132 29124 28181 29152
rect 28132 29112 28138 29124
rect 28169 29121 28181 29124
rect 28215 29121 28227 29155
rect 28169 29115 28227 29121
rect 28261 29155 28319 29161
rect 28261 29121 28273 29155
rect 28307 29154 28319 29155
rect 28307 29152 28396 29154
rect 28442 29152 28448 29164
rect 28307 29126 28448 29152
rect 28307 29121 28319 29126
rect 28368 29124 28448 29126
rect 28261 29115 28319 29121
rect 28442 29112 28448 29124
rect 28500 29112 28506 29164
rect 29380 29161 29408 29192
rect 29564 29192 38292 29220
rect 29564 29161 29592 29192
rect 38286 29180 38292 29192
rect 38344 29180 38350 29232
rect 29181 29155 29239 29161
rect 29181 29152 29193 29155
rect 28966 29124 29193 29152
rect 27154 29084 27160 29096
rect 25792 29056 27160 29084
rect 27154 29044 27160 29056
rect 27212 29044 27218 29096
rect 27706 29044 27712 29096
rect 27764 29084 27770 29096
rect 27985 29087 28043 29093
rect 27985 29084 27997 29087
rect 27764 29056 27997 29084
rect 27764 29044 27770 29056
rect 27985 29053 27997 29056
rect 28031 29053 28043 29087
rect 28966 29084 28994 29124
rect 29181 29121 29193 29124
rect 29227 29121 29239 29155
rect 29181 29115 29239 29121
rect 29365 29155 29423 29161
rect 29365 29121 29377 29155
rect 29411 29121 29423 29155
rect 29365 29115 29423 29121
rect 29549 29155 29607 29161
rect 29549 29121 29561 29155
rect 29595 29121 29607 29155
rect 29549 29115 29607 29121
rect 29733 29155 29791 29161
rect 29733 29121 29745 29155
rect 29779 29121 29791 29155
rect 29733 29115 29791 29121
rect 27985 29047 28043 29053
rect 28184 29056 28994 29084
rect 29457 29087 29515 29093
rect 25958 29016 25964 29028
rect 25919 28988 25964 29016
rect 25958 28976 25964 28988
rect 26016 28976 26022 29028
rect 27433 29019 27491 29025
rect 27433 28985 27445 29019
rect 27479 29016 27491 29019
rect 27890 29016 27896 29028
rect 27479 28988 27896 29016
rect 27479 28985 27491 28988
rect 27433 28979 27491 28985
rect 27890 28976 27896 28988
rect 27948 28976 27954 29028
rect 28077 29019 28135 29025
rect 28077 28985 28089 29019
rect 28123 29016 28135 29019
rect 28184 29016 28212 29056
rect 29457 29053 29469 29087
rect 29503 29084 29515 29087
rect 29638 29084 29644 29096
rect 29503 29056 29644 29084
rect 29503 29053 29515 29056
rect 29457 29047 29515 29053
rect 29638 29044 29644 29056
rect 29696 29044 29702 29096
rect 28123 28988 28212 29016
rect 28123 28985 28135 28988
rect 28077 28979 28135 28985
rect 28258 28976 28264 29028
rect 28316 29016 28322 29028
rect 29759 29016 29787 29115
rect 29822 29112 29828 29164
rect 29880 29152 29886 29164
rect 30374 29152 30380 29164
rect 29880 29124 30380 29152
rect 29880 29112 29886 29124
rect 30374 29112 30380 29124
rect 30432 29112 30438 29164
rect 32122 29152 32128 29164
rect 32083 29124 32128 29152
rect 32122 29112 32128 29124
rect 32180 29112 32186 29164
rect 28316 28988 29787 29016
rect 29917 29019 29975 29025
rect 28316 28976 28322 28988
rect 29917 28985 29929 29019
rect 29963 29016 29975 29019
rect 30834 29016 30840 29028
rect 29963 28988 30840 29016
rect 29963 28985 29975 28988
rect 29917 28979 29975 28985
rect 30834 28976 30840 28988
rect 30892 28976 30898 29028
rect 22649 28951 22707 28957
rect 22649 28948 22661 28951
rect 22428 28920 22661 28948
rect 22428 28908 22434 28920
rect 22649 28917 22661 28920
rect 22695 28917 22707 28951
rect 22649 28911 22707 28917
rect 27249 28951 27307 28957
rect 27249 28917 27261 28951
rect 27295 28948 27307 28951
rect 27706 28948 27712 28960
rect 27295 28920 27712 28948
rect 27295 28917 27307 28920
rect 27249 28911 27307 28917
rect 27706 28908 27712 28920
rect 27764 28908 27770 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 15838 28744 15844 28756
rect 15799 28716 15844 28744
rect 15838 28704 15844 28716
rect 15896 28704 15902 28756
rect 18230 28704 18236 28756
rect 18288 28744 18294 28756
rect 18693 28747 18751 28753
rect 18693 28744 18705 28747
rect 18288 28716 18705 28744
rect 18288 28704 18294 28716
rect 18693 28713 18705 28716
rect 18739 28744 18751 28747
rect 18739 28716 20668 28744
rect 18739 28713 18751 28716
rect 18693 28707 18751 28713
rect 20640 28676 20668 28716
rect 20714 28704 20720 28756
rect 20772 28744 20778 28756
rect 20993 28747 21051 28753
rect 20993 28744 21005 28747
rect 20772 28716 21005 28744
rect 20772 28704 20778 28716
rect 20993 28713 21005 28716
rect 21039 28713 21051 28747
rect 21542 28744 21548 28756
rect 21503 28716 21548 28744
rect 20993 28707 21051 28713
rect 21542 28704 21548 28716
rect 21600 28704 21606 28756
rect 22002 28744 22008 28756
rect 21963 28716 22008 28744
rect 22002 28704 22008 28716
rect 22060 28704 22066 28756
rect 22370 28704 22376 28756
rect 22428 28744 22434 28756
rect 22465 28747 22523 28753
rect 22465 28744 22477 28747
rect 22428 28716 22477 28744
rect 22428 28704 22434 28716
rect 22465 28713 22477 28716
rect 22511 28713 22523 28747
rect 22465 28707 22523 28713
rect 26786 28704 26792 28756
rect 26844 28744 26850 28756
rect 26881 28747 26939 28753
rect 26881 28744 26893 28747
rect 26844 28716 26893 28744
rect 26844 28704 26850 28716
rect 26881 28713 26893 28716
rect 26927 28713 26939 28747
rect 28718 28744 28724 28756
rect 26881 28707 26939 28713
rect 28000 28716 28724 28744
rect 20806 28676 20812 28688
rect 20640 28648 20812 28676
rect 20806 28636 20812 28648
rect 20864 28636 20870 28688
rect 3694 28568 3700 28620
rect 3752 28608 3758 28620
rect 9769 28611 9827 28617
rect 9769 28608 9781 28611
rect 3752 28580 9781 28608
rect 3752 28568 3758 28580
rect 9769 28577 9781 28580
rect 9815 28577 9827 28611
rect 9769 28571 9827 28577
rect 13265 28611 13323 28617
rect 13265 28577 13277 28611
rect 13311 28608 13323 28611
rect 13814 28608 13820 28620
rect 13311 28580 13820 28608
rect 13311 28577 13323 28580
rect 13265 28571 13323 28577
rect 13814 28568 13820 28580
rect 13872 28568 13878 28620
rect 14090 28608 14096 28620
rect 14051 28580 14096 28608
rect 14090 28568 14096 28580
rect 14148 28568 14154 28620
rect 16945 28611 17003 28617
rect 16945 28577 16957 28611
rect 16991 28608 17003 28611
rect 17954 28608 17960 28620
rect 16991 28580 17960 28608
rect 16991 28577 17003 28580
rect 16945 28571 17003 28577
rect 17954 28568 17960 28580
rect 18012 28608 18018 28620
rect 19521 28611 19579 28617
rect 18012 28580 19288 28608
rect 18012 28568 18018 28580
rect 19260 28552 19288 28580
rect 19521 28577 19533 28611
rect 19567 28608 19579 28611
rect 20898 28608 20904 28620
rect 19567 28580 20904 28608
rect 19567 28577 19579 28580
rect 19521 28571 19579 28577
rect 20898 28568 20904 28580
rect 20956 28568 20962 28620
rect 21729 28611 21787 28617
rect 21729 28577 21741 28611
rect 21775 28608 21787 28611
rect 22094 28608 22100 28620
rect 21775 28580 22100 28608
rect 21775 28577 21787 28580
rect 21729 28571 21787 28577
rect 22094 28568 22100 28580
rect 22152 28608 22158 28620
rect 25958 28608 25964 28620
rect 22152 28580 25964 28608
rect 22152 28568 22158 28580
rect 25958 28568 25964 28580
rect 26016 28568 26022 28620
rect 28000 28608 28028 28716
rect 28718 28704 28724 28716
rect 28776 28704 28782 28756
rect 30374 28704 30380 28756
rect 30432 28744 30438 28756
rect 32309 28747 32367 28753
rect 32309 28744 32321 28747
rect 30432 28716 32321 28744
rect 30432 28704 30438 28716
rect 32309 28713 32321 28716
rect 32355 28713 32367 28747
rect 32309 28707 32367 28713
rect 28074 28636 28080 28688
rect 28132 28676 28138 28688
rect 28132 28648 28304 28676
rect 28132 28636 28138 28648
rect 28276 28617 28304 28648
rect 28261 28611 28319 28617
rect 28000 28580 28120 28608
rect 9309 28543 9367 28549
rect 9309 28509 9321 28543
rect 9355 28509 9367 28543
rect 12066 28540 12072 28552
rect 12027 28512 12072 28540
rect 9309 28503 9367 28509
rect 9324 28404 9352 28503
rect 12066 28500 12072 28512
rect 12124 28500 12130 28552
rect 12253 28543 12311 28549
rect 12253 28509 12265 28543
rect 12299 28540 12311 28543
rect 13078 28540 13084 28552
rect 12299 28512 13084 28540
rect 12299 28509 12311 28512
rect 12253 28503 12311 28509
rect 13078 28500 13084 28512
rect 13136 28500 13142 28552
rect 13170 28500 13176 28552
rect 13228 28540 13234 28552
rect 19242 28540 19248 28552
rect 13228 28512 13273 28540
rect 19203 28512 19248 28540
rect 13228 28500 13234 28512
rect 19242 28500 19248 28512
rect 19300 28500 19306 28552
rect 21453 28543 21511 28549
rect 21453 28509 21465 28543
rect 21499 28509 21511 28543
rect 21453 28503 21511 28509
rect 9493 28475 9551 28481
rect 9493 28441 9505 28475
rect 9539 28472 9551 28475
rect 10042 28472 10048 28484
rect 9539 28444 10048 28472
rect 9539 28441 9551 28444
rect 9493 28435 9551 28441
rect 10042 28432 10048 28444
rect 10100 28432 10106 28484
rect 14369 28475 14427 28481
rect 14369 28441 14381 28475
rect 14415 28441 14427 28475
rect 14369 28435 14427 28441
rect 9950 28404 9956 28416
rect 9324 28376 9956 28404
rect 9950 28364 9956 28376
rect 10008 28364 10014 28416
rect 11790 28364 11796 28416
rect 11848 28404 11854 28416
rect 12161 28407 12219 28413
rect 12161 28404 12173 28407
rect 11848 28376 12173 28404
rect 11848 28364 11854 28376
rect 12161 28373 12173 28376
rect 12207 28373 12219 28407
rect 12161 28367 12219 28373
rect 13541 28407 13599 28413
rect 13541 28373 13553 28407
rect 13587 28404 13599 28407
rect 14384 28404 14412 28435
rect 14826 28432 14832 28484
rect 14884 28432 14890 28484
rect 17221 28475 17279 28481
rect 17221 28441 17233 28475
rect 17267 28441 17279 28475
rect 18874 28472 18880 28484
rect 18446 28444 18880 28472
rect 17221 28435 17279 28441
rect 13587 28376 14412 28404
rect 17236 28404 17264 28435
rect 18874 28432 18880 28444
rect 18932 28432 18938 28484
rect 19978 28432 19984 28484
rect 20036 28432 20042 28484
rect 21468 28472 21496 28503
rect 22186 28500 22192 28552
rect 22244 28540 22250 28552
rect 22465 28543 22523 28549
rect 22465 28540 22477 28543
rect 22244 28512 22477 28540
rect 22244 28500 22250 28512
rect 22465 28509 22477 28512
rect 22511 28509 22523 28543
rect 22646 28540 22652 28552
rect 22607 28512 22652 28540
rect 22465 28503 22523 28509
rect 22646 28500 22652 28512
rect 22704 28540 22710 28552
rect 23290 28540 23296 28552
rect 22704 28512 23296 28540
rect 22704 28500 22710 28512
rect 23290 28500 23296 28512
rect 23348 28500 23354 28552
rect 27890 28540 27896 28552
rect 27851 28512 27896 28540
rect 27890 28500 27896 28512
rect 27948 28500 27954 28552
rect 28092 28549 28120 28580
rect 28261 28577 28273 28611
rect 28307 28577 28319 28611
rect 30834 28608 30840 28620
rect 30795 28580 30840 28608
rect 28261 28571 28319 28577
rect 30834 28568 30840 28580
rect 30892 28568 30898 28620
rect 46477 28611 46535 28617
rect 46477 28577 46489 28611
rect 46523 28608 46535 28611
rect 47394 28608 47400 28620
rect 46523 28580 47400 28608
rect 46523 28577 46535 28580
rect 46477 28571 46535 28577
rect 47394 28568 47400 28580
rect 47452 28568 47458 28620
rect 47670 28608 47676 28620
rect 47631 28580 47676 28608
rect 47670 28568 47676 28580
rect 47728 28568 47734 28620
rect 28077 28543 28135 28549
rect 28077 28509 28089 28543
rect 28123 28509 28135 28543
rect 28077 28503 28135 28509
rect 28166 28500 28172 28552
rect 28224 28540 28230 28552
rect 28224 28512 28269 28540
rect 28224 28500 28230 28512
rect 28350 28500 28356 28552
rect 28408 28540 28414 28552
rect 28445 28543 28503 28549
rect 28445 28540 28457 28543
rect 28408 28512 28457 28540
rect 28408 28500 28414 28512
rect 28445 28509 28457 28512
rect 28491 28509 28503 28543
rect 28445 28503 28503 28509
rect 28534 28500 28540 28552
rect 28592 28540 28598 28552
rect 29641 28543 29699 28549
rect 29641 28540 29653 28543
rect 28592 28512 29653 28540
rect 28592 28500 28598 28512
rect 29641 28509 29653 28512
rect 29687 28509 29699 28543
rect 29641 28503 29699 28509
rect 30561 28543 30619 28549
rect 30561 28509 30573 28543
rect 30607 28509 30619 28543
rect 30561 28503 30619 28509
rect 46293 28543 46351 28549
rect 46293 28509 46305 28543
rect 46339 28509 46351 28543
rect 46293 28503 46351 28509
rect 26789 28475 26847 28481
rect 21468 28444 22094 28472
rect 18046 28404 18052 28416
rect 17236 28376 18052 28404
rect 13587 28373 13599 28376
rect 13541 28367 13599 28373
rect 18046 28364 18052 28376
rect 18104 28364 18110 28416
rect 22066 28404 22094 28444
rect 26789 28441 26801 28475
rect 26835 28472 26847 28475
rect 27430 28472 27436 28484
rect 26835 28444 27436 28472
rect 26835 28441 26847 28444
rect 26789 28435 26847 28441
rect 27430 28432 27436 28444
rect 27488 28432 27494 28484
rect 29730 28472 29736 28484
rect 28460 28444 29736 28472
rect 28460 28416 28488 28444
rect 29730 28432 29736 28444
rect 29788 28472 29794 28484
rect 29825 28475 29883 28481
rect 29825 28472 29837 28475
rect 29788 28444 29837 28472
rect 29788 28432 29794 28444
rect 29825 28441 29837 28444
rect 29871 28472 29883 28475
rect 30466 28472 30472 28484
rect 29871 28444 30472 28472
rect 29871 28441 29883 28444
rect 29825 28435 29883 28441
rect 30466 28432 30472 28444
rect 30524 28472 30530 28484
rect 30576 28472 30604 28503
rect 32214 28472 32220 28484
rect 30524 28444 30604 28472
rect 32062 28444 32220 28472
rect 30524 28432 30530 28444
rect 32214 28432 32220 28444
rect 32272 28432 32278 28484
rect 46308 28472 46336 28503
rect 46566 28472 46572 28484
rect 46308 28444 46572 28472
rect 46566 28432 46572 28444
rect 46624 28432 46630 28484
rect 22462 28404 22468 28416
rect 22066 28376 22468 28404
rect 22462 28364 22468 28376
rect 22520 28404 22526 28416
rect 22833 28407 22891 28413
rect 22833 28404 22845 28407
rect 22520 28376 22845 28404
rect 22520 28364 22526 28376
rect 22833 28373 22845 28376
rect 22879 28373 22891 28407
rect 22833 28367 22891 28373
rect 28442 28364 28448 28416
rect 28500 28364 28506 28416
rect 28629 28407 28687 28413
rect 28629 28373 28641 28407
rect 28675 28404 28687 28407
rect 28718 28404 28724 28416
rect 28675 28376 28724 28404
rect 28675 28373 28687 28376
rect 28629 28367 28687 28373
rect 28718 28364 28724 28376
rect 28776 28364 28782 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 10042 28200 10048 28212
rect 10003 28172 10048 28200
rect 10042 28160 10048 28172
rect 10100 28160 10106 28212
rect 14737 28203 14795 28209
rect 14737 28169 14749 28203
rect 14783 28200 14795 28203
rect 14826 28200 14832 28212
rect 14783 28172 14832 28200
rect 14783 28169 14795 28172
rect 14737 28163 14795 28169
rect 14826 28160 14832 28172
rect 14884 28160 14890 28212
rect 16025 28203 16083 28209
rect 16025 28169 16037 28203
rect 16071 28200 16083 28203
rect 16850 28200 16856 28212
rect 16071 28172 16856 28200
rect 16071 28169 16083 28172
rect 16025 28163 16083 28169
rect 16850 28160 16856 28172
rect 16908 28160 16914 28212
rect 18874 28160 18880 28212
rect 18932 28200 18938 28212
rect 19061 28203 19119 28209
rect 19061 28200 19073 28203
rect 18932 28172 19073 28200
rect 18932 28160 18938 28172
rect 19061 28169 19073 28172
rect 19107 28169 19119 28203
rect 19978 28200 19984 28212
rect 19939 28172 19984 28200
rect 19061 28163 19119 28169
rect 19978 28160 19984 28172
rect 20036 28160 20042 28212
rect 22094 28160 22100 28212
rect 22152 28200 22158 28212
rect 22833 28203 22891 28209
rect 22833 28200 22845 28203
rect 22152 28172 22845 28200
rect 22152 28160 22158 28172
rect 22833 28169 22845 28172
rect 22879 28200 22891 28203
rect 23198 28200 23204 28212
rect 22879 28172 23204 28200
rect 22879 28169 22891 28172
rect 22833 28163 22891 28169
rect 23198 28160 23204 28172
rect 23256 28200 23262 28212
rect 24045 28203 24103 28209
rect 24045 28200 24057 28203
rect 23256 28172 24057 28200
rect 23256 28160 23262 28172
rect 24045 28169 24057 28172
rect 24091 28169 24103 28203
rect 24045 28163 24103 28169
rect 28166 28160 28172 28212
rect 28224 28200 28230 28212
rect 30193 28203 30251 28209
rect 30193 28200 30205 28203
rect 28224 28172 30205 28200
rect 28224 28160 28230 28172
rect 30193 28169 30205 28172
rect 30239 28169 30251 28203
rect 32214 28200 32220 28212
rect 32175 28172 32220 28200
rect 30193 28163 30251 28169
rect 32214 28160 32220 28172
rect 32272 28160 32278 28212
rect 47670 28200 47676 28212
rect 35866 28172 47676 28200
rect 11790 28132 11796 28144
rect 11751 28104 11796 28132
rect 11790 28092 11796 28104
rect 11848 28092 11854 28144
rect 13909 28135 13967 28141
rect 13909 28132 13921 28135
rect 13018 28104 13921 28132
rect 13909 28101 13921 28104
rect 13955 28101 13967 28135
rect 13909 28095 13967 28101
rect 20714 28092 20720 28144
rect 20772 28132 20778 28144
rect 20993 28135 21051 28141
rect 20993 28132 21005 28135
rect 20772 28104 21005 28132
rect 20772 28092 20778 28104
rect 20993 28101 21005 28104
rect 21039 28101 21051 28135
rect 20993 28095 21051 28101
rect 23750 28092 23756 28144
rect 23808 28132 23814 28144
rect 23845 28135 23903 28141
rect 23845 28132 23857 28135
rect 23808 28104 23857 28132
rect 23808 28092 23814 28104
rect 23845 28101 23857 28104
rect 23891 28101 23903 28135
rect 23845 28095 23903 28101
rect 25501 28135 25559 28141
rect 25501 28101 25513 28135
rect 25547 28132 25559 28135
rect 25590 28132 25596 28144
rect 25547 28104 25596 28132
rect 25547 28101 25559 28104
rect 25501 28095 25559 28101
rect 25590 28092 25596 28104
rect 25648 28092 25654 28144
rect 25866 28132 25872 28144
rect 25827 28104 25872 28132
rect 25866 28092 25872 28104
rect 25924 28092 25930 28144
rect 25958 28092 25964 28144
rect 26016 28132 26022 28144
rect 28718 28132 28724 28144
rect 26016 28104 27292 28132
rect 28679 28104 28724 28132
rect 26016 28092 26022 28104
rect 9953 28067 10011 28073
rect 9953 28033 9965 28067
rect 9999 28033 10011 28067
rect 10870 28064 10876 28076
rect 10831 28036 10876 28064
rect 9953 28027 10011 28033
rect 9968 27928 9996 28027
rect 10870 28024 10876 28036
rect 10928 28024 10934 28076
rect 13817 28067 13875 28073
rect 13817 28033 13829 28067
rect 13863 28064 13875 28067
rect 14090 28064 14096 28076
rect 13863 28036 14096 28064
rect 13863 28033 13875 28036
rect 13817 28027 13875 28033
rect 14090 28024 14096 28036
rect 14148 28064 14154 28076
rect 14645 28067 14703 28073
rect 14645 28064 14657 28067
rect 14148 28036 14657 28064
rect 14148 28024 14154 28036
rect 14645 28033 14657 28036
rect 14691 28033 14703 28067
rect 14645 28027 14703 28033
rect 15933 28067 15991 28073
rect 15933 28033 15945 28067
rect 15979 28064 15991 28067
rect 15979 28036 16013 28064
rect 15979 28033 15991 28036
rect 15933 28027 15991 28033
rect 10965 27999 11023 28005
rect 10965 27965 10977 27999
rect 11011 27996 11023 27999
rect 11517 27999 11575 28005
rect 11517 27996 11529 27999
rect 11011 27968 11529 27996
rect 11011 27965 11023 27968
rect 10965 27959 11023 27965
rect 11517 27965 11529 27968
rect 11563 27965 11575 27999
rect 15948 27996 15976 28027
rect 18598 28024 18604 28076
rect 18656 28064 18662 28076
rect 18969 28067 19027 28073
rect 18969 28064 18981 28067
rect 18656 28036 18981 28064
rect 18656 28024 18662 28036
rect 18969 28033 18981 28036
rect 19015 28064 19027 28067
rect 19889 28067 19947 28073
rect 19889 28064 19901 28067
rect 19015 28036 19901 28064
rect 19015 28033 19027 28036
rect 18969 28027 19027 28033
rect 19889 28033 19901 28036
rect 19935 28033 19947 28067
rect 20806 28064 20812 28076
rect 20767 28036 20812 28064
rect 19889 28027 19947 28033
rect 20806 28024 20812 28036
rect 20864 28024 20870 28076
rect 22646 28064 22652 28076
rect 22607 28036 22652 28064
rect 22646 28024 22652 28036
rect 22704 28024 22710 28076
rect 16022 27996 16028 28008
rect 11517 27959 11575 27965
rect 11624 27968 16028 27996
rect 11624 27928 11652 27968
rect 16022 27956 16028 27968
rect 16080 27956 16086 28008
rect 16666 27996 16672 28008
rect 16627 27968 16672 27996
rect 16666 27956 16672 27968
rect 16724 27956 16730 28008
rect 16850 27996 16856 28008
rect 16811 27968 16856 27996
rect 16850 27956 16856 27968
rect 16908 27956 16914 28008
rect 17129 27999 17187 28005
rect 17129 27965 17141 27999
rect 17175 27965 17187 27999
rect 17129 27959 17187 27965
rect 17144 27928 17172 27959
rect 21082 27956 21088 28008
rect 21140 27996 21146 28008
rect 25884 27996 25912 28092
rect 26786 28024 26792 28076
rect 26844 28064 26850 28076
rect 27264 28073 27292 28104
rect 28718 28092 28724 28104
rect 28776 28092 28782 28144
rect 30834 28132 30840 28144
rect 29946 28104 30840 28132
rect 30834 28092 30840 28104
rect 30892 28092 30898 28144
rect 26973 28067 27031 28073
rect 26973 28064 26985 28067
rect 26844 28036 26985 28064
rect 26844 28024 26850 28036
rect 26973 28033 26985 28036
rect 27019 28033 27031 28067
rect 26973 28027 27031 28033
rect 27249 28067 27307 28073
rect 27249 28033 27261 28067
rect 27295 28033 27307 28067
rect 27249 28027 27307 28033
rect 27338 28024 27344 28076
rect 27396 28064 27402 28076
rect 28442 28064 28448 28076
rect 27396 28036 28448 28064
rect 27396 28024 27402 28036
rect 28442 28024 28448 28036
rect 28500 28024 28506 28076
rect 30650 28024 30656 28076
rect 30708 28064 30714 28076
rect 32122 28064 32128 28076
rect 30708 28036 32128 28064
rect 30708 28024 30714 28036
rect 32122 28024 32128 28036
rect 32180 28024 32186 28076
rect 21140 27968 25912 27996
rect 21140 27956 21146 27968
rect 27890 27956 27896 28008
rect 27948 27996 27954 28008
rect 28810 27996 28816 28008
rect 27948 27968 28816 27996
rect 27948 27956 27954 27968
rect 28810 27956 28816 27968
rect 28868 27996 28874 28008
rect 35866 27996 35894 28172
rect 47670 28160 47676 28172
rect 47728 28160 47734 28212
rect 47118 28024 47124 28076
rect 47176 28064 47182 28076
rect 47578 28064 47584 28076
rect 47176 28036 47584 28064
rect 47176 28024 47182 28036
rect 47578 28024 47584 28036
rect 47636 28024 47642 28076
rect 28868 27968 35894 27996
rect 28868 27956 28874 27968
rect 24486 27928 24492 27940
rect 9968 27900 11652 27928
rect 13188 27900 17172 27928
rect 24044 27900 24492 27928
rect 3970 27820 3976 27872
rect 4028 27860 4034 27872
rect 13188 27860 13216 27900
rect 4028 27832 13216 27860
rect 4028 27820 4034 27832
rect 13262 27820 13268 27872
rect 13320 27860 13326 27872
rect 21177 27863 21235 27869
rect 13320 27832 13365 27860
rect 13320 27820 13326 27832
rect 21177 27829 21189 27863
rect 21223 27860 21235 27863
rect 22186 27860 22192 27872
rect 21223 27832 22192 27860
rect 21223 27829 21235 27832
rect 21177 27823 21235 27829
rect 22186 27820 22192 27832
rect 22244 27820 22250 27872
rect 24044 27869 24072 27900
rect 24486 27888 24492 27900
rect 24544 27888 24550 27940
rect 24029 27863 24087 27869
rect 24029 27829 24041 27863
rect 24075 27829 24087 27863
rect 24210 27860 24216 27872
rect 24171 27832 24216 27860
rect 24029 27823 24087 27829
rect 24210 27820 24216 27832
rect 24268 27820 24274 27872
rect 27062 27860 27068 27872
rect 27023 27832 27068 27860
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 27525 27863 27583 27869
rect 27525 27829 27537 27863
rect 27571 27860 27583 27863
rect 29454 27860 29460 27872
rect 27571 27832 29460 27860
rect 27571 27829 27583 27832
rect 27525 27823 27583 27829
rect 29454 27820 29460 27832
rect 29512 27820 29518 27872
rect 47026 27860 47032 27872
rect 46987 27832 47032 27860
rect 47026 27820 47032 27832
rect 47084 27820 47090 27872
rect 47670 27860 47676 27872
rect 47631 27832 47676 27860
rect 47670 27820 47676 27832
rect 47728 27820 47734 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 12066 27616 12072 27668
rect 12124 27656 12130 27668
rect 12161 27659 12219 27665
rect 12161 27656 12173 27659
rect 12124 27628 12173 27656
rect 12124 27616 12130 27628
rect 12161 27625 12173 27628
rect 12207 27625 12219 27659
rect 13170 27656 13176 27668
rect 12161 27619 12219 27625
rect 12406 27628 13176 27656
rect 9766 27520 9772 27532
rect 9416 27492 9772 27520
rect 9416 27461 9444 27492
rect 9766 27480 9772 27492
rect 9824 27520 9830 27532
rect 10870 27520 10876 27532
rect 9824 27492 10876 27520
rect 9824 27480 9830 27492
rect 10870 27480 10876 27492
rect 10928 27480 10934 27532
rect 11977 27523 12035 27529
rect 11977 27489 11989 27523
rect 12023 27520 12035 27523
rect 12406 27520 12434 27628
rect 12023 27492 12434 27520
rect 12023 27489 12035 27492
rect 11977 27483 12035 27489
rect 9401 27455 9459 27461
rect 9401 27421 9413 27455
rect 9447 27421 9459 27455
rect 9401 27415 9459 27421
rect 10594 27412 10600 27464
rect 10652 27452 10658 27464
rect 12912 27461 12940 27628
rect 13170 27616 13176 27628
rect 13228 27656 13234 27668
rect 15838 27656 15844 27668
rect 13228 27628 15844 27656
rect 13228 27616 13234 27628
rect 13078 27548 13084 27600
rect 13136 27588 13142 27600
rect 13265 27591 13323 27597
rect 13265 27588 13277 27591
rect 13136 27560 13277 27588
rect 13136 27548 13142 27560
rect 13265 27557 13277 27560
rect 13311 27557 13323 27591
rect 13265 27551 13323 27557
rect 13998 27548 14004 27600
rect 14056 27588 14062 27600
rect 14093 27591 14151 27597
rect 14093 27588 14105 27591
rect 14056 27560 14105 27588
rect 14056 27548 14062 27560
rect 14093 27557 14105 27560
rect 14139 27557 14151 27591
rect 14093 27551 14151 27557
rect 11793 27455 11851 27461
rect 11793 27452 11805 27455
rect 10652 27424 11805 27452
rect 10652 27412 10658 27424
rect 11793 27421 11805 27424
rect 11839 27421 11851 27455
rect 11793 27415 11851 27421
rect 12161 27455 12219 27461
rect 12161 27421 12173 27455
rect 12207 27452 12219 27455
rect 12713 27455 12771 27461
rect 12207 27424 12241 27452
rect 12207 27421 12219 27424
rect 12161 27415 12219 27421
rect 12713 27421 12725 27455
rect 12759 27421 12771 27455
rect 12713 27415 12771 27421
rect 12897 27455 12955 27461
rect 12897 27421 12909 27455
rect 12943 27421 12955 27455
rect 13262 27452 13268 27464
rect 12897 27415 12955 27421
rect 13004 27424 13268 27452
rect 11974 27344 11980 27396
rect 12032 27384 12038 27396
rect 12176 27384 12204 27415
rect 12728 27384 12756 27415
rect 13004 27384 13032 27424
rect 13262 27412 13268 27424
rect 13320 27452 13326 27464
rect 14277 27455 14335 27461
rect 14277 27452 14289 27455
rect 13320 27424 14289 27452
rect 13320 27412 13326 27424
rect 14277 27421 14289 27424
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27452 14427 27455
rect 14476 27452 14504 27628
rect 15838 27616 15844 27628
rect 15896 27616 15902 27668
rect 16850 27616 16856 27668
rect 16908 27656 16914 27668
rect 17037 27659 17095 27665
rect 17037 27656 17049 27659
rect 16908 27628 17049 27656
rect 16908 27616 16914 27628
rect 17037 27625 17049 27628
rect 17083 27625 17095 27659
rect 17037 27619 17095 27625
rect 22281 27659 22339 27665
rect 22281 27625 22293 27659
rect 22327 27656 22339 27659
rect 22370 27656 22376 27668
rect 22327 27628 22376 27656
rect 22327 27625 22339 27628
rect 22281 27619 22339 27625
rect 22370 27616 22376 27628
rect 22428 27616 22434 27668
rect 26513 27659 26571 27665
rect 26513 27625 26525 27659
rect 26559 27656 26571 27659
rect 27062 27656 27068 27668
rect 26559 27628 27068 27656
rect 26559 27625 26571 27628
rect 26513 27619 26571 27625
rect 27062 27616 27068 27628
rect 27120 27616 27126 27668
rect 28350 27616 28356 27668
rect 28408 27656 28414 27668
rect 30006 27656 30012 27668
rect 28408 27628 30012 27656
rect 28408 27616 28414 27628
rect 30006 27616 30012 27628
rect 30064 27616 30070 27668
rect 43530 27616 43536 27668
rect 43588 27656 43594 27668
rect 46198 27656 46204 27668
rect 43588 27628 46204 27656
rect 43588 27616 43594 27628
rect 46198 27616 46204 27628
rect 46256 27616 46262 27668
rect 23109 27591 23167 27597
rect 23109 27588 23121 27591
rect 15580 27560 23121 27588
rect 15580 27529 15608 27560
rect 23109 27557 23121 27560
rect 23155 27588 23167 27591
rect 25590 27588 25596 27600
rect 23155 27560 25596 27588
rect 23155 27557 23167 27560
rect 23109 27551 23167 27557
rect 25590 27548 25596 27560
rect 25648 27548 25654 27600
rect 28905 27591 28963 27597
rect 28905 27557 28917 27591
rect 28951 27557 28963 27591
rect 30650 27588 30656 27600
rect 28905 27551 28963 27557
rect 29759 27560 30656 27588
rect 15565 27523 15623 27529
rect 15565 27489 15577 27523
rect 15611 27489 15623 27523
rect 22186 27520 22192 27532
rect 22147 27492 22192 27520
rect 15565 27483 15623 27489
rect 22186 27480 22192 27492
rect 22244 27480 22250 27532
rect 26881 27523 26939 27529
rect 26881 27489 26893 27523
rect 26927 27520 26939 27523
rect 27246 27520 27252 27532
rect 26927 27492 27252 27520
rect 26927 27489 26939 27492
rect 26881 27483 26939 27489
rect 27246 27480 27252 27492
rect 27304 27480 27310 27532
rect 28920 27520 28948 27551
rect 29759 27520 29787 27560
rect 30650 27548 30656 27560
rect 30708 27548 30714 27600
rect 30834 27588 30840 27600
rect 30795 27560 30840 27588
rect 30834 27548 30840 27560
rect 30892 27548 30898 27600
rect 28920 27492 29787 27520
rect 15746 27452 15752 27464
rect 14415 27424 14504 27452
rect 15707 27424 15752 27452
rect 14415 27421 14427 27424
rect 14369 27415 14427 27421
rect 15746 27412 15752 27424
rect 15804 27412 15810 27464
rect 16945 27455 17003 27461
rect 16945 27421 16957 27455
rect 16991 27452 17003 27455
rect 17770 27452 17776 27464
rect 16991 27424 17776 27452
rect 16991 27421 17003 27424
rect 16945 27415 17003 27421
rect 17770 27412 17776 27424
rect 17828 27412 17834 27464
rect 22281 27455 22339 27461
rect 22281 27421 22293 27455
rect 22327 27421 22339 27455
rect 22281 27415 22339 27421
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27421 22983 27455
rect 22925 27415 22983 27421
rect 23661 27455 23719 27461
rect 23661 27421 23673 27455
rect 23707 27452 23719 27455
rect 23750 27452 23756 27464
rect 23707 27424 23756 27452
rect 23707 27421 23719 27424
rect 23661 27415 23719 27421
rect 12032 27356 13032 27384
rect 13081 27387 13139 27393
rect 12032 27344 12038 27356
rect 13081 27353 13093 27387
rect 13127 27384 13139 27387
rect 13538 27384 13544 27396
rect 13127 27356 13544 27384
rect 13127 27353 13139 27356
rect 13081 27347 13139 27353
rect 13538 27344 13544 27356
rect 13596 27344 13602 27396
rect 13906 27344 13912 27396
rect 13964 27384 13970 27396
rect 14461 27387 14519 27393
rect 14461 27384 14473 27387
rect 13964 27356 14473 27384
rect 13964 27344 13970 27356
rect 14461 27353 14473 27356
rect 14507 27353 14519 27387
rect 14461 27347 14519 27353
rect 22005 27387 22063 27393
rect 22005 27353 22017 27387
rect 22051 27353 22063 27387
rect 22296 27384 22324 27415
rect 22738 27384 22744 27396
rect 22296 27356 22744 27384
rect 22005 27347 22063 27353
rect 9122 27276 9128 27328
rect 9180 27316 9186 27328
rect 9401 27319 9459 27325
rect 9401 27316 9413 27319
rect 9180 27288 9413 27316
rect 9180 27276 9186 27288
rect 9401 27285 9413 27288
rect 9447 27285 9459 27319
rect 9401 27279 9459 27285
rect 10870 27276 10876 27328
rect 10928 27316 10934 27328
rect 11885 27319 11943 27325
rect 11885 27316 11897 27319
rect 10928 27288 11897 27316
rect 10928 27276 10934 27288
rect 11885 27285 11897 27288
rect 11931 27316 11943 27319
rect 12989 27319 13047 27325
rect 12989 27316 13001 27319
rect 11931 27288 13001 27316
rect 11931 27285 11943 27288
rect 11885 27279 11943 27285
rect 12989 27285 13001 27288
rect 13035 27316 13047 27319
rect 13924 27316 13952 27344
rect 14642 27316 14648 27328
rect 13035 27288 13952 27316
rect 14603 27288 14648 27316
rect 13035 27285 13047 27288
rect 12989 27279 13047 27285
rect 14642 27276 14648 27288
rect 14700 27276 14706 27328
rect 15930 27316 15936 27328
rect 15891 27288 15936 27316
rect 15930 27276 15936 27288
rect 15988 27276 15994 27328
rect 22020 27316 22048 27347
rect 22738 27344 22744 27356
rect 22796 27344 22802 27396
rect 22278 27316 22284 27328
rect 22020 27288 22284 27316
rect 22278 27276 22284 27288
rect 22336 27276 22342 27328
rect 22465 27319 22523 27325
rect 22465 27285 22477 27319
rect 22511 27316 22523 27319
rect 22646 27316 22652 27328
rect 22511 27288 22652 27316
rect 22511 27285 22523 27288
rect 22465 27279 22523 27285
rect 22646 27276 22652 27288
rect 22704 27316 22710 27328
rect 22940 27316 22968 27415
rect 23750 27412 23756 27424
rect 23808 27412 23814 27464
rect 24210 27412 24216 27464
rect 24268 27452 24274 27464
rect 24489 27455 24547 27461
rect 24489 27452 24501 27455
rect 24268 27424 24501 27452
rect 24268 27412 24274 27424
rect 24489 27421 24501 27424
rect 24535 27421 24547 27455
rect 24489 27415 24547 27421
rect 26697 27455 26755 27461
rect 26697 27421 26709 27455
rect 26743 27452 26755 27455
rect 26786 27452 26792 27464
rect 26743 27424 26792 27452
rect 26743 27421 26755 27424
rect 26697 27415 26755 27421
rect 26786 27412 26792 27424
rect 26844 27412 26850 27464
rect 26970 27412 26976 27464
rect 27028 27452 27034 27464
rect 28721 27455 28779 27461
rect 27028 27424 27073 27452
rect 27028 27412 27034 27424
rect 28721 27421 28733 27455
rect 28767 27452 28779 27455
rect 28902 27452 28908 27464
rect 28767 27424 28908 27452
rect 28767 27421 28779 27424
rect 28721 27415 28779 27421
rect 28902 27412 28908 27424
rect 28960 27412 28966 27464
rect 29454 27412 29460 27464
rect 29512 27452 29518 27464
rect 29549 27455 29607 27461
rect 29828 27455 29886 27461
rect 29549 27452 29561 27455
rect 29512 27424 29561 27452
rect 29512 27412 29518 27424
rect 29549 27421 29561 27424
rect 29595 27421 29607 27455
rect 29549 27415 29607 27421
rect 29737 27449 29795 27455
rect 29737 27415 29749 27449
rect 29783 27415 29795 27449
rect 29828 27421 29840 27455
rect 29874 27421 29886 27455
rect 29828 27415 29886 27421
rect 29917 27455 29975 27461
rect 29917 27421 29929 27455
rect 29963 27421 29975 27455
rect 29917 27415 29975 27421
rect 29737 27409 29795 27415
rect 27982 27344 27988 27396
rect 28040 27384 28046 27396
rect 28166 27384 28172 27396
rect 28040 27356 28172 27384
rect 28040 27344 28046 27356
rect 28166 27344 28172 27356
rect 28224 27384 28230 27396
rect 28224 27356 28994 27384
rect 28224 27344 28230 27356
rect 22704 27288 22968 27316
rect 22704 27276 22710 27288
rect 23382 27276 23388 27328
rect 23440 27316 23446 27328
rect 23753 27319 23811 27325
rect 23753 27316 23765 27319
rect 23440 27288 23765 27316
rect 23440 27276 23446 27288
rect 23753 27285 23765 27288
rect 23799 27285 23811 27319
rect 23753 27279 23811 27285
rect 24673 27319 24731 27325
rect 24673 27285 24685 27319
rect 24719 27316 24731 27319
rect 25682 27316 25688 27328
rect 24719 27288 25688 27316
rect 24719 27285 24731 27288
rect 24673 27279 24731 27285
rect 25682 27276 25688 27288
rect 25740 27316 25746 27328
rect 25866 27316 25872 27328
rect 25740 27288 25872 27316
rect 25740 27276 25746 27288
rect 25866 27276 25872 27288
rect 25924 27276 25930 27328
rect 28966 27316 28994 27356
rect 29759 27316 29787 27409
rect 29843 27328 29871 27415
rect 29932 27384 29960 27415
rect 30006 27412 30012 27464
rect 30064 27461 30070 27464
rect 30064 27455 30113 27461
rect 30064 27421 30067 27455
rect 30101 27421 30113 27455
rect 30668 27452 30696 27548
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27520 46351 27523
rect 47026 27520 47032 27532
rect 46339 27492 47032 27520
rect 46339 27489 46351 27492
rect 46293 27483 46351 27489
rect 47026 27480 47032 27492
rect 47084 27480 47090 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 30745 27455 30803 27461
rect 30745 27452 30757 27455
rect 30668 27424 30757 27452
rect 30064 27415 30113 27421
rect 30745 27421 30757 27424
rect 30791 27421 30803 27455
rect 30745 27415 30803 27421
rect 30064 27412 30070 27415
rect 40402 27384 40408 27396
rect 29932 27356 40408 27384
rect 40402 27344 40408 27356
rect 40460 27344 40466 27396
rect 46477 27387 46535 27393
rect 46477 27353 46489 27387
rect 46523 27384 46535 27387
rect 47670 27384 47676 27396
rect 46523 27356 47676 27384
rect 46523 27353 46535 27356
rect 46477 27347 46535 27353
rect 47670 27344 47676 27356
rect 47728 27344 47734 27396
rect 28966 27288 29787 27316
rect 29822 27276 29828 27328
rect 29880 27276 29886 27328
rect 30098 27276 30104 27328
rect 30156 27316 30162 27328
rect 30285 27319 30343 27325
rect 30285 27316 30297 27319
rect 30156 27288 30297 27316
rect 30156 27276 30162 27288
rect 30285 27285 30297 27288
rect 30331 27285 30343 27319
rect 30285 27279 30343 27285
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 1762 27072 1768 27124
rect 1820 27112 1826 27124
rect 1820 27084 23612 27112
rect 1820 27072 1826 27084
rect 10410 27004 10416 27056
rect 10468 27004 10474 27056
rect 13633 27047 13691 27053
rect 13633 27044 13645 27047
rect 12820 27016 13645 27044
rect 12820 26988 12848 27016
rect 13633 27013 13645 27016
rect 13679 27013 13691 27047
rect 14642 27044 14648 27056
rect 13633 27007 13691 27013
rect 13740 27016 14648 27044
rect 9122 26976 9128 26988
rect 9083 26948 9128 26976
rect 9122 26936 9128 26948
rect 9180 26936 9186 26988
rect 12802 26976 12808 26988
rect 12715 26948 12808 26976
rect 12802 26936 12808 26948
rect 12860 26936 12866 26988
rect 12986 26976 12992 26988
rect 12947 26948 12992 26976
rect 12986 26936 12992 26948
rect 13044 26936 13050 26988
rect 13538 26976 13544 26988
rect 13499 26948 13544 26976
rect 13538 26936 13544 26948
rect 13596 26936 13602 26988
rect 13740 26985 13768 27016
rect 14642 27004 14648 27016
rect 14700 27044 14706 27056
rect 15194 27044 15200 27056
rect 14700 27016 15200 27044
rect 14700 27004 14706 27016
rect 15194 27004 15200 27016
rect 15252 27004 15258 27056
rect 16114 27004 16120 27056
rect 16172 27044 16178 27056
rect 16172 27016 17080 27044
rect 16172 27004 16178 27016
rect 13725 26979 13783 26985
rect 13725 26945 13737 26979
rect 13771 26945 13783 26979
rect 13725 26939 13783 26945
rect 13814 26936 13820 26988
rect 13872 26976 13878 26988
rect 15381 26979 15439 26985
rect 15381 26976 15393 26979
rect 13872 26948 15393 26976
rect 13872 26936 13878 26948
rect 15381 26945 15393 26948
rect 15427 26976 15439 26979
rect 15930 26976 15936 26988
rect 15427 26948 15936 26976
rect 15427 26945 15439 26948
rect 15381 26939 15439 26945
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 16574 26936 16580 26988
rect 16632 26976 16638 26988
rect 16669 26979 16727 26985
rect 16669 26976 16681 26979
rect 16632 26948 16681 26976
rect 16632 26936 16638 26948
rect 16669 26945 16681 26948
rect 16715 26945 16727 26979
rect 16669 26939 16727 26945
rect 16853 26979 16911 26985
rect 16853 26945 16865 26979
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 9398 26908 9404 26920
rect 9359 26880 9404 26908
rect 9398 26868 9404 26880
rect 9456 26868 9462 26920
rect 13081 26911 13139 26917
rect 13081 26877 13093 26911
rect 13127 26908 13139 26911
rect 13998 26908 14004 26920
rect 13127 26880 14004 26908
rect 13127 26877 13139 26880
rect 13081 26871 13139 26877
rect 13998 26868 14004 26880
rect 14056 26868 14062 26920
rect 16868 26908 16896 26939
rect 16868 26880 16988 26908
rect 10594 26800 10600 26852
rect 10652 26840 10658 26852
rect 15565 26843 15623 26849
rect 15565 26840 15577 26843
rect 10652 26812 15577 26840
rect 10652 26800 10658 26812
rect 15565 26809 15577 26812
rect 15611 26840 15623 26843
rect 15654 26840 15660 26852
rect 15611 26812 15660 26840
rect 15611 26809 15623 26812
rect 15565 26803 15623 26809
rect 15654 26800 15660 26812
rect 15712 26840 15718 26852
rect 16758 26840 16764 26852
rect 15712 26812 16764 26840
rect 15712 26800 15718 26812
rect 16758 26800 16764 26812
rect 16816 26800 16822 26852
rect 10870 26772 10876 26784
rect 10831 26744 10876 26772
rect 10870 26732 10876 26744
rect 10928 26732 10934 26784
rect 12066 26732 12072 26784
rect 12124 26772 12130 26784
rect 12621 26775 12679 26781
rect 12621 26772 12633 26775
rect 12124 26744 12633 26772
rect 12124 26732 12130 26744
rect 12621 26741 12633 26744
rect 12667 26741 12679 26775
rect 12621 26735 12679 26741
rect 16390 26732 16396 26784
rect 16448 26772 16454 26784
rect 16669 26775 16727 26781
rect 16669 26772 16681 26775
rect 16448 26744 16681 26772
rect 16448 26732 16454 26744
rect 16669 26741 16681 26744
rect 16715 26741 16727 26775
rect 16960 26772 16988 26880
rect 17052 26840 17080 27016
rect 22370 27004 22376 27056
rect 22428 27044 22434 27056
rect 22428 27016 22508 27044
rect 22428 27004 22434 27016
rect 20714 26936 20720 26988
rect 20772 26976 20778 26988
rect 22189 26979 22247 26985
rect 22189 26976 22201 26979
rect 20772 26948 22201 26976
rect 20772 26936 20778 26948
rect 22189 26945 22201 26948
rect 22235 26945 22247 26979
rect 22189 26939 22247 26945
rect 22278 26936 22284 26988
rect 22336 26976 22342 26988
rect 22480 26985 22508 27016
rect 22465 26979 22523 26985
rect 22336 26948 22381 26976
rect 22336 26936 22342 26948
rect 22465 26945 22477 26979
rect 22511 26945 22523 26979
rect 22465 26939 22523 26945
rect 22649 26979 22707 26985
rect 22649 26945 22661 26979
rect 22695 26976 22707 26979
rect 22738 26976 22744 26988
rect 22695 26948 22744 26976
rect 22695 26945 22707 26948
rect 22649 26939 22707 26945
rect 22738 26936 22744 26948
rect 22796 26936 22802 26988
rect 23477 26979 23535 26985
rect 23477 26945 23489 26979
rect 23523 26945 23535 26979
rect 23584 26976 23612 27084
rect 24210 27072 24216 27124
rect 24268 27112 24274 27124
rect 24581 27115 24639 27121
rect 24581 27112 24593 27115
rect 24268 27084 24593 27112
rect 24268 27072 24274 27084
rect 24581 27081 24593 27084
rect 24627 27081 24639 27115
rect 24581 27075 24639 27081
rect 24670 27072 24676 27124
rect 24728 27112 24734 27124
rect 29822 27112 29828 27124
rect 24728 27084 28028 27112
rect 24728 27072 24734 27084
rect 23661 27047 23719 27053
rect 23661 27013 23673 27047
rect 23707 27044 23719 27047
rect 24854 27044 24860 27056
rect 23707 27016 24860 27044
rect 23707 27013 23719 27016
rect 23661 27007 23719 27013
rect 24854 27004 24860 27016
rect 24912 27004 24918 27056
rect 26786 27004 26792 27056
rect 26844 27044 26850 27056
rect 28000 27053 28028 27084
rect 28966 27084 29828 27112
rect 27985 27047 28043 27053
rect 26844 27016 27292 27044
rect 26844 27004 26850 27016
rect 23753 26979 23811 26985
rect 23753 26976 23765 26979
rect 23584 26948 23765 26976
rect 23477 26939 23535 26945
rect 23753 26945 23765 26948
rect 23799 26945 23811 26979
rect 23753 26939 23811 26945
rect 24673 26979 24731 26985
rect 24673 26945 24685 26979
rect 24719 26976 24731 26979
rect 25774 26976 25780 26988
rect 24719 26948 25780 26976
rect 24719 26945 24731 26948
rect 24673 26939 24731 26945
rect 23492 26908 23520 26939
rect 25774 26936 25780 26948
rect 25832 26936 25838 26988
rect 26053 26979 26111 26985
rect 26053 26945 26065 26979
rect 26099 26976 26111 26979
rect 26878 26976 26884 26988
rect 26099 26948 26884 26976
rect 26099 26945 26111 26948
rect 26053 26939 26111 26945
rect 26878 26936 26884 26948
rect 26936 26936 26942 26988
rect 26970 26936 26976 26988
rect 27028 26976 27034 26988
rect 27264 26985 27292 27016
rect 27985 27013 27997 27047
rect 28031 27013 28043 27047
rect 27985 27007 28043 27013
rect 28169 27047 28227 27053
rect 28169 27013 28181 27047
rect 28215 27044 28227 27047
rect 28350 27044 28356 27056
rect 28215 27016 28356 27044
rect 28215 27013 28227 27016
rect 28169 27007 28227 27013
rect 28350 27004 28356 27016
rect 28408 27004 28414 27056
rect 28966 27044 28994 27084
rect 29822 27072 29828 27084
rect 29880 27112 29886 27124
rect 31573 27115 31631 27121
rect 31573 27112 31585 27115
rect 29880 27084 31585 27112
rect 29880 27072 29886 27084
rect 31573 27081 31585 27084
rect 31619 27081 31631 27115
rect 31573 27075 31631 27081
rect 30098 27044 30104 27056
rect 28828 27016 28994 27044
rect 30059 27016 30104 27044
rect 27249 26979 27307 26985
rect 27028 26948 27073 26976
rect 27028 26936 27034 26948
rect 27249 26945 27261 26979
rect 27295 26976 27307 26979
rect 28828 26976 28856 27016
rect 30098 27004 30104 27016
rect 30156 27004 30162 27056
rect 32217 27047 32275 27053
rect 32217 27044 32229 27047
rect 31326 27016 32229 27044
rect 32217 27013 32229 27016
rect 32263 27013 32275 27047
rect 32217 27007 32275 27013
rect 27295 26948 28856 26976
rect 27295 26945 27307 26948
rect 27249 26939 27307 26945
rect 29730 26936 29736 26988
rect 29788 26976 29794 26988
rect 29825 26979 29883 26985
rect 29825 26976 29837 26979
rect 29788 26948 29837 26976
rect 29788 26936 29794 26948
rect 29825 26945 29837 26948
rect 29871 26945 29883 26979
rect 32122 26976 32128 26988
rect 32083 26948 32128 26976
rect 29825 26939 29883 26945
rect 32122 26936 32128 26948
rect 32180 26936 32186 26988
rect 24765 26911 24823 26917
rect 23492 26880 24256 26908
rect 22094 26840 22100 26852
rect 17052 26812 22100 26840
rect 22094 26800 22100 26812
rect 22152 26800 22158 26852
rect 22186 26800 22192 26852
rect 22244 26840 22250 26852
rect 24228 26849 24256 26880
rect 24765 26877 24777 26911
rect 24811 26908 24823 26911
rect 25314 26908 25320 26920
rect 24811 26880 25320 26908
rect 24811 26877 24823 26880
rect 24765 26871 24823 26877
rect 25314 26868 25320 26880
rect 25372 26868 25378 26920
rect 26145 26911 26203 26917
rect 26145 26877 26157 26911
rect 26191 26877 26203 26911
rect 26145 26871 26203 26877
rect 27157 26911 27215 26917
rect 27157 26877 27169 26911
rect 27203 26908 27215 26911
rect 28258 26908 28264 26920
rect 27203 26880 28264 26908
rect 27203 26877 27215 26880
rect 27157 26871 27215 26877
rect 22373 26843 22431 26849
rect 22373 26840 22385 26843
rect 22244 26812 22385 26840
rect 22244 26800 22250 26812
rect 22373 26809 22385 26812
rect 22419 26809 22431 26843
rect 22373 26803 22431 26809
rect 24213 26843 24271 26849
rect 24213 26809 24225 26843
rect 24259 26809 24271 26843
rect 26160 26840 26188 26871
rect 28258 26868 28264 26880
rect 28316 26868 28322 26920
rect 27246 26840 27252 26852
rect 26160 26812 27252 26840
rect 24213 26803 24271 26809
rect 27246 26800 27252 26812
rect 27304 26800 27310 26852
rect 27430 26840 27436 26852
rect 27391 26812 27436 26840
rect 27430 26800 27436 26812
rect 27488 26800 27494 26852
rect 20806 26772 20812 26784
rect 16960 26744 20812 26772
rect 16669 26735 16727 26741
rect 20806 26732 20812 26744
rect 20864 26772 20870 26784
rect 21913 26775 21971 26781
rect 21913 26772 21925 26775
rect 20864 26744 21925 26772
rect 20864 26732 20870 26744
rect 21913 26741 21925 26744
rect 21959 26741 21971 26775
rect 21913 26735 21971 26741
rect 23293 26775 23351 26781
rect 23293 26741 23305 26775
rect 23339 26772 23351 26775
rect 23750 26772 23756 26784
rect 23339 26744 23756 26772
rect 23339 26741 23351 26744
rect 23293 26735 23351 26741
rect 23750 26732 23756 26744
rect 23808 26732 23814 26784
rect 25682 26732 25688 26784
rect 25740 26772 25746 26784
rect 26329 26775 26387 26781
rect 26329 26772 26341 26775
rect 25740 26744 26341 26772
rect 25740 26732 25746 26744
rect 26329 26741 26341 26744
rect 26375 26741 26387 26775
rect 26329 26735 26387 26741
rect 26878 26732 26884 26784
rect 26936 26772 26942 26784
rect 26973 26775 27031 26781
rect 26973 26772 26985 26775
rect 26936 26744 26985 26772
rect 26936 26732 26942 26744
rect 26973 26741 26985 26744
rect 27019 26741 27031 26775
rect 26973 26735 27031 26741
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 9398 26528 9404 26580
rect 9456 26568 9462 26580
rect 10229 26571 10287 26577
rect 10229 26568 10241 26571
rect 9456 26540 10241 26568
rect 9456 26528 9462 26540
rect 10229 26537 10241 26540
rect 10275 26537 10287 26571
rect 10229 26531 10287 26537
rect 13541 26571 13599 26577
rect 13541 26537 13553 26571
rect 13587 26568 13599 26571
rect 13998 26568 14004 26580
rect 13587 26540 14004 26568
rect 13587 26537 13599 26540
rect 13541 26531 13599 26537
rect 13998 26528 14004 26540
rect 14056 26528 14062 26580
rect 15381 26571 15439 26577
rect 15381 26537 15393 26571
rect 15427 26568 15439 26571
rect 16574 26568 16580 26580
rect 15427 26540 16580 26568
rect 15427 26537 15439 26540
rect 15381 26531 15439 26537
rect 16574 26528 16580 26540
rect 16632 26528 16638 26580
rect 22097 26571 22155 26577
rect 22097 26537 22109 26571
rect 22143 26568 22155 26571
rect 22278 26568 22284 26580
rect 22143 26540 22284 26568
rect 22143 26537 22155 26540
rect 22097 26531 22155 26537
rect 22278 26528 22284 26540
rect 22336 26528 22342 26580
rect 24946 26568 24952 26580
rect 24907 26540 24952 26568
rect 24946 26528 24952 26540
rect 25004 26528 25010 26580
rect 26602 26528 26608 26580
rect 26660 26568 26666 26580
rect 27617 26571 27675 26577
rect 26660 26540 27568 26568
rect 26660 26528 26666 26540
rect 20533 26503 20591 26509
rect 20533 26469 20545 26503
rect 20579 26469 20591 26503
rect 23658 26500 23664 26512
rect 20533 26463 20591 26469
rect 21192 26472 23664 26500
rect 9953 26435 10011 26441
rect 9953 26401 9965 26435
rect 9999 26432 10011 26435
rect 10594 26432 10600 26444
rect 9999 26404 10600 26432
rect 9999 26401 10011 26404
rect 9953 26395 10011 26401
rect 10594 26392 10600 26404
rect 10652 26392 10658 26444
rect 12066 26432 12072 26444
rect 12027 26404 12072 26432
rect 12066 26392 12072 26404
rect 12124 26392 12130 26444
rect 16022 26432 16028 26444
rect 15396 26404 16028 26432
rect 9861 26367 9919 26373
rect 9861 26333 9873 26367
rect 9907 26364 9919 26367
rect 10870 26364 10876 26376
rect 9907 26336 10876 26364
rect 9907 26333 9919 26336
rect 9861 26327 9919 26333
rect 10870 26324 10876 26336
rect 10928 26324 10934 26376
rect 11793 26367 11851 26373
rect 11793 26333 11805 26367
rect 11839 26333 11851 26367
rect 14090 26364 14096 26376
rect 14051 26336 14096 26364
rect 11793 26327 11851 26333
rect 11808 26296 11836 26327
rect 14090 26324 14096 26336
rect 14148 26324 14154 26376
rect 15396 26373 15424 26404
rect 16022 26392 16028 26404
rect 16080 26392 16086 26444
rect 16390 26432 16396 26444
rect 16351 26404 16396 26432
rect 16390 26392 16396 26404
rect 16448 26392 16454 26444
rect 15381 26367 15439 26373
rect 15381 26333 15393 26367
rect 15427 26333 15439 26367
rect 15654 26364 15660 26376
rect 15615 26336 15660 26364
rect 15381 26327 15439 26333
rect 15654 26324 15660 26336
rect 15712 26324 15718 26376
rect 16117 26367 16175 26373
rect 16117 26333 16129 26367
rect 16163 26333 16175 26367
rect 16117 26327 16175 26333
rect 14185 26299 14243 26305
rect 14185 26296 14197 26299
rect 11808 26268 12434 26296
rect 13294 26268 14197 26296
rect 12406 26228 12434 26268
rect 14185 26265 14197 26268
rect 14231 26265 14243 26299
rect 14185 26259 14243 26265
rect 15565 26299 15623 26305
rect 15565 26265 15577 26299
rect 15611 26296 15623 26299
rect 16132 26296 16160 26327
rect 17494 26324 17500 26376
rect 17552 26324 17558 26376
rect 18322 26364 18328 26376
rect 18283 26336 18328 26364
rect 18322 26324 18328 26336
rect 18380 26324 18386 26376
rect 19889 26367 19947 26373
rect 19889 26333 19901 26367
rect 19935 26364 19947 26367
rect 20548 26364 20576 26463
rect 21192 26441 21220 26472
rect 23658 26460 23664 26472
rect 23716 26500 23722 26512
rect 24670 26500 24676 26512
rect 23716 26472 24676 26500
rect 23716 26460 23722 26472
rect 24670 26460 24676 26472
rect 24728 26460 24734 26512
rect 27154 26500 27160 26512
rect 25240 26472 27160 26500
rect 21177 26435 21235 26441
rect 21177 26401 21189 26435
rect 21223 26401 21235 26435
rect 21177 26395 21235 26401
rect 23382 26392 23388 26444
rect 23440 26432 23446 26444
rect 24765 26435 24823 26441
rect 24765 26432 24777 26435
rect 23440 26404 24777 26432
rect 23440 26392 23446 26404
rect 24765 26401 24777 26404
rect 24811 26401 24823 26435
rect 24765 26395 24823 26401
rect 19935 26336 20576 26364
rect 20901 26367 20959 26373
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 20901 26333 20913 26367
rect 20947 26364 20959 26367
rect 21634 26364 21640 26376
rect 20947 26336 21640 26364
rect 20947 26333 20959 26336
rect 20901 26327 20959 26333
rect 21634 26324 21640 26336
rect 21692 26324 21698 26376
rect 22094 26324 22100 26376
rect 22152 26364 22158 26376
rect 24397 26367 24455 26373
rect 24397 26364 24409 26367
rect 22152 26336 24409 26364
rect 22152 26324 22158 26336
rect 24397 26333 24409 26336
rect 24443 26333 24455 26367
rect 24397 26327 24455 26333
rect 24555 26367 24613 26373
rect 24555 26333 24567 26367
rect 24601 26364 24613 26367
rect 25240 26364 25268 26472
rect 27154 26460 27160 26472
rect 27212 26500 27218 26512
rect 27430 26500 27436 26512
rect 27212 26472 27436 26500
rect 27212 26460 27218 26472
rect 27430 26460 27436 26472
rect 27488 26460 27494 26512
rect 27540 26500 27568 26540
rect 27617 26537 27629 26571
rect 27663 26568 27675 26571
rect 28629 26571 28687 26577
rect 28629 26568 28641 26571
rect 27663 26540 28641 26568
rect 27663 26537 27675 26540
rect 27617 26531 27675 26537
rect 28629 26537 28641 26540
rect 28675 26537 28687 26571
rect 28629 26531 28687 26537
rect 47118 26500 47124 26512
rect 27540 26472 47124 26500
rect 25314 26392 25320 26444
rect 25372 26432 25378 26444
rect 26970 26432 26976 26444
rect 25372 26404 26976 26432
rect 25372 26392 25378 26404
rect 26970 26392 26976 26404
rect 27028 26432 27034 26444
rect 32324 26441 32352 26472
rect 47118 26460 47124 26472
rect 47176 26460 47182 26512
rect 32309 26435 32367 26441
rect 27028 26404 28488 26432
rect 27028 26392 27034 26404
rect 25682 26364 25688 26376
rect 24601 26336 25268 26364
rect 25643 26336 25688 26364
rect 24601 26333 24613 26336
rect 24555 26327 24613 26333
rect 25682 26324 25688 26336
rect 25740 26324 25746 26376
rect 25774 26324 25780 26376
rect 25832 26364 25838 26376
rect 26053 26367 26111 26373
rect 26053 26364 26065 26367
rect 25832 26336 26065 26364
rect 25832 26324 25838 26336
rect 26053 26333 26065 26336
rect 26099 26333 26111 26367
rect 27246 26364 27252 26376
rect 27207 26336 27252 26364
rect 26053 26327 26111 26333
rect 27246 26324 27252 26336
rect 27304 26324 27310 26376
rect 27430 26324 27436 26376
rect 27488 26364 27494 26376
rect 27525 26367 27583 26373
rect 27525 26364 27537 26367
rect 27488 26336 27537 26364
rect 27488 26324 27494 26336
rect 27525 26333 27537 26336
rect 27571 26333 27583 26367
rect 28258 26364 28264 26376
rect 28219 26336 28264 26364
rect 27525 26327 27583 26333
rect 28258 26324 28264 26336
rect 28316 26324 28322 26376
rect 28460 26373 28488 26404
rect 32309 26401 32321 26435
rect 32355 26401 32367 26435
rect 32309 26395 32367 26401
rect 46293 26435 46351 26441
rect 46293 26401 46305 26435
rect 46339 26432 46351 26435
rect 46934 26432 46940 26444
rect 46339 26404 46940 26432
rect 46339 26401 46351 26404
rect 46293 26395 46351 26401
rect 46934 26392 46940 26404
rect 46992 26392 46998 26444
rect 47762 26432 47768 26444
rect 47723 26404 47768 26432
rect 47762 26392 47768 26404
rect 47820 26392 47826 26444
rect 28445 26367 28503 26373
rect 28445 26333 28457 26367
rect 28491 26333 28503 26367
rect 28445 26327 28503 26333
rect 31297 26367 31355 26373
rect 31297 26333 31309 26367
rect 31343 26364 31355 26367
rect 32033 26367 32091 26373
rect 32033 26364 32045 26367
rect 31343 26336 32045 26364
rect 31343 26333 31355 26336
rect 31297 26327 31355 26333
rect 32033 26333 32045 26336
rect 32079 26364 32091 26367
rect 32122 26364 32128 26376
rect 32079 26336 32128 26364
rect 32079 26333 32091 26336
rect 32033 26327 32091 26333
rect 32122 26324 32128 26336
rect 32180 26324 32186 26376
rect 16666 26296 16672 26308
rect 15611 26268 16068 26296
rect 16132 26268 16672 26296
rect 15611 26265 15623 26268
rect 15565 26259 15623 26265
rect 12710 26228 12716 26240
rect 12406 26200 12716 26228
rect 12710 26188 12716 26200
rect 12768 26188 12774 26240
rect 16040 26228 16068 26268
rect 16666 26256 16672 26268
rect 16724 26256 16730 26308
rect 21266 26256 21272 26308
rect 21324 26296 21330 26308
rect 21729 26299 21787 26305
rect 21729 26296 21741 26299
rect 21324 26268 21741 26296
rect 21324 26256 21330 26268
rect 21729 26265 21741 26268
rect 21775 26265 21787 26299
rect 21729 26259 21787 26265
rect 21818 26256 21824 26308
rect 21876 26296 21882 26308
rect 21913 26299 21971 26305
rect 21913 26296 21925 26299
rect 21876 26268 21925 26296
rect 21876 26256 21882 26268
rect 21913 26265 21925 26268
rect 21959 26265 21971 26299
rect 25866 26296 25872 26308
rect 25827 26268 25872 26296
rect 21913 26259 21971 26265
rect 25866 26256 25872 26268
rect 25924 26256 25930 26308
rect 25961 26299 26019 26305
rect 25961 26265 25973 26299
rect 26007 26296 26019 26299
rect 26878 26296 26884 26308
rect 26007 26268 26884 26296
rect 26007 26265 26019 26268
rect 25961 26259 26019 26265
rect 26878 26256 26884 26268
rect 26936 26256 26942 26308
rect 31389 26299 31447 26305
rect 31389 26265 31401 26299
rect 31435 26296 31447 26299
rect 32306 26296 32312 26308
rect 31435 26268 32312 26296
rect 31435 26265 31447 26268
rect 31389 26259 31447 26265
rect 32306 26256 32312 26268
rect 32364 26256 32370 26308
rect 43438 26256 43444 26308
rect 43496 26296 43502 26308
rect 46290 26296 46296 26308
rect 43496 26268 46296 26296
rect 43496 26256 43502 26268
rect 46290 26256 46296 26268
rect 46348 26256 46354 26308
rect 46477 26299 46535 26305
rect 46477 26265 46489 26299
rect 46523 26296 46535 26299
rect 48038 26296 48044 26308
rect 46523 26268 48044 26296
rect 46523 26265 46535 26268
rect 46477 26259 46535 26265
rect 48038 26256 48044 26268
rect 48096 26256 48102 26308
rect 16758 26228 16764 26240
rect 16040 26200 16764 26228
rect 16758 26188 16764 26200
rect 16816 26188 16822 26240
rect 17862 26228 17868 26240
rect 17823 26200 17868 26228
rect 17862 26188 17868 26200
rect 17920 26188 17926 26240
rect 18417 26231 18475 26237
rect 18417 26197 18429 26231
rect 18463 26228 18475 26231
rect 18506 26228 18512 26240
rect 18463 26200 18512 26228
rect 18463 26197 18475 26200
rect 18417 26191 18475 26197
rect 18506 26188 18512 26200
rect 18564 26188 18570 26240
rect 19426 26188 19432 26240
rect 19484 26228 19490 26240
rect 19705 26231 19763 26237
rect 19705 26228 19717 26231
rect 19484 26200 19717 26228
rect 19484 26188 19490 26200
rect 19705 26197 19717 26200
rect 19751 26197 19763 26231
rect 19705 26191 19763 26197
rect 20990 26188 20996 26240
rect 21048 26228 21054 26240
rect 26234 26228 26240 26240
rect 21048 26200 21093 26228
rect 26195 26200 26240 26228
rect 21048 26188 21054 26200
rect 26234 26188 26240 26200
rect 26292 26188 26298 26240
rect 27801 26231 27859 26237
rect 27801 26197 27813 26231
rect 27847 26228 27859 26231
rect 27982 26228 27988 26240
rect 27847 26200 27988 26228
rect 27847 26197 27859 26200
rect 27801 26191 27859 26197
rect 27982 26188 27988 26200
rect 28040 26188 28046 26240
rect 32030 26188 32036 26240
rect 32088 26228 32094 26240
rect 45646 26228 45652 26240
rect 32088 26200 45652 26228
rect 32088 26188 32094 26200
rect 45646 26188 45652 26200
rect 45704 26188 45710 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 10321 26027 10379 26033
rect 10321 25993 10333 26027
rect 10367 26024 10379 26027
rect 10410 26024 10416 26036
rect 10367 25996 10416 26024
rect 10367 25993 10379 25996
rect 10321 25987 10379 25993
rect 10410 25984 10416 25996
rect 10468 25984 10474 26036
rect 12710 26024 12716 26036
rect 12671 25996 12716 26024
rect 12710 25984 12716 25996
rect 12768 25984 12774 26036
rect 15746 26024 15752 26036
rect 15707 25996 15752 26024
rect 15746 25984 15752 25996
rect 15804 25984 15810 26036
rect 16758 25984 16764 26036
rect 16816 26024 16822 26036
rect 17037 26027 17095 26033
rect 17037 26024 17049 26027
rect 16816 25996 17049 26024
rect 16816 25984 16822 25996
rect 17037 25993 17049 25996
rect 17083 25993 17095 26027
rect 17037 25987 17095 25993
rect 17221 26027 17279 26033
rect 17221 25993 17233 26027
rect 17267 26024 17279 26027
rect 20714 26024 20720 26036
rect 17267 25996 20720 26024
rect 17267 25993 17279 25996
rect 17221 25987 17279 25993
rect 20714 25984 20720 25996
rect 20772 25984 20778 26036
rect 46198 26024 46204 26036
rect 22066 25996 46204 26024
rect 16022 25916 16028 25968
rect 16080 25956 16086 25968
rect 16574 25956 16580 25968
rect 16080 25928 16580 25956
rect 16080 25916 16086 25928
rect 16574 25916 16580 25928
rect 16632 25956 16638 25968
rect 16669 25959 16727 25965
rect 16669 25956 16681 25959
rect 16632 25928 16681 25956
rect 16632 25916 16638 25928
rect 16669 25925 16681 25928
rect 16715 25956 16727 25959
rect 17862 25956 17868 25968
rect 16715 25928 17868 25956
rect 16715 25925 16727 25928
rect 16669 25919 16727 25925
rect 17862 25916 17868 25928
rect 17920 25916 17926 25968
rect 18506 25956 18512 25968
rect 18467 25928 18512 25956
rect 18506 25916 18512 25928
rect 18564 25916 18570 25968
rect 20165 25959 20223 25965
rect 20165 25925 20177 25959
rect 20211 25956 20223 25959
rect 22066 25956 22094 25996
rect 46198 25984 46204 25996
rect 46256 25984 46262 26036
rect 26970 25956 26976 25968
rect 20211 25928 22094 25956
rect 26931 25928 26976 25956
rect 20211 25925 20223 25928
rect 20165 25919 20223 25925
rect 26970 25916 26976 25928
rect 27028 25916 27034 25968
rect 27246 25916 27252 25968
rect 27304 25956 27310 25968
rect 27341 25959 27399 25965
rect 27341 25956 27353 25959
rect 27304 25928 27353 25956
rect 27304 25916 27310 25928
rect 27341 25925 27353 25928
rect 27387 25925 27399 25959
rect 27341 25919 27399 25925
rect 28350 25916 28356 25968
rect 28408 25956 28414 25968
rect 28408 25928 28580 25956
rect 28408 25916 28414 25928
rect 10226 25888 10232 25900
rect 10187 25860 10232 25888
rect 10226 25848 10232 25860
rect 10284 25848 10290 25900
rect 12621 25891 12679 25897
rect 12621 25857 12633 25891
rect 12667 25888 12679 25891
rect 13446 25888 13452 25900
rect 12667 25860 13452 25888
rect 12667 25857 12679 25860
rect 12621 25851 12679 25857
rect 13446 25848 13452 25860
rect 13504 25848 13510 25900
rect 15562 25888 15568 25900
rect 15523 25860 15568 25888
rect 15562 25848 15568 25860
rect 15620 25848 15626 25900
rect 16853 25891 16911 25897
rect 16853 25886 16865 25891
rect 16776 25858 16865 25886
rect 15102 25780 15108 25832
rect 15160 25820 15166 25832
rect 15381 25823 15439 25829
rect 15381 25820 15393 25823
rect 15160 25792 15393 25820
rect 15160 25780 15166 25792
rect 15381 25789 15393 25792
rect 15427 25820 15439 25823
rect 16776 25820 16804 25858
rect 16853 25857 16865 25858
rect 16899 25857 16911 25891
rect 16853 25851 16911 25857
rect 16945 25891 17003 25897
rect 16945 25857 16957 25891
rect 16991 25857 17003 25891
rect 16945 25851 17003 25857
rect 20993 25891 21051 25897
rect 20993 25857 21005 25891
rect 21039 25888 21051 25891
rect 21726 25888 21732 25900
rect 21039 25860 21732 25888
rect 21039 25857 21051 25860
rect 20993 25851 21051 25857
rect 15427 25792 16804 25820
rect 15427 25789 15439 25792
rect 15381 25783 15439 25789
rect 15562 25712 15568 25764
rect 15620 25752 15626 25764
rect 16960 25752 16988 25851
rect 21726 25848 21732 25860
rect 21784 25848 21790 25900
rect 21818 25848 21824 25900
rect 21876 25888 21882 25900
rect 22281 25891 22339 25897
rect 22281 25888 22293 25891
rect 21876 25860 21921 25888
rect 22066 25860 22293 25888
rect 21876 25848 21882 25860
rect 18322 25820 18328 25832
rect 18283 25792 18328 25820
rect 18322 25780 18328 25792
rect 18380 25780 18386 25832
rect 21266 25820 21272 25832
rect 21227 25792 21272 25820
rect 21266 25780 21272 25792
rect 21324 25820 21330 25832
rect 22066 25820 22094 25860
rect 22281 25857 22293 25860
rect 22327 25857 22339 25891
rect 22281 25851 22339 25857
rect 27157 25891 27215 25897
rect 27157 25857 27169 25891
rect 27203 25857 27215 25891
rect 27982 25888 27988 25900
rect 27943 25860 27988 25888
rect 27157 25851 27215 25857
rect 21324 25792 22094 25820
rect 22189 25823 22247 25829
rect 21324 25780 21330 25792
rect 22189 25789 22201 25823
rect 22235 25820 22247 25823
rect 22462 25820 22468 25832
rect 22235 25792 22468 25820
rect 22235 25789 22247 25792
rect 22189 25783 22247 25789
rect 15620 25724 16988 25752
rect 21085 25755 21143 25761
rect 15620 25712 15626 25724
rect 21085 25721 21097 25755
rect 21131 25752 21143 25755
rect 22094 25752 22100 25764
rect 21131 25724 22100 25752
rect 21131 25721 21143 25724
rect 21085 25715 21143 25721
rect 22094 25712 22100 25724
rect 22152 25752 22158 25764
rect 22204 25752 22232 25783
rect 22462 25780 22468 25792
rect 22520 25780 22526 25832
rect 27172 25820 27200 25851
rect 27982 25848 27988 25860
rect 28040 25848 28046 25900
rect 28166 25888 28172 25900
rect 28127 25860 28172 25888
rect 28166 25848 28172 25860
rect 28224 25848 28230 25900
rect 28552 25897 28580 25928
rect 32122 25916 32128 25968
rect 32180 25916 32186 25968
rect 32306 25956 32312 25968
rect 32267 25928 32312 25956
rect 32306 25916 32312 25928
rect 32364 25916 32370 25968
rect 33965 25959 34023 25965
rect 33965 25925 33977 25959
rect 34011 25956 34023 25959
rect 43438 25956 43444 25968
rect 34011 25928 43444 25956
rect 34011 25925 34023 25928
rect 33965 25919 34023 25925
rect 43438 25916 43444 25928
rect 43496 25916 43502 25968
rect 28537 25891 28595 25897
rect 28537 25857 28549 25891
rect 28583 25857 28595 25891
rect 28537 25851 28595 25857
rect 30929 25891 30987 25897
rect 30929 25857 30941 25891
rect 30975 25888 30987 25891
rect 32140 25888 32168 25916
rect 30975 25860 32168 25888
rect 30975 25857 30987 25860
rect 30929 25851 30987 25857
rect 45646 25848 45652 25900
rect 45704 25888 45710 25900
rect 46569 25891 46627 25897
rect 46569 25888 46581 25891
rect 45704 25860 46581 25888
rect 45704 25848 45710 25860
rect 46569 25857 46581 25860
rect 46615 25857 46627 25891
rect 46569 25851 46627 25857
rect 28258 25820 28264 25832
rect 27172 25792 28264 25820
rect 28258 25780 28264 25792
rect 28316 25780 28322 25832
rect 28350 25780 28356 25832
rect 28408 25820 28414 25832
rect 31294 25820 31300 25832
rect 28408 25792 28453 25820
rect 31255 25792 31300 25820
rect 28408 25780 28414 25792
rect 31294 25780 31300 25792
rect 31352 25780 31358 25832
rect 32125 25823 32183 25829
rect 32125 25789 32137 25823
rect 32171 25789 32183 25823
rect 47394 25820 47400 25832
rect 32125 25783 32183 25789
rect 35866 25792 47400 25820
rect 23382 25752 23388 25764
rect 22152 25724 22245 25752
rect 22296 25724 23388 25752
rect 22152 25712 22158 25724
rect 22296 25696 22324 25724
rect 23382 25712 23388 25724
rect 23440 25712 23446 25764
rect 24026 25712 24032 25764
rect 24084 25752 24090 25764
rect 32140 25752 32168 25783
rect 24084 25724 32168 25752
rect 24084 25712 24090 25724
rect 21174 25684 21180 25696
rect 21135 25656 21180 25684
rect 21174 25644 21180 25656
rect 21232 25644 21238 25696
rect 22278 25684 22284 25696
rect 22191 25656 22284 25684
rect 22278 25644 22284 25656
rect 22336 25644 22342 25696
rect 22465 25687 22523 25693
rect 22465 25653 22477 25687
rect 22511 25684 22523 25687
rect 22738 25684 22744 25696
rect 22511 25656 22744 25684
rect 22511 25653 22523 25656
rect 22465 25647 22523 25653
rect 22738 25644 22744 25656
rect 22796 25644 22802 25696
rect 27522 25644 27528 25696
rect 27580 25684 27586 25696
rect 28721 25687 28779 25693
rect 28721 25684 28733 25687
rect 27580 25656 28733 25684
rect 27580 25644 27586 25656
rect 28721 25653 28733 25656
rect 28767 25653 28779 25687
rect 28721 25647 28779 25653
rect 31294 25644 31300 25696
rect 31352 25684 31358 25696
rect 35866 25684 35894 25792
rect 47394 25780 47400 25792
rect 47452 25780 47458 25832
rect 46290 25712 46296 25764
rect 46348 25752 46354 25764
rect 47765 25755 47823 25761
rect 47765 25752 47777 25755
rect 46348 25724 47777 25752
rect 46348 25712 46354 25724
rect 47765 25721 47777 25724
rect 47811 25721 47823 25755
rect 47765 25715 47823 25721
rect 31352 25656 35894 25684
rect 31352 25644 31358 25656
rect 46474 25644 46480 25696
rect 46532 25684 46538 25696
rect 46661 25687 46719 25693
rect 46661 25684 46673 25687
rect 46532 25656 46673 25684
rect 46532 25644 46538 25656
rect 46661 25653 46673 25656
rect 46707 25653 46719 25687
rect 46661 25647 46719 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 16666 25480 16672 25492
rect 16627 25452 16672 25480
rect 16666 25440 16672 25452
rect 16724 25440 16730 25492
rect 17494 25440 17500 25492
rect 17552 25480 17558 25492
rect 17589 25483 17647 25489
rect 17589 25480 17601 25483
rect 17552 25452 17601 25480
rect 17552 25440 17558 25452
rect 17589 25449 17601 25452
rect 17635 25449 17647 25483
rect 17589 25443 17647 25449
rect 20990 25440 20996 25492
rect 21048 25480 21054 25492
rect 21453 25483 21511 25489
rect 21453 25480 21465 25483
rect 21048 25452 21465 25480
rect 21048 25440 21054 25452
rect 21453 25449 21465 25452
rect 21499 25449 21511 25483
rect 22278 25480 22284 25492
rect 21453 25443 21511 25449
rect 21744 25452 22284 25480
rect 21744 25424 21772 25452
rect 22278 25440 22284 25452
rect 22336 25440 22342 25492
rect 28258 25440 28264 25492
rect 28316 25480 28322 25492
rect 28997 25483 29055 25489
rect 28997 25480 29009 25483
rect 28316 25452 29009 25480
rect 28316 25440 28322 25452
rect 28997 25449 29009 25452
rect 29043 25449 29055 25483
rect 28997 25443 29055 25449
rect 21726 25412 21732 25424
rect 21687 25384 21732 25412
rect 21726 25372 21732 25384
rect 21784 25372 21790 25424
rect 21821 25415 21879 25421
rect 21821 25381 21833 25415
rect 21867 25412 21879 25415
rect 22094 25412 22100 25424
rect 21867 25384 22100 25412
rect 21867 25381 21879 25384
rect 21821 25375 21879 25381
rect 22094 25372 22100 25384
rect 22152 25372 22158 25424
rect 22465 25415 22523 25421
rect 22465 25381 22477 25415
rect 22511 25412 22523 25415
rect 22554 25412 22560 25424
rect 22511 25384 22560 25412
rect 22511 25381 22523 25384
rect 22465 25375 22523 25381
rect 22554 25372 22560 25384
rect 22612 25372 22618 25424
rect 12713 25347 12771 25353
rect 12713 25313 12725 25347
rect 12759 25344 12771 25347
rect 12802 25344 12808 25356
rect 12759 25316 12808 25344
rect 12759 25313 12771 25316
rect 12713 25307 12771 25313
rect 12802 25304 12808 25316
rect 12860 25304 12866 25356
rect 18322 25344 18328 25356
rect 15764 25316 18328 25344
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 9858 25276 9864 25288
rect 9819 25248 9864 25276
rect 9858 25236 9864 25248
rect 9916 25236 9922 25288
rect 12342 25236 12348 25288
rect 12400 25276 12406 25288
rect 12621 25279 12679 25285
rect 12621 25276 12633 25279
rect 12400 25248 12633 25276
rect 12400 25236 12406 25248
rect 12621 25245 12633 25248
rect 12667 25245 12679 25279
rect 12621 25239 12679 25245
rect 15470 25236 15476 25288
rect 15528 25276 15534 25288
rect 15764 25285 15792 25316
rect 18322 25304 18328 25316
rect 18380 25304 18386 25356
rect 20993 25347 21051 25353
rect 20993 25313 21005 25347
rect 21039 25344 21051 25347
rect 26234 25344 26240 25356
rect 21039 25316 21772 25344
rect 21039 25313 21051 25316
rect 20993 25307 21051 25313
rect 21744 25288 21772 25316
rect 25332 25316 26240 25344
rect 15749 25279 15807 25285
rect 15749 25276 15761 25279
rect 15528 25248 15761 25276
rect 15528 25236 15534 25248
rect 15749 25245 15761 25248
rect 15795 25245 15807 25279
rect 15749 25239 15807 25245
rect 15838 25236 15844 25288
rect 15896 25276 15902 25288
rect 16025 25279 16083 25285
rect 16025 25276 16037 25279
rect 15896 25248 16037 25276
rect 15896 25236 15902 25248
rect 16025 25245 16037 25248
rect 16071 25245 16083 25279
rect 16574 25276 16580 25288
rect 16535 25248 16580 25276
rect 16025 25239 16083 25245
rect 16574 25236 16580 25248
rect 16632 25236 16638 25288
rect 17494 25276 17500 25288
rect 17455 25248 17500 25276
rect 17494 25236 17500 25248
rect 17552 25236 17558 25288
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25276 18567 25279
rect 18598 25276 18604 25288
rect 18555 25248 18604 25276
rect 18555 25245 18567 25248
rect 18509 25239 18567 25245
rect 18598 25236 18604 25248
rect 18656 25236 18662 25288
rect 19242 25276 19248 25288
rect 19203 25248 19248 25276
rect 19242 25236 19248 25248
rect 19300 25236 19306 25288
rect 21266 25236 21272 25288
rect 21324 25276 21330 25288
rect 21637 25279 21695 25285
rect 21637 25276 21649 25279
rect 21324 25248 21649 25276
rect 21324 25236 21330 25248
rect 21637 25245 21649 25248
rect 21683 25245 21695 25279
rect 21637 25239 21695 25245
rect 21726 25236 21732 25288
rect 21784 25236 21790 25288
rect 21902 25279 21960 25285
rect 21902 25245 21914 25279
rect 21948 25245 21960 25279
rect 22738 25276 22744 25288
rect 22699 25248 22744 25276
rect 21902 25239 21960 25245
rect 1670 25208 1676 25220
rect 1631 25180 1676 25208
rect 1670 25168 1676 25180
rect 1728 25168 1734 25220
rect 10134 25208 10140 25220
rect 10095 25180 10140 25208
rect 10134 25168 10140 25180
rect 10192 25168 10198 25220
rect 11422 25208 11428 25220
rect 11362 25180 11428 25208
rect 11422 25168 11428 25180
rect 11480 25168 11486 25220
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 19521 25211 19579 25217
rect 19521 25208 19533 25211
rect 19484 25180 19533 25208
rect 19484 25168 19490 25180
rect 19521 25177 19533 25180
rect 19567 25177 19579 25211
rect 21744 25208 21772 25236
rect 21928 25208 21956 25239
rect 22738 25236 22744 25248
rect 22796 25236 22802 25288
rect 25332 25285 25360 25316
rect 26234 25304 26240 25316
rect 26292 25304 26298 25356
rect 46474 25344 46480 25356
rect 46435 25316 46480 25344
rect 46474 25304 46480 25316
rect 46532 25304 46538 25356
rect 48130 25344 48136 25356
rect 48091 25316 48136 25344
rect 48130 25304 48136 25316
rect 48188 25304 48194 25356
rect 25317 25279 25375 25285
rect 25317 25245 25329 25279
rect 25363 25245 25375 25279
rect 25590 25276 25596 25288
rect 25551 25248 25596 25276
rect 25317 25239 25375 25245
rect 25590 25236 25596 25248
rect 25648 25236 25654 25288
rect 27246 25276 27252 25288
rect 27207 25248 27252 25276
rect 27246 25236 27252 25248
rect 27304 25236 27310 25288
rect 31481 25279 31539 25285
rect 31481 25245 31493 25279
rect 31527 25276 31539 25279
rect 32122 25276 32128 25288
rect 31527 25248 32128 25276
rect 31527 25245 31539 25248
rect 31481 25239 31539 25245
rect 32122 25236 32128 25248
rect 32180 25236 32186 25288
rect 45646 25276 45652 25288
rect 45607 25248 45652 25276
rect 45646 25236 45652 25248
rect 45704 25236 45710 25288
rect 46293 25279 46351 25285
rect 46293 25245 46305 25279
rect 46339 25245 46351 25279
rect 46293 25239 46351 25245
rect 19521 25171 19579 25177
rect 19628 25180 20010 25208
rect 21744 25180 21956 25208
rect 22465 25211 22523 25217
rect 11054 25100 11060 25152
rect 11112 25140 11118 25152
rect 11609 25143 11667 25149
rect 11609 25140 11621 25143
rect 11112 25112 11621 25140
rect 11112 25100 11118 25112
rect 11609 25109 11621 25112
rect 11655 25109 11667 25143
rect 12986 25140 12992 25152
rect 12947 25112 12992 25140
rect 11609 25103 11667 25109
rect 12986 25100 12992 25112
rect 13044 25100 13050 25152
rect 15562 25140 15568 25152
rect 15523 25112 15568 25140
rect 15562 25100 15568 25112
rect 15620 25100 15626 25152
rect 15654 25100 15660 25152
rect 15712 25140 15718 25152
rect 15933 25143 15991 25149
rect 15933 25140 15945 25143
rect 15712 25112 15945 25140
rect 15712 25100 15718 25112
rect 15933 25109 15945 25112
rect 15979 25109 15991 25143
rect 15933 25103 15991 25109
rect 18601 25143 18659 25149
rect 18601 25109 18613 25143
rect 18647 25140 18659 25143
rect 19628 25140 19656 25180
rect 22465 25177 22477 25211
rect 22511 25208 22523 25211
rect 22830 25208 22836 25220
rect 22511 25180 22836 25208
rect 22511 25177 22523 25180
rect 22465 25171 22523 25177
rect 22830 25168 22836 25180
rect 22888 25208 22894 25220
rect 24854 25208 24860 25220
rect 22888 25180 24860 25208
rect 22888 25168 22894 25180
rect 24854 25168 24860 25180
rect 24912 25208 24918 25220
rect 25501 25211 25559 25217
rect 25501 25208 25513 25211
rect 24912 25180 25513 25208
rect 24912 25168 24918 25180
rect 25501 25177 25513 25180
rect 25547 25177 25559 25211
rect 27522 25208 27528 25220
rect 27483 25180 27528 25208
rect 25501 25171 25559 25177
rect 27522 25168 27528 25180
rect 27580 25168 27586 25220
rect 28074 25168 28080 25220
rect 28132 25168 28138 25220
rect 31202 25168 31208 25220
rect 31260 25208 31266 25220
rect 31297 25211 31355 25217
rect 31297 25208 31309 25211
rect 31260 25180 31309 25208
rect 31260 25168 31266 25180
rect 31297 25177 31309 25180
rect 31343 25208 31355 25211
rect 32766 25208 32772 25220
rect 31343 25180 31754 25208
rect 32679 25180 32772 25208
rect 31343 25177 31355 25180
rect 31297 25171 31355 25177
rect 18647 25112 19656 25140
rect 18647 25109 18659 25112
rect 18601 25103 18659 25109
rect 21174 25100 21180 25152
rect 21232 25140 21238 25152
rect 22649 25143 22707 25149
rect 22649 25140 22661 25143
rect 21232 25112 22661 25140
rect 21232 25100 21238 25112
rect 22649 25109 22661 25112
rect 22695 25109 22707 25143
rect 22649 25103 22707 25109
rect 25133 25143 25191 25149
rect 25133 25109 25145 25143
rect 25179 25140 25191 25143
rect 25406 25140 25412 25152
rect 25179 25112 25412 25140
rect 25179 25109 25191 25112
rect 25133 25103 25191 25109
rect 25406 25100 25412 25112
rect 25464 25100 25470 25152
rect 31726 25140 31754 25180
rect 32766 25168 32772 25180
rect 32824 25208 32830 25220
rect 43070 25208 43076 25220
rect 32824 25180 43076 25208
rect 32824 25168 32830 25180
rect 43070 25168 43076 25180
rect 43128 25168 43134 25220
rect 46308 25208 46336 25239
rect 46566 25208 46572 25220
rect 46308 25180 46572 25208
rect 46566 25168 46572 25180
rect 46624 25168 46630 25220
rect 41230 25140 41236 25152
rect 31726 25112 41236 25140
rect 41230 25100 41236 25112
rect 41288 25140 41294 25152
rect 45554 25140 45560 25152
rect 41288 25112 45560 25140
rect 41288 25100 41294 25112
rect 45554 25100 45560 25112
rect 45612 25100 45618 25152
rect 45741 25143 45799 25149
rect 45741 25109 45753 25143
rect 45787 25140 45799 25143
rect 46014 25140 46020 25152
rect 45787 25112 46020 25140
rect 45787 25109 45799 25112
rect 45741 25103 45799 25109
rect 46014 25100 46020 25112
rect 46072 25100 46078 25152
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 9858 24936 9864 24948
rect 9819 24908 9864 24936
rect 9858 24896 9864 24908
rect 9916 24896 9922 24948
rect 10134 24896 10140 24948
rect 10192 24936 10198 24948
rect 10505 24939 10563 24945
rect 10505 24936 10517 24939
rect 10192 24908 10517 24936
rect 10192 24896 10198 24908
rect 10505 24905 10517 24908
rect 10551 24905 10563 24939
rect 10505 24899 10563 24905
rect 11698 24896 11704 24948
rect 11756 24936 11762 24948
rect 12342 24936 12348 24948
rect 11756 24908 12348 24936
rect 11756 24896 11762 24908
rect 12342 24896 12348 24908
rect 12400 24936 12406 24948
rect 14553 24939 14611 24945
rect 14553 24936 14565 24939
rect 12400 24908 14565 24936
rect 12400 24896 12406 24908
rect 14553 24905 14565 24908
rect 14599 24936 14611 24939
rect 15286 24936 15292 24948
rect 14599 24908 15292 24936
rect 14599 24905 14611 24908
rect 14553 24899 14611 24905
rect 15286 24896 15292 24908
rect 15344 24936 15350 24948
rect 15749 24939 15807 24945
rect 15749 24936 15761 24939
rect 15344 24908 15761 24936
rect 15344 24896 15350 24908
rect 15749 24905 15761 24908
rect 15795 24905 15807 24939
rect 15749 24899 15807 24905
rect 16758 24896 16764 24948
rect 16816 24896 16822 24948
rect 18322 24896 18328 24948
rect 18380 24936 18386 24948
rect 18417 24939 18475 24945
rect 18417 24936 18429 24939
rect 18380 24908 18429 24936
rect 18380 24896 18386 24908
rect 18417 24905 18429 24908
rect 18463 24905 18475 24939
rect 21266 24936 21272 24948
rect 21227 24908 21272 24936
rect 18417 24899 18475 24905
rect 21266 24896 21272 24908
rect 21324 24896 21330 24948
rect 22741 24939 22799 24945
rect 22741 24905 22753 24939
rect 22787 24936 22799 24939
rect 22830 24936 22836 24948
rect 22787 24908 22836 24936
rect 22787 24905 22799 24908
rect 22741 24899 22799 24905
rect 22830 24896 22836 24908
rect 22888 24896 22894 24948
rect 25225 24939 25283 24945
rect 25225 24905 25237 24939
rect 25271 24936 25283 24939
rect 25314 24936 25320 24948
rect 25271 24908 25320 24936
rect 25271 24905 25283 24908
rect 25225 24899 25283 24905
rect 25314 24896 25320 24908
rect 25372 24896 25378 24948
rect 12986 24828 12992 24880
rect 13044 24868 13050 24880
rect 13081 24871 13139 24877
rect 13081 24868 13093 24871
rect 13044 24840 13093 24868
rect 13044 24828 13050 24840
rect 13081 24837 13093 24840
rect 13127 24837 13139 24871
rect 13081 24831 13139 24837
rect 13538 24828 13544 24880
rect 13596 24828 13602 24880
rect 15470 24868 15476 24880
rect 15431 24840 15476 24868
rect 15470 24828 15476 24840
rect 15528 24828 15534 24880
rect 15654 24868 15660 24880
rect 15615 24840 15660 24868
rect 15654 24828 15660 24840
rect 15712 24828 15718 24880
rect 16776 24868 16804 24896
rect 16592 24840 16804 24868
rect 9766 24800 9772 24812
rect 9727 24772 9772 24800
rect 9766 24760 9772 24772
rect 9824 24760 9830 24812
rect 10410 24800 10416 24812
rect 10371 24772 10416 24800
rect 10410 24760 10416 24772
rect 10468 24760 10474 24812
rect 10594 24800 10600 24812
rect 10555 24772 10600 24800
rect 10594 24760 10600 24772
rect 10652 24760 10658 24812
rect 11517 24803 11575 24809
rect 11517 24800 11529 24803
rect 10796 24772 11529 24800
rect 10226 24692 10232 24744
rect 10284 24732 10290 24744
rect 10796 24732 10824 24772
rect 11517 24769 11529 24772
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 15841 24803 15899 24809
rect 15841 24800 15853 24803
rect 15252 24772 15853 24800
rect 15252 24760 15258 24772
rect 15841 24769 15853 24772
rect 15887 24769 15899 24803
rect 15841 24763 15899 24769
rect 16025 24803 16083 24809
rect 16025 24769 16037 24803
rect 16071 24800 16083 24803
rect 16592 24800 16620 24840
rect 17678 24828 17684 24880
rect 17736 24828 17742 24880
rect 20438 24828 20444 24880
rect 20496 24828 20502 24880
rect 24486 24828 24492 24880
rect 24544 24828 24550 24880
rect 22554 24800 22560 24812
rect 16071 24772 16620 24800
rect 22515 24772 22560 24800
rect 16071 24769 16083 24772
rect 16025 24763 16083 24769
rect 22554 24760 22560 24772
rect 22612 24760 22618 24812
rect 22833 24803 22891 24809
rect 22833 24769 22845 24803
rect 22879 24800 22891 24803
rect 23106 24800 23112 24812
rect 22879 24772 23112 24800
rect 22879 24769 22891 24772
rect 22833 24763 22891 24769
rect 23106 24760 23112 24772
rect 23164 24760 23170 24812
rect 25038 24760 25044 24812
rect 25096 24800 25102 24812
rect 26145 24803 26203 24809
rect 26145 24800 26157 24803
rect 25096 24772 26157 24800
rect 25096 24760 25102 24772
rect 26145 24769 26157 24772
rect 26191 24800 26203 24803
rect 27985 24803 28043 24809
rect 27985 24800 27997 24803
rect 26191 24772 27997 24800
rect 26191 24769 26203 24772
rect 26145 24763 26203 24769
rect 27985 24769 27997 24772
rect 28031 24769 28043 24803
rect 27985 24763 28043 24769
rect 28074 24760 28080 24812
rect 28132 24800 28138 24812
rect 32122 24800 32128 24812
rect 28132 24772 28177 24800
rect 32083 24772 32128 24800
rect 28132 24760 28138 24772
rect 32122 24760 32128 24772
rect 32180 24760 32186 24812
rect 10284 24704 10824 24732
rect 10284 24692 10290 24704
rect 11422 24692 11428 24744
rect 11480 24732 11486 24744
rect 11609 24735 11667 24741
rect 11609 24732 11621 24735
rect 11480 24704 11621 24732
rect 11480 24692 11486 24704
rect 11609 24701 11621 24704
rect 11655 24701 11667 24735
rect 11609 24695 11667 24701
rect 12805 24735 12863 24741
rect 12805 24701 12817 24735
rect 12851 24732 12863 24735
rect 14090 24732 14096 24744
rect 12851 24704 14096 24732
rect 12851 24701 12863 24704
rect 12805 24695 12863 24701
rect 14090 24692 14096 24704
rect 14148 24692 14154 24744
rect 16666 24732 16672 24744
rect 16627 24704 16672 24732
rect 16666 24692 16672 24704
rect 16724 24692 16730 24744
rect 16942 24732 16948 24744
rect 16903 24704 16948 24732
rect 16942 24692 16948 24704
rect 17000 24692 17006 24744
rect 19242 24692 19248 24744
rect 19300 24732 19306 24744
rect 19521 24735 19579 24741
rect 19521 24732 19533 24735
rect 19300 24704 19533 24732
rect 19300 24692 19306 24704
rect 19521 24701 19533 24704
rect 19567 24701 19579 24735
rect 19521 24695 19579 24701
rect 19797 24735 19855 24741
rect 19797 24701 19809 24735
rect 19843 24732 19855 24735
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 19843 24704 22385 24732
rect 19843 24701 19855 24704
rect 19797 24695 19855 24701
rect 22373 24701 22385 24704
rect 22419 24701 22431 24735
rect 22373 24695 22431 24701
rect 23477 24735 23535 24741
rect 23477 24701 23489 24735
rect 23523 24701 23535 24735
rect 23750 24732 23756 24744
rect 23711 24704 23756 24732
rect 23477 24695 23535 24701
rect 3510 24624 3516 24676
rect 3568 24664 3574 24676
rect 12526 24664 12532 24676
rect 3568 24636 12532 24664
rect 3568 24624 3574 24636
rect 12526 24624 12532 24636
rect 12584 24624 12590 24676
rect 14108 24636 16804 24664
rect 12434 24556 12440 24608
rect 12492 24596 12498 24608
rect 14108 24596 14136 24636
rect 12492 24568 14136 24596
rect 16776 24596 16804 24636
rect 18414 24596 18420 24608
rect 16776 24568 18420 24596
rect 12492 24556 12498 24568
rect 18414 24556 18420 24568
rect 18472 24556 18478 24608
rect 19536 24596 19564 24695
rect 23492 24664 23520 24695
rect 23750 24692 23756 24704
rect 23808 24692 23814 24744
rect 25222 24692 25228 24744
rect 25280 24692 25286 24744
rect 29270 24692 29276 24744
rect 29328 24732 29334 24744
rect 29365 24735 29423 24741
rect 29365 24732 29377 24735
rect 29328 24704 29377 24732
rect 29328 24692 29334 24704
rect 29365 24701 29377 24704
rect 29411 24701 29423 24735
rect 29365 24695 29423 24701
rect 29549 24735 29607 24741
rect 29549 24701 29561 24735
rect 29595 24732 29607 24735
rect 29638 24732 29644 24744
rect 29595 24704 29644 24732
rect 29595 24701 29607 24704
rect 29549 24695 29607 24701
rect 29638 24692 29644 24704
rect 29696 24692 29702 24744
rect 29822 24732 29828 24744
rect 29783 24704 29828 24732
rect 29822 24692 29828 24704
rect 29880 24692 29886 24744
rect 32030 24692 32036 24744
rect 32088 24732 32094 24744
rect 32309 24735 32367 24741
rect 32309 24732 32321 24735
rect 32088 24704 32321 24732
rect 32088 24692 32094 24704
rect 32309 24701 32321 24704
rect 32355 24701 32367 24735
rect 32309 24695 32367 24701
rect 45189 24735 45247 24741
rect 45189 24701 45201 24735
rect 45235 24701 45247 24735
rect 45370 24732 45376 24744
rect 45331 24704 45376 24732
rect 45189 24695 45247 24701
rect 20824 24636 23520 24664
rect 25240 24664 25268 24692
rect 45002 24664 45008 24676
rect 25240 24636 45008 24664
rect 20824 24596 20852 24636
rect 45002 24624 45008 24636
rect 45060 24624 45066 24676
rect 19536 24568 20852 24596
rect 26237 24599 26295 24605
rect 26237 24565 26249 24599
rect 26283 24596 26295 24599
rect 26418 24596 26424 24608
rect 26283 24568 26424 24596
rect 26283 24565 26295 24568
rect 26237 24559 26295 24565
rect 26418 24556 26424 24568
rect 26476 24556 26482 24608
rect 45204 24596 45232 24695
rect 45370 24692 45376 24704
rect 45428 24692 45434 24744
rect 46842 24732 46848 24744
rect 46803 24704 46848 24732
rect 46842 24692 46848 24704
rect 46900 24692 46906 24744
rect 45278 24624 45284 24676
rect 45336 24664 45342 24676
rect 46198 24664 46204 24676
rect 45336 24636 46204 24664
rect 45336 24624 45342 24636
rect 46198 24624 46204 24636
rect 46256 24624 46262 24676
rect 47765 24599 47823 24605
rect 47765 24596 47777 24599
rect 45204 24568 47777 24596
rect 47765 24565 47777 24568
rect 47811 24565 47823 24599
rect 47765 24559 47823 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 10321 24395 10379 24401
rect 10321 24361 10333 24395
rect 10367 24392 10379 24395
rect 10410 24392 10416 24404
rect 10367 24364 10416 24392
rect 10367 24361 10379 24364
rect 10321 24355 10379 24361
rect 10410 24352 10416 24364
rect 10468 24352 10474 24404
rect 12406 24364 22094 24392
rect 3878 24284 3884 24336
rect 3936 24324 3942 24336
rect 12406 24324 12434 24364
rect 3936 24296 12434 24324
rect 13449 24327 13507 24333
rect 3936 24284 3942 24296
rect 13449 24293 13461 24327
rect 13495 24324 13507 24327
rect 13538 24324 13544 24336
rect 13495 24296 13544 24324
rect 13495 24293 13507 24296
rect 13449 24287 13507 24293
rect 13538 24284 13544 24296
rect 13596 24284 13602 24336
rect 14090 24324 14096 24336
rect 14051 24296 14096 24324
rect 14090 24284 14096 24296
rect 14148 24284 14154 24336
rect 15286 24324 15292 24336
rect 15247 24296 15292 24324
rect 15286 24284 15292 24296
rect 15344 24284 15350 24336
rect 16485 24327 16543 24333
rect 15488 24296 16436 24324
rect 1946 24216 1952 24268
rect 2004 24256 2010 24268
rect 12434 24256 12440 24268
rect 2004 24228 12440 24256
rect 2004 24216 2010 24228
rect 12434 24216 12440 24228
rect 12492 24216 12498 24268
rect 12526 24216 12532 24268
rect 12584 24256 12590 24268
rect 15488 24256 15516 24296
rect 12584 24228 12629 24256
rect 14108 24228 15516 24256
rect 12584 24216 12590 24228
rect 9125 24191 9183 24197
rect 9125 24157 9137 24191
rect 9171 24188 9183 24191
rect 9582 24188 9588 24200
rect 9171 24160 9588 24188
rect 9171 24157 9183 24160
rect 9125 24151 9183 24157
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 9677 24191 9735 24197
rect 9677 24157 9689 24191
rect 9723 24157 9735 24191
rect 9677 24151 9735 24157
rect 9692 24120 9720 24151
rect 10134 24148 10140 24200
rect 10192 24188 10198 24200
rect 10597 24191 10655 24197
rect 10597 24188 10609 24191
rect 10192 24160 10609 24188
rect 10192 24148 10198 24160
rect 10597 24157 10609 24160
rect 10643 24157 10655 24191
rect 11054 24188 11060 24200
rect 11015 24160 11060 24188
rect 10597 24151 10655 24157
rect 11054 24148 11060 24160
rect 11112 24148 11118 24200
rect 12710 24148 12716 24200
rect 12768 24188 12774 24200
rect 13357 24191 13415 24197
rect 13357 24188 13369 24191
rect 12768 24160 13369 24188
rect 12768 24148 12774 24160
rect 13357 24157 13369 24160
rect 13403 24188 13415 24191
rect 13998 24188 14004 24200
rect 13403 24160 14004 24188
rect 13403 24157 13415 24160
rect 13357 24151 13415 24157
rect 13998 24148 14004 24160
rect 14056 24148 14062 24200
rect 14108 24197 14136 24228
rect 15562 24216 15568 24268
rect 15620 24256 15626 24268
rect 16301 24259 16359 24265
rect 16301 24256 16313 24259
rect 15620 24228 16313 24256
rect 15620 24216 15626 24228
rect 16301 24225 16313 24228
rect 16347 24225 16359 24259
rect 16408 24256 16436 24296
rect 16485 24293 16497 24327
rect 16531 24324 16543 24327
rect 16942 24324 16948 24336
rect 16531 24296 16948 24324
rect 16531 24293 16543 24296
rect 16485 24287 16543 24293
rect 16942 24284 16948 24296
rect 17000 24284 17006 24336
rect 17678 24284 17684 24336
rect 17736 24324 17742 24336
rect 17773 24327 17831 24333
rect 17773 24324 17785 24327
rect 17736 24296 17785 24324
rect 17736 24284 17742 24296
rect 17773 24293 17785 24296
rect 17819 24293 17831 24327
rect 20438 24324 20444 24336
rect 20399 24296 20444 24324
rect 17773 24287 17831 24293
rect 20438 24284 20444 24296
rect 20496 24284 20502 24336
rect 22066 24324 22094 24364
rect 24486 24352 24492 24404
rect 24544 24392 24550 24404
rect 24581 24395 24639 24401
rect 24581 24392 24593 24395
rect 24544 24364 24593 24392
rect 24544 24352 24550 24364
rect 24581 24361 24593 24364
rect 24627 24361 24639 24395
rect 24581 24355 24639 24361
rect 24688 24364 31754 24392
rect 24688 24324 24716 24364
rect 26878 24324 26884 24336
rect 22066 24296 24716 24324
rect 26839 24296 26884 24324
rect 26878 24284 26884 24296
rect 26936 24284 26942 24336
rect 29638 24324 29644 24336
rect 29599 24296 29644 24324
rect 29638 24284 29644 24296
rect 29696 24284 29702 24336
rect 31726 24324 31754 24364
rect 33134 24324 33140 24336
rect 31726 24296 33140 24324
rect 33134 24284 33140 24296
rect 33192 24284 33198 24336
rect 16574 24256 16580 24268
rect 16408 24228 16580 24256
rect 16301 24219 16359 24225
rect 16574 24216 16580 24228
rect 16632 24216 16638 24268
rect 18598 24216 18604 24268
rect 18656 24256 18662 24268
rect 25133 24259 25191 24265
rect 18656 24228 20392 24256
rect 18656 24216 18662 24228
rect 14093 24191 14151 24197
rect 14093 24157 14105 24191
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 15657 24191 15715 24197
rect 15657 24157 15669 24191
rect 15703 24188 15715 24191
rect 15746 24188 15752 24200
rect 15703 24160 15752 24188
rect 15703 24157 15715 24160
rect 15657 24151 15715 24157
rect 10226 24120 10232 24132
rect 9692 24092 10232 24120
rect 10226 24080 10232 24092
rect 10284 24080 10290 24132
rect 10321 24123 10379 24129
rect 10321 24089 10333 24123
rect 10367 24120 10379 24123
rect 11072 24120 11100 24148
rect 11238 24120 11244 24132
rect 10367 24092 11100 24120
rect 11199 24092 11244 24120
rect 10367 24089 10379 24092
rect 10321 24083 10379 24089
rect 11238 24080 11244 24092
rect 11296 24080 11302 24132
rect 13446 24080 13452 24132
rect 13504 24120 13510 24132
rect 14108 24120 14136 24151
rect 15746 24148 15752 24160
rect 15804 24148 15810 24200
rect 16761 24191 16819 24197
rect 16761 24157 16773 24191
rect 16807 24188 16819 24191
rect 16850 24188 16856 24200
rect 16807 24160 16856 24188
rect 16807 24157 16819 24160
rect 16761 24151 16819 24157
rect 16850 24148 16856 24160
rect 16908 24148 16914 24200
rect 17494 24148 17500 24200
rect 17552 24188 17558 24200
rect 17681 24191 17739 24197
rect 17681 24188 17693 24191
rect 17552 24160 17693 24188
rect 17552 24148 17558 24160
rect 17681 24157 17693 24160
rect 17727 24157 17739 24191
rect 19426 24188 19432 24200
rect 19387 24160 19432 24188
rect 17681 24151 17739 24157
rect 13504 24092 14136 24120
rect 13504 24080 13510 24092
rect 15194 24080 15200 24132
rect 15252 24120 15258 24132
rect 15565 24123 15623 24129
rect 15565 24120 15577 24123
rect 15252 24092 15577 24120
rect 15252 24080 15258 24092
rect 15565 24089 15577 24092
rect 15611 24089 15623 24123
rect 15565 24083 15623 24089
rect 15930 24080 15936 24132
rect 15988 24120 15994 24132
rect 17696 24120 17724 24151
rect 19426 24148 19432 24160
rect 19484 24148 19490 24200
rect 20364 24197 20392 24228
rect 25133 24225 25145 24259
rect 25179 24256 25191 24259
rect 27246 24256 27252 24268
rect 25179 24228 27252 24256
rect 25179 24225 25191 24228
rect 25133 24219 25191 24225
rect 27246 24216 27252 24228
rect 27304 24216 27310 24268
rect 46014 24256 46020 24268
rect 45975 24228 46020 24256
rect 46014 24216 46020 24228
rect 46072 24216 46078 24268
rect 47302 24256 47308 24268
rect 47263 24228 47308 24256
rect 47302 24216 47308 24228
rect 47360 24216 47366 24268
rect 20349 24191 20407 24197
rect 20349 24157 20361 24191
rect 20395 24157 20407 24191
rect 20349 24151 20407 24157
rect 24489 24191 24547 24197
rect 24489 24157 24501 24191
rect 24535 24188 24547 24191
rect 25038 24188 25044 24200
rect 24535 24160 25044 24188
rect 24535 24157 24547 24160
rect 24489 24151 24547 24157
rect 25038 24148 25044 24160
rect 25096 24148 25102 24200
rect 29178 24148 29184 24200
rect 29236 24188 29242 24200
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 29236 24160 29561 24188
rect 29236 24148 29242 24160
rect 29549 24157 29561 24160
rect 29595 24188 29607 24191
rect 30190 24188 30196 24200
rect 29595 24160 30196 24188
rect 29595 24157 29607 24160
rect 29549 24151 29607 24157
rect 30190 24148 30196 24160
rect 30248 24148 30254 24200
rect 45833 24191 45891 24197
rect 45833 24157 45845 24191
rect 45879 24157 45891 24191
rect 45833 24151 45891 24157
rect 20070 24120 20076 24132
rect 15988 24092 16896 24120
rect 17696 24092 20076 24120
rect 15988 24080 15994 24092
rect 8202 24012 8208 24064
rect 8260 24052 8266 24064
rect 9125 24055 9183 24061
rect 9125 24052 9137 24055
rect 8260 24024 9137 24052
rect 8260 24012 8266 24024
rect 9125 24021 9137 24024
rect 9171 24021 9183 24055
rect 9766 24052 9772 24064
rect 9727 24024 9772 24052
rect 9125 24015 9183 24021
rect 9766 24012 9772 24024
rect 9824 24012 9830 24064
rect 10502 24052 10508 24064
rect 10463 24024 10508 24052
rect 10502 24012 10508 24024
rect 10560 24012 10566 24064
rect 15470 24052 15476 24064
rect 15431 24024 15476 24052
rect 15470 24012 15476 24024
rect 15528 24012 15534 24064
rect 15838 24052 15844 24064
rect 15799 24024 15844 24052
rect 15838 24012 15844 24024
rect 15896 24012 15902 24064
rect 16669 24055 16727 24061
rect 16669 24021 16681 24055
rect 16715 24052 16727 24055
rect 16758 24052 16764 24064
rect 16715 24024 16764 24052
rect 16715 24021 16727 24024
rect 16669 24015 16727 24021
rect 16758 24012 16764 24024
rect 16816 24012 16822 24064
rect 16868 24052 16896 24092
rect 20070 24080 20076 24092
rect 20128 24080 20134 24132
rect 25406 24120 25412 24132
rect 25367 24092 25412 24120
rect 25406 24080 25412 24092
rect 25464 24080 25470 24132
rect 26418 24080 26424 24132
rect 26476 24080 26482 24132
rect 45848 24120 45876 24151
rect 47026 24120 47032 24132
rect 45848 24092 47032 24120
rect 47026 24080 47032 24092
rect 47084 24080 47090 24132
rect 21910 24052 21916 24064
rect 16868 24024 21916 24052
rect 21910 24012 21916 24024
rect 21968 24012 21974 24064
rect 45554 24012 45560 24064
rect 45612 24052 45618 24064
rect 45830 24052 45836 24064
rect 45612 24024 45836 24052
rect 45612 24012 45618 24024
rect 45830 24012 45836 24024
rect 45888 24012 45894 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1946 23848 1952 23860
rect 1907 23820 1952 23848
rect 1946 23808 1952 23820
rect 2004 23808 2010 23860
rect 3418 23808 3424 23860
rect 3476 23848 3482 23860
rect 29822 23848 29828 23860
rect 3476 23820 9904 23848
rect 3476 23808 3482 23820
rect 9766 23780 9772 23792
rect 9706 23752 9772 23780
rect 9766 23740 9772 23752
rect 9824 23740 9830 23792
rect 9876 23780 9904 23820
rect 10060 23820 29828 23848
rect 10060 23780 10088 23820
rect 29822 23808 29828 23820
rect 29880 23808 29886 23860
rect 45370 23808 45376 23860
rect 45428 23848 45434 23860
rect 47673 23851 47731 23857
rect 47673 23848 47685 23851
rect 45428 23820 47685 23848
rect 45428 23808 45434 23820
rect 47673 23817 47685 23820
rect 47719 23817 47731 23851
rect 47673 23811 47731 23817
rect 9876 23752 10088 23780
rect 11054 23740 11060 23792
rect 11112 23780 11118 23792
rect 12161 23783 12219 23789
rect 12161 23780 12173 23783
rect 11112 23752 12173 23780
rect 11112 23740 11118 23752
rect 12161 23749 12173 23752
rect 12207 23749 12219 23783
rect 12161 23743 12219 23749
rect 12377 23783 12435 23789
rect 12377 23749 12389 23783
rect 12423 23780 12435 23783
rect 14550 23780 14556 23792
rect 12423 23752 14556 23780
rect 12423 23749 12435 23752
rect 12377 23743 12435 23749
rect 14550 23740 14556 23752
rect 14608 23740 14614 23792
rect 19352 23752 21864 23780
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 8202 23712 8208 23724
rect 8163 23684 8208 23712
rect 8202 23672 8208 23684
rect 8260 23672 8266 23724
rect 12986 23672 12992 23724
rect 13044 23712 13050 23724
rect 13265 23715 13323 23721
rect 13265 23712 13277 23715
rect 13044 23684 13277 23712
rect 13044 23672 13050 23684
rect 13265 23681 13277 23684
rect 13311 23681 13323 23715
rect 15286 23712 15292 23724
rect 15199 23684 15292 23712
rect 13265 23675 13323 23681
rect 15286 23672 15292 23684
rect 15344 23712 15350 23724
rect 16114 23712 16120 23724
rect 15344 23684 16120 23712
rect 15344 23672 15350 23684
rect 16114 23672 16120 23684
rect 16172 23672 16178 23724
rect 16574 23672 16580 23724
rect 16632 23712 16638 23724
rect 16669 23715 16727 23721
rect 16669 23712 16681 23715
rect 16632 23684 16681 23712
rect 16632 23672 16638 23684
rect 16669 23681 16681 23684
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 17586 23672 17592 23724
rect 17644 23712 17650 23724
rect 19352 23721 19380 23752
rect 21836 23721 21864 23752
rect 21910 23740 21916 23792
rect 21968 23780 21974 23792
rect 25961 23783 26019 23789
rect 21968 23752 25912 23780
rect 21968 23740 21974 23752
rect 18693 23715 18751 23721
rect 18693 23712 18705 23715
rect 17644 23684 18705 23712
rect 17644 23672 17650 23684
rect 18693 23681 18705 23684
rect 18739 23681 18751 23715
rect 18693 23675 18751 23681
rect 19337 23715 19395 23721
rect 19337 23681 19349 23715
rect 19383 23681 19395 23715
rect 20073 23715 20131 23721
rect 20073 23712 20085 23715
rect 19337 23675 19395 23681
rect 19536 23684 20085 23712
rect 8478 23644 8484 23656
rect 8439 23616 8484 23644
rect 8478 23604 8484 23616
rect 8536 23604 8542 23656
rect 9950 23644 9956 23656
rect 9911 23616 9956 23644
rect 9950 23604 9956 23616
rect 10008 23604 10014 23656
rect 15470 23604 15476 23656
rect 15528 23644 15534 23656
rect 15565 23647 15623 23653
rect 15565 23644 15577 23647
rect 15528 23616 15577 23644
rect 15528 23604 15534 23616
rect 15565 23613 15577 23616
rect 15611 23613 15623 23647
rect 15565 23607 15623 23613
rect 17678 23604 17684 23656
rect 17736 23644 17742 23656
rect 17862 23644 17868 23656
rect 17736 23616 17868 23644
rect 17736 23604 17742 23616
rect 17862 23604 17868 23616
rect 17920 23644 17926 23656
rect 19352 23644 19380 23675
rect 17920 23616 19380 23644
rect 17920 23604 17926 23616
rect 9674 23536 9680 23588
rect 9732 23576 9738 23588
rect 10594 23576 10600 23588
rect 9732 23548 10600 23576
rect 9732 23536 9738 23548
rect 10594 23536 10600 23548
rect 10652 23536 10658 23588
rect 12529 23579 12587 23585
rect 12529 23545 12541 23579
rect 12575 23576 12587 23579
rect 15102 23576 15108 23588
rect 12575 23548 15108 23576
rect 12575 23545 12587 23548
rect 12529 23539 12587 23545
rect 15102 23536 15108 23548
rect 15160 23536 15166 23588
rect 16666 23576 16672 23588
rect 16627 23548 16672 23576
rect 16666 23536 16672 23548
rect 16724 23536 16730 23588
rect 18598 23536 18604 23588
rect 18656 23576 18662 23588
rect 19536 23585 19564 23684
rect 20073 23681 20085 23684
rect 20119 23681 20131 23715
rect 20073 23675 20131 23681
rect 21821 23715 21879 23721
rect 21821 23681 21833 23715
rect 21867 23681 21879 23715
rect 22925 23715 22983 23721
rect 22925 23712 22937 23715
rect 21821 23675 21879 23681
rect 22066 23684 22937 23712
rect 22066 23644 22094 23684
rect 22925 23681 22937 23684
rect 22971 23681 22983 23715
rect 22925 23675 22983 23681
rect 23474 23672 23480 23724
rect 23532 23712 23538 23724
rect 25884 23721 25912 23752
rect 25961 23749 25973 23783
rect 26007 23780 26019 23783
rect 27157 23783 27215 23789
rect 27157 23780 27169 23783
rect 26007 23752 27169 23780
rect 26007 23749 26019 23752
rect 25961 23743 26019 23749
rect 27157 23749 27169 23752
rect 27203 23749 27215 23783
rect 27157 23743 27215 23749
rect 28813 23783 28871 23789
rect 28813 23749 28825 23783
rect 28859 23780 28871 23783
rect 37274 23780 37280 23792
rect 28859 23752 37280 23780
rect 28859 23749 28871 23752
rect 28813 23743 28871 23749
rect 37274 23740 37280 23752
rect 37332 23740 37338 23792
rect 23569 23715 23627 23721
rect 23569 23712 23581 23715
rect 23532 23684 23581 23712
rect 23532 23672 23538 23684
rect 23569 23681 23581 23684
rect 23615 23681 23627 23715
rect 23569 23675 23627 23681
rect 23753 23715 23811 23721
rect 23753 23681 23765 23715
rect 23799 23681 23811 23715
rect 23753 23675 23811 23681
rect 25869 23715 25927 23721
rect 25869 23681 25881 23715
rect 25915 23681 25927 23715
rect 25869 23675 25927 23681
rect 20088 23616 22094 23644
rect 20088 23588 20116 23616
rect 23382 23604 23388 23656
rect 23440 23644 23446 23656
rect 23768 23644 23796 23675
rect 28718 23672 28724 23724
rect 28776 23712 28782 23724
rect 30377 23715 30435 23721
rect 30377 23712 30389 23715
rect 28776 23684 30389 23712
rect 28776 23672 28782 23684
rect 30377 23681 30389 23684
rect 30423 23681 30435 23715
rect 30377 23675 30435 23681
rect 31205 23715 31263 23721
rect 31205 23681 31217 23715
rect 31251 23712 31263 23715
rect 45830 23712 45836 23724
rect 31251 23684 31754 23712
rect 45791 23684 45836 23712
rect 31251 23681 31263 23684
rect 31205 23675 31263 23681
rect 23440 23616 23796 23644
rect 23440 23604 23446 23616
rect 23842 23604 23848 23656
rect 23900 23644 23906 23656
rect 26418 23644 26424 23656
rect 23900 23616 26424 23644
rect 23900 23604 23906 23616
rect 26418 23604 26424 23616
rect 26476 23644 26482 23656
rect 26973 23647 27031 23653
rect 26973 23644 26985 23647
rect 26476 23616 26985 23644
rect 26476 23604 26482 23616
rect 26973 23613 26985 23616
rect 27019 23613 27031 23647
rect 31110 23644 31116 23656
rect 31071 23616 31116 23644
rect 26973 23607 27031 23613
rect 31110 23604 31116 23616
rect 31168 23604 31174 23656
rect 31726 23644 31754 23684
rect 45830 23672 45836 23684
rect 45888 23672 45894 23724
rect 46201 23715 46259 23721
rect 46201 23681 46213 23715
rect 46247 23712 46259 23715
rect 46658 23712 46664 23724
rect 46247 23684 46664 23712
rect 46247 23681 46259 23684
rect 46201 23675 46259 23681
rect 46658 23672 46664 23684
rect 46716 23672 46722 23724
rect 47486 23672 47492 23724
rect 47544 23712 47550 23724
rect 47581 23715 47639 23721
rect 47581 23712 47593 23715
rect 47544 23684 47593 23712
rect 47544 23672 47550 23684
rect 47581 23681 47593 23684
rect 47627 23681 47639 23715
rect 47581 23675 47639 23681
rect 32217 23647 32275 23653
rect 32217 23644 32229 23647
rect 31726 23616 32229 23644
rect 32217 23613 32229 23616
rect 32263 23613 32275 23647
rect 32217 23607 32275 23613
rect 32401 23647 32459 23653
rect 32401 23613 32413 23647
rect 32447 23644 32459 23647
rect 33042 23644 33048 23656
rect 32447 23616 33048 23644
rect 32447 23613 32459 23616
rect 32401 23607 32459 23613
rect 19521 23579 19579 23585
rect 19521 23576 19533 23579
rect 18656 23548 19533 23576
rect 18656 23536 18662 23548
rect 19521 23545 19533 23548
rect 19567 23545 19579 23579
rect 19521 23539 19579 23545
rect 20070 23536 20076 23588
rect 20128 23536 20134 23588
rect 22005 23579 22063 23585
rect 22005 23545 22017 23579
rect 22051 23576 22063 23579
rect 23198 23576 23204 23588
rect 22051 23548 23204 23576
rect 22051 23545 22063 23548
rect 22005 23539 22063 23545
rect 23198 23536 23204 23548
rect 23256 23576 23262 23588
rect 28902 23576 28908 23588
rect 23256 23548 28908 23576
rect 23256 23536 23262 23548
rect 28902 23536 28908 23548
rect 28960 23536 28966 23588
rect 30469 23579 30527 23585
rect 30469 23545 30481 23579
rect 30515 23576 30527 23579
rect 31754 23576 31760 23588
rect 30515 23548 31760 23576
rect 30515 23545 30527 23548
rect 30469 23539 30527 23545
rect 31754 23536 31760 23548
rect 31812 23536 31818 23588
rect 32232 23576 32260 23607
rect 33042 23604 33048 23616
rect 33100 23604 33106 23656
rect 33134 23604 33140 23656
rect 33192 23644 33198 23656
rect 44453 23647 44511 23653
rect 33192 23616 33237 23644
rect 33192 23604 33198 23616
rect 44453 23613 44465 23647
rect 44499 23613 44511 23647
rect 44726 23644 44732 23656
rect 44687 23616 44732 23644
rect 44453 23607 44511 23613
rect 32490 23576 32496 23588
rect 32232 23548 32496 23576
rect 32490 23536 32496 23548
rect 32548 23536 32554 23588
rect 44468 23576 44496 23607
rect 44726 23604 44732 23616
rect 44784 23604 44790 23656
rect 46382 23604 46388 23656
rect 46440 23644 46446 23656
rect 46753 23647 46811 23653
rect 46753 23644 46765 23647
rect 46440 23616 46765 23644
rect 46440 23604 46446 23616
rect 46753 23613 46765 23616
rect 46799 23613 46811 23647
rect 46753 23607 46811 23613
rect 46842 23576 46848 23588
rect 44468 23548 46848 23576
rect 46842 23536 46848 23548
rect 46900 23536 46906 23588
rect 10502 23468 10508 23520
rect 10560 23508 10566 23520
rect 12345 23511 12403 23517
rect 12345 23508 12357 23511
rect 10560 23480 12357 23508
rect 10560 23468 10566 23480
rect 12345 23477 12357 23480
rect 12391 23477 12403 23511
rect 13446 23508 13452 23520
rect 13407 23480 13452 23508
rect 12345 23471 12403 23477
rect 13446 23468 13452 23480
rect 13504 23468 13510 23520
rect 18785 23511 18843 23517
rect 18785 23477 18797 23511
rect 18831 23508 18843 23511
rect 19334 23508 19340 23520
rect 18831 23480 19340 23508
rect 18831 23477 18843 23480
rect 18785 23471 18843 23477
rect 19334 23468 19340 23480
rect 19392 23468 19398 23520
rect 20162 23508 20168 23520
rect 20123 23480 20168 23508
rect 20162 23468 20168 23480
rect 20220 23468 20226 23520
rect 23014 23508 23020 23520
rect 22975 23480 23020 23508
rect 23014 23468 23020 23480
rect 23072 23468 23078 23520
rect 23566 23508 23572 23520
rect 23527 23480 23572 23508
rect 23566 23468 23572 23480
rect 23624 23468 23630 23520
rect 31573 23511 31631 23517
rect 31573 23477 31585 23511
rect 31619 23508 31631 23511
rect 32030 23508 32036 23520
rect 31619 23480 32036 23508
rect 31619 23477 31631 23480
rect 31573 23471 31631 23477
rect 32030 23468 32036 23480
rect 32088 23468 32094 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 8478 23264 8484 23316
rect 8536 23304 8542 23316
rect 9033 23307 9091 23313
rect 9033 23304 9045 23307
rect 8536 23276 9045 23304
rect 8536 23264 8542 23276
rect 9033 23273 9045 23276
rect 9079 23273 9091 23307
rect 9033 23267 9091 23273
rect 9585 23307 9643 23313
rect 9585 23273 9597 23307
rect 9631 23304 9643 23307
rect 9950 23304 9956 23316
rect 9631 23276 9956 23304
rect 9631 23273 9643 23276
rect 9585 23267 9643 23273
rect 9950 23264 9956 23276
rect 10008 23264 10014 23316
rect 10226 23264 10232 23316
rect 10284 23304 10290 23316
rect 10321 23307 10379 23313
rect 10321 23304 10333 23307
rect 10284 23276 10333 23304
rect 10284 23264 10290 23276
rect 10321 23273 10333 23276
rect 10367 23273 10379 23307
rect 10502 23304 10508 23316
rect 10463 23276 10508 23304
rect 10321 23267 10379 23273
rect 10502 23264 10508 23276
rect 10560 23264 10566 23316
rect 11238 23264 11244 23316
rect 11296 23304 11302 23316
rect 11609 23307 11667 23313
rect 11609 23304 11621 23307
rect 11296 23276 11621 23304
rect 11296 23264 11302 23276
rect 11609 23273 11621 23276
rect 11655 23273 11667 23307
rect 14550 23304 14556 23316
rect 14511 23276 14556 23304
rect 11609 23267 11667 23273
rect 14550 23264 14556 23276
rect 14608 23264 14614 23316
rect 18230 23304 18236 23316
rect 18191 23276 18236 23304
rect 18230 23264 18236 23276
rect 18288 23264 18294 23316
rect 20254 23264 20260 23316
rect 20312 23304 20318 23316
rect 47578 23304 47584 23316
rect 20312 23276 47584 23304
rect 20312 23264 20318 23276
rect 47578 23264 47584 23276
rect 47636 23264 47642 23316
rect 10520 23168 10548 23264
rect 10686 23196 10692 23248
rect 10744 23236 10750 23248
rect 14737 23239 14795 23245
rect 14737 23236 14749 23239
rect 10744 23208 14749 23236
rect 10744 23196 10750 23208
rect 14737 23205 14749 23208
rect 14783 23205 14795 23239
rect 15838 23236 15844 23248
rect 14737 23199 14795 23205
rect 15488 23208 15844 23236
rect 9508 23140 10548 23168
rect 9214 23103 9272 23109
rect 9214 23069 9226 23103
rect 9260 23100 9272 23103
rect 9508 23100 9536 23140
rect 10594 23128 10600 23180
rect 10652 23168 10658 23180
rect 15488 23177 15516 23208
rect 15838 23196 15844 23208
rect 15896 23196 15902 23248
rect 33505 23239 33563 23245
rect 33505 23236 33517 23239
rect 33060 23208 33517 23236
rect 13357 23171 13415 23177
rect 13357 23168 13369 23171
rect 10652 23140 13369 23168
rect 10652 23128 10658 23140
rect 13357 23137 13369 23140
rect 13403 23137 13415 23171
rect 13357 23131 13415 23137
rect 15473 23171 15531 23177
rect 15473 23137 15485 23171
rect 15519 23137 15531 23171
rect 15746 23168 15752 23180
rect 15707 23140 15752 23168
rect 15473 23131 15531 23137
rect 15746 23128 15752 23140
rect 15804 23128 15810 23180
rect 19245 23171 19303 23177
rect 19245 23137 19257 23171
rect 19291 23168 19303 23171
rect 19426 23168 19432 23180
rect 19291 23140 19432 23168
rect 19291 23137 19303 23140
rect 19245 23131 19303 23137
rect 19426 23128 19432 23140
rect 19484 23128 19490 23180
rect 22281 23171 22339 23177
rect 22281 23137 22293 23171
rect 22327 23168 22339 23171
rect 23566 23168 23572 23180
rect 22327 23140 23572 23168
rect 22327 23137 22339 23140
rect 22281 23131 22339 23137
rect 23566 23128 23572 23140
rect 23624 23128 23630 23180
rect 23753 23171 23811 23177
rect 23753 23137 23765 23171
rect 23799 23168 23811 23171
rect 24118 23168 24124 23180
rect 23799 23140 24124 23168
rect 23799 23137 23811 23140
rect 23753 23131 23811 23137
rect 24118 23128 24124 23140
rect 24176 23128 24182 23180
rect 30282 23128 30288 23180
rect 30340 23168 30346 23180
rect 31297 23171 31355 23177
rect 31297 23168 31309 23171
rect 30340 23140 31309 23168
rect 30340 23128 30346 23140
rect 31297 23137 31309 23140
rect 31343 23137 31355 23171
rect 31754 23168 31760 23180
rect 31715 23140 31760 23168
rect 31297 23131 31355 23137
rect 31754 23128 31760 23140
rect 31812 23128 31818 23180
rect 32030 23168 32036 23180
rect 31991 23140 32036 23168
rect 32030 23128 32036 23140
rect 32088 23128 32094 23180
rect 32490 23128 32496 23180
rect 32548 23168 32554 23180
rect 33060 23168 33088 23208
rect 33505 23205 33517 23208
rect 33551 23205 33563 23239
rect 33505 23199 33563 23205
rect 41506 23168 41512 23180
rect 32548 23140 33088 23168
rect 33336 23140 41512 23168
rect 32548 23128 32554 23140
rect 9260 23072 9536 23100
rect 9677 23103 9735 23109
rect 9260 23069 9272 23072
rect 9214 23063 9272 23069
rect 9677 23069 9689 23103
rect 9723 23100 9735 23103
rect 9766 23100 9772 23112
rect 9723 23072 9772 23100
rect 9723 23069 9735 23072
rect 9677 23063 9735 23069
rect 9766 23060 9772 23072
rect 9824 23060 9830 23112
rect 11054 23060 11060 23112
rect 11112 23100 11118 23112
rect 11517 23103 11575 23109
rect 11517 23100 11529 23103
rect 11112 23072 11529 23100
rect 11112 23060 11118 23072
rect 11517 23069 11529 23072
rect 11563 23069 11575 23103
rect 11517 23063 11575 23069
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23100 15439 23103
rect 15654 23100 15660 23112
rect 15427 23072 15660 23100
rect 15427 23069 15439 23072
rect 15381 23063 15439 23069
rect 15654 23060 15660 23072
rect 15712 23100 15718 23112
rect 16114 23100 16120 23112
rect 15712 23072 16120 23100
rect 15712 23060 15718 23072
rect 16114 23060 16120 23072
rect 16172 23060 16178 23112
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23100 18107 23103
rect 22005 23103 22063 23109
rect 18095 23072 19288 23100
rect 18095 23069 18107 23072
rect 18049 23063 18107 23069
rect 9950 22992 9956 23044
rect 10008 23032 10014 23044
rect 10137 23035 10195 23041
rect 10137 23032 10149 23035
rect 10008 23004 10149 23032
rect 10008 22992 10014 23004
rect 10137 23001 10149 23004
rect 10183 23001 10195 23035
rect 10137 22995 10195 23001
rect 12986 22992 12992 23044
rect 13044 23032 13050 23044
rect 13081 23035 13139 23041
rect 13081 23032 13093 23035
rect 13044 23004 13093 23032
rect 13044 22992 13050 23004
rect 13081 23001 13093 23004
rect 13127 23001 13139 23035
rect 13081 22995 13139 23001
rect 14369 23035 14427 23041
rect 14369 23001 14381 23035
rect 14415 23032 14427 23035
rect 15286 23032 15292 23044
rect 14415 23004 15292 23032
rect 14415 23001 14427 23004
rect 14369 22995 14427 23001
rect 15286 22992 15292 23004
rect 15344 22992 15350 23044
rect 9217 22967 9275 22973
rect 9217 22933 9229 22967
rect 9263 22964 9275 22967
rect 10042 22964 10048 22976
rect 9263 22936 10048 22964
rect 9263 22933 9275 22936
rect 9217 22927 9275 22933
rect 10042 22924 10048 22936
rect 10100 22924 10106 22976
rect 10318 22924 10324 22976
rect 10376 22973 10382 22976
rect 10376 22967 10395 22973
rect 10383 22933 10395 22967
rect 10376 22927 10395 22933
rect 14579 22967 14637 22973
rect 14579 22933 14591 22967
rect 14625 22964 14637 22967
rect 15194 22964 15200 22976
rect 14625 22936 15200 22964
rect 14625 22933 14637 22936
rect 14579 22927 14637 22933
rect 10376 22924 10382 22927
rect 15194 22924 15200 22936
rect 15252 22964 15258 22976
rect 15378 22964 15384 22976
rect 15252 22936 15384 22964
rect 15252 22924 15258 22936
rect 15378 22924 15384 22936
rect 15436 22924 15442 22976
rect 19260 22964 19288 23072
rect 22005 23069 22017 23103
rect 22051 23069 22063 23103
rect 22005 23063 22063 23069
rect 19426 23032 19432 23044
rect 19387 23004 19432 23032
rect 19426 22992 19432 23004
rect 19484 22992 19490 23044
rect 21085 23035 21143 23041
rect 21085 23001 21097 23035
rect 21131 23032 21143 23035
rect 21174 23032 21180 23044
rect 21131 23004 21180 23032
rect 21131 23001 21143 23004
rect 21085 22995 21143 23001
rect 21174 22992 21180 23004
rect 21232 22992 21238 23044
rect 22020 23032 22048 23063
rect 28534 23060 28540 23112
rect 28592 23100 28598 23112
rect 29549 23103 29607 23109
rect 29549 23100 29561 23103
rect 28592 23072 29561 23100
rect 28592 23060 28598 23072
rect 29549 23069 29561 23072
rect 29595 23069 29607 23103
rect 31478 23100 31484 23112
rect 30958 23072 31484 23100
rect 29549 23063 29607 23069
rect 31478 23060 31484 23072
rect 31536 23060 31542 23112
rect 22278 23032 22284 23044
rect 22020 23004 22284 23032
rect 22278 22992 22284 23004
rect 22336 22992 22342 23044
rect 23014 22992 23020 23044
rect 23072 22992 23078 23044
rect 29822 23032 29828 23044
rect 23682 23004 23888 23032
rect 29783 23004 29828 23032
rect 19978 22964 19984 22976
rect 19260 22936 19984 22964
rect 19978 22924 19984 22936
rect 20036 22964 20042 22976
rect 23682 22964 23710 23004
rect 20036 22936 23710 22964
rect 23860 22964 23888 23004
rect 29822 22992 29828 23004
rect 29880 22992 29886 23044
rect 31128 23004 31754 23032
rect 31128 22964 31156 23004
rect 23860 22936 31156 22964
rect 31726 22964 31754 23004
rect 32490 22992 32496 23044
rect 32548 22992 32554 23044
rect 33336 22964 33364 23140
rect 41506 23128 41512 23140
rect 41564 23128 41570 23180
rect 41782 23168 41788 23180
rect 41743 23140 41788 23168
rect 41782 23128 41788 23140
rect 41840 23128 41846 23180
rect 46290 23168 46296 23180
rect 46251 23140 46296 23168
rect 46290 23128 46296 23140
rect 46348 23128 46354 23180
rect 46750 23168 46756 23180
rect 46711 23140 46756 23168
rect 46750 23128 46756 23140
rect 46808 23128 46814 23180
rect 33410 23060 33416 23112
rect 33468 23100 33474 23112
rect 33965 23103 34023 23109
rect 33965 23100 33977 23103
rect 33468 23072 33977 23100
rect 33468 23060 33474 23072
rect 33965 23069 33977 23072
rect 34011 23100 34023 23103
rect 39758 23100 39764 23112
rect 34011 23072 39764 23100
rect 34011 23069 34023 23072
rect 33965 23063 34023 23069
rect 39758 23060 39764 23072
rect 39816 23060 39822 23112
rect 39942 23100 39948 23112
rect 39903 23072 39948 23100
rect 39942 23060 39948 23072
rect 40000 23060 40006 23112
rect 45833 23103 45891 23109
rect 45833 23069 45845 23103
rect 45879 23100 45891 23103
rect 46014 23100 46020 23112
rect 45879 23072 46020 23100
rect 45879 23069 45891 23072
rect 45833 23063 45891 23069
rect 46014 23060 46020 23072
rect 46072 23060 46078 23112
rect 40126 23032 40132 23044
rect 40087 23004 40132 23032
rect 40126 22992 40132 23004
rect 40184 22992 40190 23044
rect 46477 23035 46535 23041
rect 46477 23001 46489 23035
rect 46523 23032 46535 23035
rect 47670 23032 47676 23044
rect 46523 23004 47676 23032
rect 46523 23001 46535 23004
rect 46477 22995 46535 23001
rect 47670 22992 47676 23004
rect 47728 22992 47734 23044
rect 31726 22936 33364 22964
rect 20036 22924 20042 22936
rect 33870 22924 33876 22976
rect 33928 22964 33934 22976
rect 34057 22967 34115 22973
rect 34057 22964 34069 22967
rect 33928 22936 34069 22964
rect 33928 22924 33934 22936
rect 34057 22933 34069 22936
rect 34103 22933 34115 22967
rect 34057 22927 34115 22933
rect 42794 22924 42800 22976
rect 42852 22964 42858 22976
rect 45649 22967 45707 22973
rect 45649 22964 45661 22967
rect 42852 22936 45661 22964
rect 42852 22924 42858 22936
rect 45649 22933 45661 22936
rect 45695 22933 45707 22967
rect 45649 22927 45707 22933
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 9766 22760 9772 22772
rect 9324 22732 9772 22760
rect 9324 22701 9352 22732
rect 9766 22720 9772 22732
rect 9824 22760 9830 22772
rect 10597 22763 10655 22769
rect 10597 22760 10609 22763
rect 9824 22732 10609 22760
rect 9824 22720 9830 22732
rect 10597 22729 10609 22732
rect 10643 22729 10655 22763
rect 12710 22760 12716 22772
rect 12671 22732 12716 22760
rect 10597 22723 10655 22729
rect 12710 22720 12716 22732
rect 12768 22760 12774 22772
rect 13354 22760 13360 22772
rect 12768 22732 13360 22760
rect 12768 22720 12774 22732
rect 13354 22720 13360 22732
rect 13412 22720 13418 22772
rect 15746 22760 15752 22772
rect 14384 22732 15752 22760
rect 9309 22695 9367 22701
rect 9309 22661 9321 22695
rect 9355 22661 9367 22695
rect 9309 22655 9367 22661
rect 9674 22652 9680 22704
rect 9732 22692 9738 22704
rect 10226 22692 10232 22704
rect 9732 22664 10232 22692
rect 9732 22652 9738 22664
rect 10226 22652 10232 22664
rect 10284 22652 10290 22704
rect 10445 22695 10503 22701
rect 10445 22661 10457 22695
rect 10491 22692 10503 22695
rect 10686 22692 10692 22704
rect 10491 22664 10692 22692
rect 10491 22661 10503 22664
rect 10445 22655 10503 22661
rect 10686 22652 10692 22664
rect 10744 22652 10750 22704
rect 14384 22701 14412 22732
rect 15746 22720 15752 22732
rect 15804 22720 15810 22772
rect 22465 22763 22523 22769
rect 22465 22729 22477 22763
rect 22511 22760 22523 22763
rect 22922 22760 22928 22772
rect 22511 22732 22928 22760
rect 22511 22729 22523 22732
rect 22465 22723 22523 22729
rect 22922 22720 22928 22732
rect 22980 22720 22986 22772
rect 24118 22760 24124 22772
rect 23032 22732 24124 22760
rect 14369 22695 14427 22701
rect 14369 22661 14381 22695
rect 14415 22661 14427 22695
rect 14369 22655 14427 22661
rect 15378 22652 15384 22704
rect 15436 22652 15442 22704
rect 23032 22701 23060 22732
rect 24118 22720 24124 22732
rect 24176 22760 24182 22772
rect 28534 22760 28540 22772
rect 24176 22732 25176 22760
rect 28495 22732 28540 22760
rect 24176 22720 24182 22732
rect 17681 22695 17739 22701
rect 17681 22661 17693 22695
rect 17727 22692 17739 22695
rect 22281 22695 22339 22701
rect 17727 22664 22094 22692
rect 17727 22661 17739 22664
rect 17681 22655 17739 22661
rect 11885 22627 11943 22633
rect 11885 22593 11897 22627
rect 11931 22624 11943 22627
rect 12529 22627 12587 22633
rect 11931 22596 12434 22624
rect 11931 22593 11943 22596
rect 11885 22587 11943 22593
rect 9490 22448 9496 22500
rect 9548 22488 9554 22500
rect 9585 22491 9643 22497
rect 9585 22488 9597 22491
rect 9548 22460 9597 22488
rect 9548 22448 9554 22460
rect 9585 22457 9597 22460
rect 9631 22457 9643 22491
rect 9585 22451 9643 22457
rect 9766 22420 9772 22432
rect 9727 22392 9772 22420
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 9858 22380 9864 22432
rect 9916 22420 9922 22432
rect 10318 22420 10324 22432
rect 9916 22392 10324 22420
rect 9916 22380 9922 22392
rect 10318 22380 10324 22392
rect 10376 22420 10382 22432
rect 10413 22423 10471 22429
rect 10413 22420 10425 22423
rect 10376 22392 10425 22420
rect 10376 22380 10382 22392
rect 10413 22389 10425 22392
rect 10459 22389 10471 22423
rect 10413 22383 10471 22389
rect 11882 22380 11888 22432
rect 11940 22420 11946 22432
rect 11977 22423 12035 22429
rect 11977 22420 11989 22423
rect 11940 22392 11989 22420
rect 11940 22380 11946 22392
rect 11977 22389 11989 22392
rect 12023 22389 12035 22423
rect 12406 22420 12434 22596
rect 12529 22593 12541 22627
rect 12575 22593 12587 22627
rect 12529 22587 12587 22593
rect 13357 22627 13415 22633
rect 13357 22593 13369 22627
rect 13403 22624 13415 22627
rect 13403 22596 13952 22624
rect 13403 22593 13415 22596
rect 13357 22587 13415 22593
rect 12544 22556 12572 22587
rect 13446 22556 13452 22568
rect 12544 22528 13452 22556
rect 13446 22516 13452 22528
rect 13504 22556 13510 22568
rect 13541 22559 13599 22565
rect 13541 22556 13553 22559
rect 13504 22528 13553 22556
rect 13504 22516 13510 22528
rect 13541 22525 13553 22528
rect 13587 22525 13599 22559
rect 13541 22519 13599 22525
rect 13924 22488 13952 22596
rect 16666 22584 16672 22636
rect 16724 22624 16730 22636
rect 16761 22627 16819 22633
rect 16761 22624 16773 22627
rect 16724 22596 16773 22624
rect 16724 22584 16730 22596
rect 16761 22593 16773 22596
rect 16807 22624 16819 22627
rect 18230 22624 18236 22636
rect 16807 22596 18236 22624
rect 16807 22593 16819 22596
rect 16761 22587 16819 22593
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22593 18475 22627
rect 18782 22624 18788 22636
rect 18743 22596 18788 22624
rect 18417 22587 18475 22593
rect 14090 22556 14096 22568
rect 14051 22528 14096 22556
rect 14090 22516 14096 22528
rect 14148 22516 14154 22568
rect 17678 22556 17684 22568
rect 14200 22528 17684 22556
rect 14200 22488 14228 22528
rect 17678 22516 17684 22528
rect 17736 22516 17742 22568
rect 18432 22556 18460 22587
rect 18782 22584 18788 22596
rect 18840 22584 18846 22636
rect 19613 22627 19671 22633
rect 19613 22593 19625 22627
rect 19659 22624 19671 22627
rect 19978 22624 19984 22636
rect 19659 22596 19984 22624
rect 19659 22593 19671 22596
rect 19613 22587 19671 22593
rect 19628 22556 19656 22587
rect 19978 22584 19984 22596
rect 20036 22584 20042 22636
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22624 20223 22627
rect 20254 22624 20260 22636
rect 20211 22596 20260 22624
rect 20211 22593 20223 22596
rect 20165 22587 20223 22593
rect 20254 22584 20260 22596
rect 20312 22584 20318 22636
rect 20898 22624 20904 22636
rect 20859 22596 20904 22624
rect 20898 22584 20904 22596
rect 20956 22584 20962 22636
rect 22066 22624 22094 22664
rect 22281 22661 22293 22695
rect 22327 22692 22339 22695
rect 23017 22695 23075 22701
rect 23017 22692 23029 22695
rect 22327 22664 23029 22692
rect 22327 22661 22339 22664
rect 22281 22655 22339 22661
rect 23017 22661 23029 22664
rect 23063 22661 23075 22695
rect 23233 22695 23291 22701
rect 23233 22692 23245 22695
rect 23017 22655 23075 22661
rect 23216 22661 23245 22692
rect 23279 22692 23291 22695
rect 25148 22692 25176 22732
rect 28534 22720 28540 22732
rect 28592 22720 28598 22772
rect 30742 22760 30748 22772
rect 30703 22732 30748 22760
rect 30742 22720 30748 22732
rect 30800 22720 30806 22772
rect 30929 22763 30987 22769
rect 30929 22729 30941 22763
rect 30975 22760 30987 22763
rect 31110 22760 31116 22772
rect 30975 22732 31116 22760
rect 30975 22729 30987 22732
rect 30929 22723 30987 22729
rect 31110 22720 31116 22732
rect 31168 22720 31174 22772
rect 31478 22760 31484 22772
rect 31439 22732 31484 22760
rect 31478 22720 31484 22732
rect 31536 22720 31542 22772
rect 32217 22763 32275 22769
rect 32217 22729 32229 22763
rect 32263 22760 32275 22763
rect 32490 22760 32496 22772
rect 32263 22732 32496 22760
rect 32263 22729 32275 22732
rect 32217 22723 32275 22729
rect 32490 22720 32496 22732
rect 32548 22720 32554 22772
rect 33042 22760 33048 22772
rect 33003 22732 33048 22760
rect 33042 22720 33048 22732
rect 33100 22720 33106 22772
rect 40126 22760 40132 22772
rect 40087 22732 40132 22760
rect 40126 22720 40132 22732
rect 40184 22720 40190 22772
rect 45189 22763 45247 22769
rect 45189 22729 45201 22763
rect 45235 22760 45247 22763
rect 45830 22760 45836 22772
rect 45235 22732 45836 22760
rect 45235 22729 45247 22732
rect 45189 22723 45247 22729
rect 45830 22720 45836 22732
rect 45888 22720 45894 22772
rect 47670 22760 47676 22772
rect 47631 22732 47676 22760
rect 47670 22720 47676 22732
rect 47728 22720 47734 22772
rect 39942 22692 39948 22704
rect 23279 22664 25084 22692
rect 25148 22664 39948 22692
rect 23279 22661 23291 22664
rect 23216 22655 23291 22661
rect 22370 22624 22376 22636
rect 22066 22596 22376 22624
rect 22370 22584 22376 22596
rect 22428 22584 22434 22636
rect 22557 22627 22615 22633
rect 22557 22593 22569 22627
rect 22603 22624 22615 22627
rect 23216 22624 23244 22655
rect 23842 22624 23848 22636
rect 22603 22596 23244 22624
rect 23803 22596 23848 22624
rect 22603 22593 22615 22596
rect 22557 22587 22615 22593
rect 20806 22556 20812 22568
rect 18432 22528 19656 22556
rect 20767 22528 20812 22556
rect 20806 22516 20812 22528
rect 20864 22556 20870 22568
rect 22572 22556 22600 22587
rect 23842 22584 23848 22596
rect 23900 22584 23906 22636
rect 23934 22584 23940 22636
rect 23992 22624 23998 22636
rect 25056 22633 25084 22664
rect 39942 22652 39948 22664
rect 40000 22652 40006 22704
rect 41506 22692 41512 22704
rect 41467 22664 41512 22692
rect 41506 22652 41512 22664
rect 41564 22652 41570 22704
rect 45020 22664 45876 22692
rect 24029 22627 24087 22633
rect 24029 22624 24041 22627
rect 23992 22596 24041 22624
rect 23992 22584 23998 22596
rect 24029 22593 24041 22596
rect 24075 22593 24087 22627
rect 24029 22587 24087 22593
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22593 24271 22627
rect 24213 22587 24271 22593
rect 25041 22627 25099 22633
rect 25041 22593 25053 22627
rect 25087 22593 25099 22627
rect 25041 22587 25099 22593
rect 25869 22627 25927 22633
rect 25869 22593 25881 22627
rect 25915 22624 25927 22627
rect 25958 22624 25964 22636
rect 25915 22596 25964 22624
rect 25915 22593 25927 22596
rect 25869 22587 25927 22593
rect 23474 22556 23480 22568
rect 20864 22528 22600 22556
rect 22940 22528 23480 22556
rect 20864 22516 20870 22528
rect 15930 22488 15936 22500
rect 13924 22460 14228 22488
rect 15396 22460 15936 22488
rect 15396 22420 15424 22460
rect 15930 22448 15936 22460
rect 15988 22448 15994 22500
rect 17862 22488 17868 22500
rect 17823 22460 17868 22488
rect 17862 22448 17868 22460
rect 17920 22448 17926 22500
rect 22830 22488 22836 22500
rect 22066 22460 22836 22488
rect 12406 22392 15424 22420
rect 15841 22423 15899 22429
rect 11977 22383 12035 22389
rect 15841 22389 15853 22423
rect 15887 22420 15899 22423
rect 16114 22420 16120 22432
rect 15887 22392 16120 22420
rect 15887 22389 15899 22392
rect 15841 22383 15899 22389
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 16850 22420 16856 22432
rect 16811 22392 16856 22420
rect 16850 22380 16856 22392
rect 16908 22380 16914 22432
rect 20806 22380 20812 22432
rect 20864 22420 20870 22432
rect 21082 22420 21088 22432
rect 20864 22392 21088 22420
rect 20864 22380 20870 22392
rect 21082 22380 21088 22392
rect 21140 22380 21146 22432
rect 21266 22420 21272 22432
rect 21227 22392 21272 22420
rect 21266 22380 21272 22392
rect 21324 22380 21330 22432
rect 21818 22380 21824 22432
rect 21876 22420 21882 22432
rect 22066 22420 22094 22460
rect 22830 22448 22836 22460
rect 22888 22448 22894 22500
rect 21876 22392 22094 22420
rect 22281 22423 22339 22429
rect 21876 22380 21882 22392
rect 22281 22389 22293 22423
rect 22327 22420 22339 22423
rect 22940 22420 22968 22528
rect 23474 22516 23480 22528
rect 23532 22516 23538 22568
rect 23382 22488 23388 22500
rect 23343 22460 23388 22488
rect 23382 22448 23388 22460
rect 23440 22448 23446 22500
rect 22327 22392 22968 22420
rect 22327 22389 22339 22392
rect 22281 22383 22339 22389
rect 23014 22380 23020 22432
rect 23072 22420 23078 22432
rect 23201 22423 23259 22429
rect 23201 22420 23213 22423
rect 23072 22392 23213 22420
rect 23072 22380 23078 22392
rect 23201 22389 23213 22392
rect 23247 22420 23259 22423
rect 24228 22420 24256 22587
rect 25958 22584 25964 22596
rect 26016 22584 26022 22636
rect 28534 22624 28540 22636
rect 28447 22596 28540 22624
rect 28534 22584 28540 22596
rect 28592 22624 28598 22636
rect 28718 22624 28724 22636
rect 28592 22596 28724 22624
rect 28592 22584 28598 22596
rect 28718 22584 28724 22596
rect 28776 22584 28782 22636
rect 29270 22624 29276 22636
rect 29231 22596 29276 22624
rect 29270 22584 29276 22596
rect 29328 22624 29334 22636
rect 30282 22624 30288 22636
rect 29328 22596 30288 22624
rect 29328 22584 29334 22596
rect 30282 22584 30288 22596
rect 30340 22624 30346 22636
rect 30377 22627 30435 22633
rect 30377 22624 30389 22627
rect 30340 22596 30389 22624
rect 30340 22584 30346 22596
rect 30377 22593 30389 22596
rect 30423 22593 30435 22627
rect 30558 22624 30564 22636
rect 30519 22596 30564 22624
rect 30377 22587 30435 22593
rect 30558 22584 30564 22596
rect 30616 22584 30622 22636
rect 30653 22627 30711 22633
rect 30653 22593 30665 22627
rect 30699 22593 30711 22627
rect 31386 22624 31392 22636
rect 31347 22596 31392 22624
rect 30653 22587 30711 22593
rect 24397 22559 24455 22565
rect 24397 22525 24409 22559
rect 24443 22556 24455 22559
rect 24857 22559 24915 22565
rect 24857 22556 24869 22559
rect 24443 22528 24869 22556
rect 24443 22525 24455 22528
rect 24397 22519 24455 22525
rect 24857 22525 24869 22528
rect 24903 22525 24915 22559
rect 24857 22519 24915 22525
rect 29365 22559 29423 22565
rect 29365 22525 29377 22559
rect 29411 22525 29423 22559
rect 29365 22519 29423 22525
rect 29641 22559 29699 22565
rect 29641 22525 29653 22559
rect 29687 22556 29699 22559
rect 29822 22556 29828 22568
rect 29687 22528 29828 22556
rect 29687 22525 29699 22528
rect 29641 22519 29699 22525
rect 29380 22488 29408 22519
rect 29822 22516 29828 22528
rect 29880 22516 29886 22568
rect 30668 22556 30696 22587
rect 31386 22584 31392 22596
rect 31444 22624 31450 22636
rect 32125 22627 32183 22633
rect 32125 22624 32137 22627
rect 31444 22596 32137 22624
rect 31444 22584 31450 22596
rect 32125 22593 32137 22596
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 32953 22627 33011 22633
rect 32953 22593 32965 22627
rect 32999 22624 33011 22627
rect 33410 22624 33416 22636
rect 32999 22596 33416 22624
rect 32999 22593 33011 22596
rect 32953 22587 33011 22593
rect 33410 22584 33416 22596
rect 33468 22584 33474 22636
rect 39758 22584 39764 22636
rect 39816 22624 39822 22636
rect 40037 22627 40095 22633
rect 40037 22624 40049 22627
rect 39816 22596 40049 22624
rect 39816 22584 39822 22596
rect 40037 22593 40049 22596
rect 40083 22593 40095 22627
rect 41524 22624 41552 22652
rect 45020 22633 45048 22664
rect 45848 22636 45876 22664
rect 42429 22627 42487 22633
rect 42429 22624 42441 22627
rect 41524 22596 42441 22624
rect 40037 22587 40095 22593
rect 42429 22593 42441 22596
rect 42475 22593 42487 22627
rect 42429 22587 42487 22593
rect 45005 22627 45063 22633
rect 45005 22593 45017 22627
rect 45051 22593 45063 22627
rect 45005 22587 45063 22593
rect 45189 22627 45247 22633
rect 45189 22593 45201 22627
rect 45235 22624 45247 22627
rect 45235 22596 45692 22624
rect 45235 22593 45247 22596
rect 45189 22587 45247 22593
rect 31110 22556 31116 22568
rect 30668 22528 31116 22556
rect 31110 22516 31116 22528
rect 31168 22556 31174 22568
rect 33689 22559 33747 22565
rect 33689 22556 33701 22559
rect 31168 22528 33701 22556
rect 31168 22516 31174 22528
rect 33689 22525 33701 22528
rect 33735 22525 33747 22559
rect 33870 22556 33876 22568
rect 33831 22528 33876 22556
rect 33689 22519 33747 22525
rect 33870 22516 33876 22528
rect 33928 22516 33934 22568
rect 35529 22559 35587 22565
rect 35529 22525 35541 22559
rect 35575 22556 35587 22559
rect 40052 22556 40080 22587
rect 41598 22556 41604 22568
rect 35575 22528 35894 22556
rect 40052 22528 41604 22556
rect 35575 22525 35587 22528
rect 35529 22519 35587 22525
rect 30282 22488 30288 22500
rect 29380 22460 30288 22488
rect 30282 22448 30288 22460
rect 30340 22448 30346 22500
rect 35866 22488 35894 22528
rect 41598 22516 41604 22528
rect 41656 22516 41662 22568
rect 45664 22565 45692 22596
rect 45830 22584 45836 22636
rect 45888 22624 45894 22636
rect 46385 22627 46443 22633
rect 46385 22624 46397 22627
rect 45888 22596 46397 22624
rect 45888 22584 45894 22596
rect 46385 22593 46397 22596
rect 46431 22593 46443 22627
rect 47578 22624 47584 22636
rect 47539 22596 47584 22624
rect 46385 22587 46443 22593
rect 47578 22584 47584 22596
rect 47636 22584 47642 22636
rect 42705 22559 42763 22565
rect 42705 22525 42717 22559
rect 42751 22556 42763 22559
rect 45649 22559 45707 22565
rect 42751 22528 45554 22556
rect 42751 22525 42763 22528
rect 42705 22519 42763 22525
rect 43530 22488 43536 22500
rect 35866 22460 43536 22488
rect 43530 22448 43536 22460
rect 43588 22448 43594 22500
rect 25222 22420 25228 22432
rect 23247 22392 24256 22420
rect 25183 22392 25228 22420
rect 23247 22389 23259 22392
rect 23201 22383 23259 22389
rect 25222 22380 25228 22392
rect 25280 22380 25286 22432
rect 25682 22420 25688 22432
rect 25643 22392 25688 22420
rect 25682 22380 25688 22392
rect 25740 22380 25746 22432
rect 26234 22380 26240 22432
rect 26292 22420 26298 22432
rect 31202 22420 31208 22432
rect 26292 22392 31208 22420
rect 26292 22380 26298 22392
rect 31202 22380 31208 22392
rect 31260 22380 31266 22432
rect 41598 22420 41604 22432
rect 41559 22392 41604 22420
rect 41598 22380 41604 22392
rect 41656 22380 41662 22432
rect 45526 22420 45554 22528
rect 45649 22525 45661 22559
rect 45695 22556 45707 22559
rect 46198 22556 46204 22568
rect 45695 22528 46204 22556
rect 45695 22525 45707 22528
rect 45649 22519 45707 22525
rect 46198 22516 46204 22528
rect 46256 22516 46262 22568
rect 46750 22556 46756 22568
rect 46711 22528 46756 22556
rect 46750 22516 46756 22528
rect 46808 22516 46814 22568
rect 45922 22488 45928 22500
rect 45883 22460 45928 22488
rect 45922 22448 45928 22460
rect 45980 22448 45986 22500
rect 47486 22420 47492 22432
rect 45526 22392 47492 22420
rect 47486 22380 47492 22392
rect 47544 22380 47550 22432
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 9490 22216 9496 22228
rect 9451 22188 9496 22216
rect 9490 22176 9496 22188
rect 9548 22176 9554 22228
rect 14090 22216 14096 22228
rect 14051 22188 14096 22216
rect 14090 22176 14096 22188
rect 14148 22176 14154 22228
rect 20244 22219 20302 22225
rect 20244 22185 20256 22219
rect 20290 22216 20302 22219
rect 21266 22216 21272 22228
rect 20290 22188 21272 22216
rect 20290 22185 20302 22188
rect 20244 22179 20302 22185
rect 21266 22176 21272 22188
rect 21324 22176 21330 22228
rect 22278 22216 22284 22228
rect 22239 22188 22284 22216
rect 22278 22176 22284 22188
rect 22336 22176 22342 22228
rect 22370 22176 22376 22228
rect 22428 22216 22434 22228
rect 26234 22216 26240 22228
rect 22428 22188 26240 22216
rect 22428 22176 22434 22188
rect 26234 22176 26240 22188
rect 26292 22176 26298 22228
rect 26418 22216 26424 22228
rect 26379 22188 26424 22216
rect 26418 22176 26424 22188
rect 26476 22176 26482 22228
rect 30193 22219 30251 22225
rect 30193 22216 30205 22219
rect 29472 22188 30205 22216
rect 11716 22120 12020 22148
rect 9766 22080 9772 22092
rect 8404 22052 9772 22080
rect 8404 22021 8432 22052
rect 9766 22040 9772 22052
rect 9824 22040 9830 22092
rect 10042 22040 10048 22092
rect 10100 22080 10106 22092
rect 11716 22080 11744 22120
rect 11882 22080 11888 22092
rect 10100 22052 11744 22080
rect 11843 22052 11888 22080
rect 10100 22040 10106 22052
rect 11882 22040 11888 22052
rect 11940 22040 11946 22092
rect 11992 22080 12020 22120
rect 17788 22120 18092 22148
rect 12161 22083 12219 22089
rect 12161 22080 12173 22083
rect 11992 22052 12173 22080
rect 12161 22049 12173 22052
rect 12207 22049 12219 22083
rect 12161 22043 12219 22049
rect 13354 22040 13360 22092
rect 13412 22080 13418 22092
rect 14921 22083 14979 22089
rect 13412 22052 14872 22080
rect 13412 22040 13418 22052
rect 8389 22015 8447 22021
rect 8389 21981 8401 22015
rect 8435 21981 8447 22015
rect 8389 21975 8447 21981
rect 9677 22015 9735 22021
rect 9677 21981 9689 22015
rect 9723 21981 9735 22015
rect 10597 22015 10655 22021
rect 9677 21975 9735 21981
rect 9963 21993 10021 21999
rect 9692 21944 9720 21975
rect 9963 21959 9975 21993
rect 10009 21990 10021 21993
rect 10009 21962 10088 21990
rect 10597 21981 10609 22015
rect 10643 22012 10655 22015
rect 10686 22012 10692 22024
rect 10643 21984 10692 22012
rect 10643 21981 10655 21984
rect 10597 21975 10655 21981
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 11698 22012 11704 22024
rect 11659 21984 11704 22012
rect 11698 21972 11704 21984
rect 11756 21972 11762 22024
rect 13538 21972 13544 22024
rect 13596 22012 13602 22024
rect 14844 22021 14872 22052
rect 14921 22049 14933 22083
rect 14967 22080 14979 22083
rect 15378 22080 15384 22092
rect 14967 22052 15384 22080
rect 14967 22049 14979 22052
rect 14921 22043 14979 22049
rect 15378 22040 15384 22052
rect 15436 22040 15442 22092
rect 17788 22080 17816 22120
rect 17954 22080 17960 22092
rect 15488 22052 17816 22080
rect 17915 22052 17960 22080
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13596 21984 14105 22012
rect 13596 21972 13602 21984
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 14829 22015 14887 22021
rect 14829 21981 14841 22015
rect 14875 21981 14887 22015
rect 14829 21975 14887 21981
rect 10009 21959 10021 21962
rect 9766 21944 9772 21956
rect 9692 21916 9772 21944
rect 9766 21904 9772 21916
rect 9824 21904 9830 21956
rect 9963 21953 10021 21959
rect 10060 21944 10088 21962
rect 10134 21944 10140 21956
rect 10060 21916 10140 21944
rect 10134 21904 10140 21916
rect 10192 21944 10198 21956
rect 10781 21947 10839 21953
rect 10781 21944 10793 21947
rect 10192 21916 10793 21944
rect 10192 21904 10198 21916
rect 10781 21913 10793 21916
rect 10827 21944 10839 21947
rect 11422 21944 11428 21956
rect 10827 21916 11428 21944
rect 10827 21913 10839 21916
rect 10781 21907 10839 21913
rect 11422 21904 11428 21916
rect 11480 21904 11486 21956
rect 13446 21904 13452 21956
rect 13504 21944 13510 21956
rect 15488 21944 15516 22052
rect 17954 22040 17960 22052
rect 18012 22040 18018 22092
rect 18064 22080 18092 22120
rect 23842 22108 23848 22160
rect 23900 22108 23906 22160
rect 20898 22080 20904 22092
rect 18064 22052 19288 22080
rect 19260 22024 19288 22052
rect 19352 22052 20904 22080
rect 16761 22015 16819 22021
rect 16761 21981 16773 22015
rect 16807 21981 16819 22015
rect 19242 22012 19248 22024
rect 19203 21984 19248 22012
rect 16761 21975 16819 21981
rect 13504 21916 15516 21944
rect 13504 21904 13510 21916
rect 8202 21876 8208 21888
rect 8163 21848 8208 21876
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 9861 21879 9919 21885
rect 9861 21845 9873 21879
rect 9907 21876 9919 21879
rect 9950 21876 9956 21888
rect 9907 21848 9956 21876
rect 9907 21845 9919 21848
rect 9861 21839 9919 21845
rect 9950 21836 9956 21848
rect 10008 21876 10014 21888
rect 10594 21876 10600 21888
rect 10008 21848 10600 21876
rect 10008 21836 10014 21848
rect 10594 21836 10600 21848
rect 10652 21836 10658 21888
rect 16776 21876 16804 21975
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 16942 21944 16948 21956
rect 16903 21916 16948 21944
rect 16942 21904 16948 21916
rect 17000 21904 17006 21956
rect 19352 21876 19380 22052
rect 20898 22040 20904 22052
rect 20956 22080 20962 22092
rect 21726 22080 21732 22092
rect 20956 22052 21732 22080
rect 20956 22040 20962 22052
rect 21726 22040 21732 22052
rect 21784 22040 21790 22092
rect 23860 22080 23888 22108
rect 23584 22052 23888 22080
rect 24673 22083 24731 22089
rect 19978 22012 19984 22024
rect 19939 21984 19984 22012
rect 19978 21972 19984 21984
rect 20036 21972 20042 22024
rect 22465 22015 22523 22021
rect 22465 21981 22477 22015
rect 22511 22012 22523 22015
rect 22554 22012 22560 22024
rect 22511 21984 22560 22012
rect 22511 21981 22523 21984
rect 22465 21975 22523 21981
rect 22554 21972 22560 21984
rect 22612 21972 22618 22024
rect 23584 22021 23612 22052
rect 24673 22049 24685 22083
rect 24719 22080 24731 22083
rect 25682 22080 25688 22092
rect 24719 22052 25688 22080
rect 24719 22049 24731 22052
rect 24673 22043 24731 22049
rect 25682 22040 25688 22052
rect 25740 22040 25746 22092
rect 27157 22083 27215 22089
rect 27157 22049 27169 22083
rect 27203 22080 27215 22083
rect 27706 22080 27712 22092
rect 27203 22052 27712 22080
rect 27203 22049 27215 22052
rect 27157 22043 27215 22049
rect 27706 22040 27712 22052
rect 27764 22040 27770 22092
rect 29472 22080 29500 22188
rect 30193 22185 30205 22188
rect 30239 22185 30251 22219
rect 30193 22179 30251 22185
rect 30208 22148 30236 22179
rect 30282 22176 30288 22228
rect 30340 22216 30346 22228
rect 30377 22219 30435 22225
rect 30377 22216 30389 22219
rect 30340 22188 30389 22216
rect 30340 22176 30346 22188
rect 30377 22185 30389 22188
rect 30423 22185 30435 22219
rect 30377 22179 30435 22185
rect 41417 22219 41475 22225
rect 41417 22185 41429 22219
rect 41463 22216 41475 22219
rect 41506 22216 41512 22228
rect 41463 22188 41512 22216
rect 41463 22185 41475 22188
rect 41417 22179 41475 22185
rect 41506 22176 41512 22188
rect 41564 22176 41570 22228
rect 45830 22216 45836 22228
rect 45791 22188 45836 22216
rect 45830 22176 45836 22188
rect 45888 22176 45894 22228
rect 31110 22148 31116 22160
rect 30208 22120 31116 22148
rect 31110 22108 31116 22120
rect 31168 22108 31174 22160
rect 28644 22052 29500 22080
rect 23569 22015 23627 22021
rect 23569 21981 23581 22015
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 23658 21972 23664 22024
rect 23716 22012 23722 22024
rect 23845 22015 23903 22021
rect 23845 22012 23857 22015
rect 23716 21984 23857 22012
rect 23716 21972 23722 21984
rect 23845 21981 23857 21984
rect 23891 21981 23903 22015
rect 26878 22012 26884 22024
rect 26839 21984 26884 22012
rect 23845 21975 23903 21981
rect 26878 21972 26884 21984
rect 26936 21972 26942 22024
rect 28258 21972 28264 22024
rect 28316 21972 28322 22024
rect 20990 21904 20996 21956
rect 21048 21904 21054 21956
rect 24670 21944 24676 21956
rect 23676 21916 24676 21944
rect 16776 21848 19380 21876
rect 19429 21879 19487 21885
rect 19429 21845 19441 21879
rect 19475 21876 19487 21879
rect 20070 21876 20076 21888
rect 19475 21848 20076 21876
rect 19475 21845 19487 21848
rect 19429 21839 19487 21845
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 21818 21836 21824 21888
rect 21876 21876 21882 21888
rect 23290 21876 23296 21888
rect 21876 21848 23296 21876
rect 21876 21836 21882 21848
rect 23290 21836 23296 21848
rect 23348 21836 23354 21888
rect 23676 21885 23704 21916
rect 24670 21904 24676 21916
rect 24728 21904 24734 21956
rect 24854 21904 24860 21956
rect 24912 21944 24918 21956
rect 24949 21947 25007 21953
rect 24949 21944 24961 21947
rect 24912 21916 24961 21944
rect 24912 21904 24918 21916
rect 24949 21913 24961 21916
rect 24995 21913 25007 21947
rect 26234 21944 26240 21956
rect 26174 21916 26240 21944
rect 24949 21907 25007 21913
rect 26234 21904 26240 21916
rect 26292 21904 26298 21956
rect 23667 21879 23725 21885
rect 23667 21845 23679 21879
rect 23713 21845 23725 21879
rect 23667 21839 23725 21845
rect 23753 21879 23811 21885
rect 23753 21845 23765 21879
rect 23799 21876 23811 21879
rect 23934 21876 23940 21888
rect 23799 21848 23940 21876
rect 23799 21845 23811 21848
rect 23753 21839 23811 21845
rect 23934 21836 23940 21848
rect 23992 21836 23998 21888
rect 27338 21836 27344 21888
rect 27396 21876 27402 21888
rect 28644 21885 28672 22052
rect 44726 22040 44732 22092
rect 44784 22080 44790 22092
rect 46477 22083 46535 22089
rect 46477 22080 46489 22083
rect 44784 22052 46489 22080
rect 44784 22040 44790 22052
rect 46477 22049 46489 22052
rect 46523 22049 46535 22083
rect 47762 22080 47768 22092
rect 47723 22052 47768 22080
rect 46477 22043 46535 22049
rect 47762 22040 47768 22052
rect 47820 22040 47826 22092
rect 30742 22012 30748 22024
rect 29932 21984 30748 22012
rect 29932 21888 29960 21984
rect 30742 21972 30748 21984
rect 30800 22012 30806 22024
rect 31113 22015 31171 22021
rect 31113 22012 31125 22015
rect 30800 21984 31125 22012
rect 30800 21972 30806 21984
rect 31113 21981 31125 21984
rect 31159 21981 31171 22015
rect 41230 22012 41236 22024
rect 41191 21984 41236 22012
rect 31113 21975 31171 21981
rect 41230 21972 41236 21984
rect 41288 21972 41294 22024
rect 43901 22015 43959 22021
rect 43901 21981 43913 22015
rect 43947 22012 43959 22015
rect 45554 22012 45560 22024
rect 43947 21984 45560 22012
rect 43947 21981 43959 21984
rect 43901 21975 43959 21981
rect 45554 21972 45560 21984
rect 45612 21972 45618 22024
rect 45830 21972 45836 22024
rect 45888 22012 45894 22024
rect 46290 22012 46296 22024
rect 45888 21984 46296 22012
rect 45888 21972 45894 21984
rect 46290 21972 46296 21984
rect 46348 21972 46354 22024
rect 30009 21947 30067 21953
rect 30009 21913 30021 21947
rect 30055 21944 30067 21947
rect 30558 21944 30564 21956
rect 30055 21916 30564 21944
rect 30055 21913 30067 21916
rect 30009 21907 30067 21913
rect 30558 21904 30564 21916
rect 30616 21944 30622 21956
rect 30837 21947 30895 21953
rect 30837 21944 30849 21947
rect 30616 21916 30849 21944
rect 30616 21904 30622 21916
rect 30837 21913 30849 21916
rect 30883 21944 30895 21947
rect 31938 21944 31944 21956
rect 30883 21916 31944 21944
rect 30883 21913 30895 21916
rect 30837 21907 30895 21913
rect 31938 21904 31944 21916
rect 31996 21904 32002 21956
rect 45465 21947 45523 21953
rect 45465 21913 45477 21947
rect 45511 21913 45523 21947
rect 45465 21907 45523 21913
rect 45649 21947 45707 21953
rect 45649 21913 45661 21947
rect 45695 21944 45707 21947
rect 45695 21916 46336 21944
rect 45695 21913 45707 21916
rect 45649 21907 45707 21913
rect 28629 21879 28687 21885
rect 28629 21876 28641 21879
rect 27396 21848 28641 21876
rect 27396 21836 27402 21848
rect 28629 21845 28641 21848
rect 28675 21845 28687 21879
rect 28629 21839 28687 21845
rect 29914 21836 29920 21888
rect 29972 21876 29978 21888
rect 30209 21879 30267 21885
rect 30209 21876 30221 21879
rect 29972 21848 30221 21876
rect 29972 21836 29978 21848
rect 30209 21845 30221 21848
rect 30255 21845 30267 21879
rect 30209 21839 30267 21845
rect 30374 21836 30380 21888
rect 30432 21876 30438 21888
rect 30935 21879 30993 21885
rect 30935 21876 30947 21879
rect 30432 21848 30947 21876
rect 30432 21836 30438 21848
rect 30935 21845 30947 21848
rect 30981 21845 30993 21879
rect 30935 21839 30993 21845
rect 31021 21879 31079 21885
rect 31021 21845 31033 21879
rect 31067 21876 31079 21879
rect 31110 21876 31116 21888
rect 31067 21848 31116 21876
rect 31067 21845 31079 21848
rect 31021 21839 31079 21845
rect 31110 21836 31116 21848
rect 31168 21836 31174 21888
rect 43990 21876 43996 21888
rect 43951 21848 43996 21876
rect 43990 21836 43996 21848
rect 44048 21836 44054 21888
rect 45480 21876 45508 21907
rect 46308 21888 46336 21916
rect 45922 21876 45928 21888
rect 45480 21848 45928 21876
rect 45922 21836 45928 21848
rect 45980 21836 45986 21888
rect 46290 21836 46296 21888
rect 46348 21836 46354 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 4614 21632 4620 21684
rect 4672 21672 4678 21684
rect 10042 21672 10048 21684
rect 4672 21644 10048 21672
rect 4672 21632 4678 21644
rect 10042 21632 10048 21644
rect 10100 21632 10106 21684
rect 16025 21675 16083 21681
rect 16025 21641 16037 21675
rect 16071 21672 16083 21675
rect 16942 21672 16948 21684
rect 16071 21644 16948 21672
rect 16071 21641 16083 21644
rect 16025 21635 16083 21641
rect 16942 21632 16948 21644
rect 17000 21632 17006 21684
rect 20438 21632 20444 21684
rect 20496 21672 20502 21684
rect 20993 21675 21051 21681
rect 20993 21672 21005 21675
rect 20496 21644 21005 21672
rect 20496 21632 20502 21644
rect 20993 21641 21005 21644
rect 21039 21672 21051 21675
rect 22554 21672 22560 21684
rect 21039 21644 22560 21672
rect 21039 21641 21051 21644
rect 20993 21635 21051 21641
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 23290 21632 23296 21684
rect 23348 21672 23354 21684
rect 24854 21672 24860 21684
rect 23348 21644 23796 21672
rect 24815 21644 24860 21672
rect 23348 21632 23354 21644
rect 8202 21564 8208 21616
rect 8260 21604 8266 21616
rect 9401 21607 9459 21613
rect 9401 21604 9413 21607
rect 8260 21576 9413 21604
rect 8260 21564 8266 21576
rect 9401 21573 9413 21576
rect 9447 21573 9459 21607
rect 9401 21567 9459 21573
rect 10134 21564 10140 21616
rect 10192 21564 10198 21616
rect 16666 21604 16672 21616
rect 15304 21576 16672 21604
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 13173 21539 13231 21545
rect 13173 21536 13185 21539
rect 11931 21508 13185 21536
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 13173 21505 13185 21508
rect 13219 21536 13231 21539
rect 13446 21536 13452 21548
rect 13219 21508 13452 21536
rect 13219 21505 13231 21508
rect 13173 21499 13231 21505
rect 13446 21496 13452 21508
rect 13504 21496 13510 21548
rect 15304 21545 15332 21576
rect 16666 21564 16672 21576
rect 16724 21564 16730 21616
rect 16850 21604 16856 21616
rect 16811 21576 16856 21604
rect 16850 21564 16856 21576
rect 16908 21564 16914 21616
rect 19242 21564 19248 21616
rect 19300 21604 19306 21616
rect 22278 21604 22284 21616
rect 19300 21576 22284 21604
rect 19300 21564 19306 21576
rect 22278 21564 22284 21576
rect 22336 21564 22342 21616
rect 22462 21564 22468 21616
rect 22520 21604 22526 21616
rect 22520 21576 23704 21604
rect 22520 21564 22526 21576
rect 15289 21539 15347 21545
rect 15289 21505 15301 21539
rect 15335 21505 15347 21539
rect 15930 21536 15936 21548
rect 15891 21508 15936 21536
rect 15289 21499 15347 21505
rect 15930 21496 15936 21508
rect 15988 21496 15994 21548
rect 19886 21496 19892 21548
rect 19944 21536 19950 21548
rect 19981 21539 20039 21545
rect 19981 21536 19993 21539
rect 19944 21508 19993 21536
rect 19944 21496 19950 21508
rect 19981 21505 19993 21508
rect 20027 21536 20039 21539
rect 20809 21539 20867 21545
rect 20809 21536 20821 21539
rect 20027 21508 20821 21536
rect 20027 21505 20039 21508
rect 19981 21499 20039 21505
rect 20809 21505 20821 21508
rect 20855 21505 20867 21539
rect 22186 21536 22192 21548
rect 22147 21508 22192 21536
rect 20809 21499 20867 21505
rect 22186 21496 22192 21508
rect 22244 21496 22250 21548
rect 22554 21496 22560 21548
rect 22612 21536 22618 21548
rect 23201 21539 23259 21545
rect 23201 21536 23213 21539
rect 22612 21508 23213 21536
rect 22612 21496 22618 21508
rect 23201 21505 23213 21508
rect 23247 21536 23259 21539
rect 23247 21508 23520 21536
rect 23247 21505 23259 21508
rect 23201 21499 23259 21505
rect 9122 21468 9128 21480
rect 9083 21440 9128 21468
rect 9122 21428 9128 21440
rect 9180 21428 9186 21480
rect 9766 21428 9772 21480
rect 9824 21468 9830 21480
rect 10873 21471 10931 21477
rect 10873 21468 10885 21471
rect 9824 21440 10885 21468
rect 9824 21428 9830 21440
rect 10873 21437 10885 21440
rect 10919 21468 10931 21471
rect 16669 21471 16727 21477
rect 16669 21468 16681 21471
rect 10919 21440 16681 21468
rect 10919 21437 10931 21440
rect 10873 21431 10931 21437
rect 16669 21437 16681 21440
rect 16715 21437 16727 21471
rect 18322 21468 18328 21480
rect 18283 21440 18328 21468
rect 16669 21431 16727 21437
rect 18322 21428 18328 21440
rect 18380 21428 18386 21480
rect 22281 21471 22339 21477
rect 22281 21437 22293 21471
rect 22327 21468 22339 21471
rect 23382 21468 23388 21480
rect 22327 21440 23388 21468
rect 22327 21437 22339 21440
rect 22281 21431 22339 21437
rect 23382 21428 23388 21440
rect 23440 21428 23446 21480
rect 22094 21360 22100 21412
rect 22152 21400 22158 21412
rect 23017 21403 23075 21409
rect 23017 21400 23029 21403
rect 22152 21372 23029 21400
rect 22152 21360 22158 21372
rect 23017 21369 23029 21372
rect 23063 21369 23075 21403
rect 23492 21400 23520 21508
rect 23676 21468 23704 21576
rect 23768 21545 23796 21644
rect 24854 21632 24860 21644
rect 24912 21632 24918 21684
rect 26234 21672 26240 21684
rect 26195 21644 26240 21672
rect 26234 21632 26240 21644
rect 26292 21632 26298 21684
rect 28258 21672 28264 21684
rect 28219 21644 28264 21672
rect 28258 21632 28264 21644
rect 28316 21632 28322 21684
rect 28350 21632 28356 21684
rect 28408 21672 28414 21684
rect 28408 21644 35894 21672
rect 28408 21632 28414 21644
rect 29914 21604 29920 21616
rect 25240 21576 29920 21604
rect 25240 21548 25268 21576
rect 23753 21539 23811 21545
rect 23753 21505 23765 21539
rect 23799 21505 23811 21539
rect 23753 21499 23811 21505
rect 24670 21496 24676 21548
rect 24728 21536 24734 21548
rect 24765 21539 24823 21545
rect 24765 21536 24777 21539
rect 24728 21508 24777 21536
rect 24728 21496 24734 21508
rect 24765 21505 24777 21508
rect 24811 21505 24823 21539
rect 24765 21499 24823 21505
rect 24949 21539 25007 21545
rect 24949 21505 24961 21539
rect 24995 21536 25007 21539
rect 25222 21536 25228 21548
rect 24995 21508 25228 21536
rect 24995 21505 25007 21508
rect 24949 21499 25007 21505
rect 25222 21496 25228 21508
rect 25280 21496 25286 21548
rect 25409 21539 25467 21545
rect 25409 21505 25421 21539
rect 25455 21505 25467 21539
rect 25409 21499 25467 21505
rect 26145 21539 26203 21545
rect 26145 21505 26157 21539
rect 26191 21505 26203 21539
rect 26145 21499 26203 21505
rect 25424 21468 25452 21499
rect 23676 21440 25452 21468
rect 25958 21400 25964 21412
rect 23492 21372 25964 21400
rect 23017 21363 23075 21369
rect 25958 21360 25964 21372
rect 26016 21360 26022 21412
rect 26160 21400 26188 21499
rect 27172 21468 27200 21576
rect 29914 21564 29920 21576
rect 29972 21564 29978 21616
rect 30374 21604 30380 21616
rect 30116 21576 30380 21604
rect 27338 21536 27344 21548
rect 27299 21508 27344 21536
rect 27338 21496 27344 21508
rect 27396 21496 27402 21548
rect 30116 21545 30144 21576
rect 30374 21564 30380 21576
rect 30432 21564 30438 21616
rect 28169 21539 28227 21545
rect 28169 21505 28181 21539
rect 28215 21505 28227 21539
rect 28169 21499 28227 21505
rect 30101 21539 30159 21545
rect 30101 21505 30113 21539
rect 30147 21505 30159 21539
rect 30282 21536 30288 21548
rect 30243 21508 30288 21536
rect 30101 21499 30159 21505
rect 27249 21471 27307 21477
rect 27249 21468 27261 21471
rect 27172 21440 27261 21468
rect 27249 21437 27261 21440
rect 27295 21437 27307 21471
rect 27706 21468 27712 21480
rect 27667 21440 27712 21468
rect 27249 21431 27307 21437
rect 27706 21428 27712 21440
rect 27764 21428 27770 21480
rect 28184 21468 28212 21499
rect 30282 21496 30288 21508
rect 30340 21496 30346 21548
rect 31205 21539 31263 21545
rect 31205 21505 31217 21539
rect 31251 21536 31263 21539
rect 31386 21536 31392 21548
rect 31251 21508 31392 21536
rect 31251 21505 31263 21508
rect 31205 21499 31263 21505
rect 31220 21468 31248 21499
rect 31386 21496 31392 21508
rect 31444 21496 31450 21548
rect 28184 21440 31248 21468
rect 28184 21400 28212 21440
rect 26160 21372 28212 21400
rect 35866 21400 35894 21644
rect 42058 21632 42064 21684
rect 42116 21672 42122 21684
rect 46198 21672 46204 21684
rect 42116 21644 44128 21672
rect 46159 21644 46204 21672
rect 42116 21632 42122 21644
rect 43990 21604 43996 21616
rect 43951 21576 43996 21604
rect 43990 21564 43996 21576
rect 44048 21564 44054 21616
rect 44100 21604 44128 21644
rect 46198 21632 46204 21644
rect 46256 21632 46262 21684
rect 47946 21604 47952 21616
rect 44100 21576 46704 21604
rect 47907 21576 47952 21604
rect 46676 21548 46704 21576
rect 47946 21564 47952 21576
rect 48004 21564 48010 21616
rect 45830 21536 45836 21548
rect 45204 21508 45836 21536
rect 43809 21471 43867 21477
rect 43809 21437 43821 21471
rect 43855 21468 43867 21471
rect 45204 21468 45232 21508
rect 45830 21496 45836 21508
rect 45888 21496 45894 21548
rect 45922 21496 45928 21548
rect 45980 21536 45986 21548
rect 46109 21539 46167 21545
rect 46109 21536 46121 21539
rect 45980 21508 46121 21536
rect 45980 21496 45986 21508
rect 46109 21505 46121 21508
rect 46155 21505 46167 21539
rect 46290 21536 46296 21548
rect 46251 21508 46296 21536
rect 46109 21499 46167 21505
rect 46290 21496 46296 21508
rect 46348 21496 46354 21548
rect 46658 21496 46664 21548
rect 46716 21536 46722 21548
rect 46845 21539 46903 21545
rect 46845 21536 46857 21539
rect 46716 21508 46857 21536
rect 46716 21496 46722 21508
rect 46845 21505 46857 21508
rect 46891 21505 46903 21539
rect 46845 21499 46903 21505
rect 45370 21468 45376 21480
rect 43855 21440 45232 21468
rect 45331 21440 45376 21468
rect 43855 21437 43867 21440
rect 43809 21431 43867 21437
rect 45370 21428 45376 21440
rect 45428 21428 45434 21480
rect 48133 21403 48191 21409
rect 48133 21400 48145 21403
rect 35866 21372 48145 21400
rect 10410 21292 10416 21344
rect 10468 21332 10474 21344
rect 12069 21335 12127 21341
rect 12069 21332 12081 21335
rect 10468 21304 12081 21332
rect 10468 21292 10474 21304
rect 12069 21301 12081 21304
rect 12115 21301 12127 21335
rect 13354 21332 13360 21344
rect 13315 21304 13360 21332
rect 12069 21295 12127 21301
rect 13354 21292 13360 21304
rect 13412 21292 13418 21344
rect 15381 21335 15439 21341
rect 15381 21301 15393 21335
rect 15427 21332 15439 21335
rect 15838 21332 15844 21344
rect 15427 21304 15844 21332
rect 15427 21301 15439 21304
rect 15381 21295 15439 21301
rect 15838 21292 15844 21304
rect 15896 21292 15902 21344
rect 20257 21335 20315 21341
rect 20257 21301 20269 21335
rect 20303 21332 20315 21335
rect 21082 21332 21088 21344
rect 20303 21304 21088 21332
rect 20303 21301 20315 21304
rect 20257 21295 20315 21301
rect 21082 21292 21088 21304
rect 21140 21292 21146 21344
rect 22370 21292 22376 21344
rect 22428 21332 22434 21344
rect 22557 21335 22615 21341
rect 22557 21332 22569 21335
rect 22428 21304 22569 21332
rect 22428 21292 22434 21304
rect 22557 21301 22569 21304
rect 22603 21301 22615 21335
rect 22557 21295 22615 21301
rect 23658 21292 23664 21344
rect 23716 21332 23722 21344
rect 23845 21335 23903 21341
rect 23845 21332 23857 21335
rect 23716 21304 23857 21332
rect 23716 21292 23722 21304
rect 23845 21301 23857 21304
rect 23891 21301 23903 21335
rect 23845 21295 23903 21301
rect 25593 21335 25651 21341
rect 25593 21301 25605 21335
rect 25639 21332 25651 21335
rect 26160 21332 26188 21372
rect 48133 21369 48145 21372
rect 48179 21369 48191 21403
rect 48133 21363 48191 21369
rect 25639 21304 26188 21332
rect 30101 21335 30159 21341
rect 25639 21301 25651 21304
rect 25593 21295 25651 21301
rect 30101 21301 30113 21335
rect 30147 21332 30159 21335
rect 30466 21332 30472 21344
rect 30147 21304 30472 21332
rect 30147 21301 30159 21304
rect 30101 21295 30159 21301
rect 30466 21292 30472 21304
rect 30524 21292 30530 21344
rect 31202 21292 31208 21344
rect 31260 21332 31266 21344
rect 31297 21335 31355 21341
rect 31297 21332 31309 21335
rect 31260 21304 31309 21332
rect 31260 21292 31266 21304
rect 31297 21301 31309 21304
rect 31343 21301 31355 21335
rect 31297 21295 31355 21301
rect 46474 21292 46480 21344
rect 46532 21332 46538 21344
rect 46937 21335 46995 21341
rect 46937 21332 46949 21335
rect 46532 21304 46949 21332
rect 46532 21292 46538 21304
rect 46937 21301 46949 21304
rect 46983 21301 46995 21335
rect 46937 21295 46995 21301
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 9122 21088 9128 21140
rect 9180 21128 9186 21140
rect 9217 21131 9275 21137
rect 9217 21128 9229 21131
rect 9180 21100 9229 21128
rect 9180 21088 9186 21100
rect 9217 21097 9229 21100
rect 9263 21097 9275 21131
rect 9217 21091 9275 21097
rect 10134 21088 10140 21140
rect 10192 21128 10198 21140
rect 10229 21131 10287 21137
rect 10229 21128 10241 21131
rect 10192 21100 10241 21128
rect 10192 21088 10198 21100
rect 10229 21097 10241 21100
rect 10275 21097 10287 21131
rect 10229 21091 10287 21097
rect 15930 21088 15936 21140
rect 15988 21128 15994 21140
rect 18141 21131 18199 21137
rect 18141 21128 18153 21131
rect 15988 21100 18153 21128
rect 15988 21088 15994 21100
rect 18141 21097 18153 21100
rect 18187 21097 18199 21131
rect 18141 21091 18199 21097
rect 19978 21088 19984 21140
rect 20036 21128 20042 21140
rect 20257 21131 20315 21137
rect 20257 21128 20269 21131
rect 20036 21100 20269 21128
rect 20036 21088 20042 21100
rect 20257 21097 20269 21100
rect 20303 21097 20315 21131
rect 20257 21091 20315 21097
rect 20990 21088 20996 21140
rect 21048 21128 21054 21140
rect 21085 21131 21143 21137
rect 21085 21128 21097 21131
rect 21048 21100 21097 21128
rect 21048 21088 21054 21100
rect 21085 21097 21097 21100
rect 21131 21097 21143 21131
rect 21085 21091 21143 21097
rect 22066 21100 31754 21128
rect 22066 21060 22094 21100
rect 17512 21032 22094 21060
rect 26053 21063 26111 21069
rect 11977 20995 12035 21001
rect 11977 20992 11989 20995
rect 2746 20964 11989 20992
rect 14 20816 20 20868
rect 72 20856 78 20868
rect 2746 20856 2774 20964
rect 11977 20961 11989 20964
rect 12023 20961 12035 20995
rect 15838 20992 15844 21004
rect 15799 20964 15844 20992
rect 11977 20955 12035 20961
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 17512 21001 17540 21032
rect 26053 21029 26065 21063
rect 26099 21060 26111 21063
rect 26878 21060 26884 21072
rect 26099 21032 26884 21060
rect 26099 21029 26111 21032
rect 26053 21023 26111 21029
rect 26878 21020 26884 21032
rect 26936 21020 26942 21072
rect 17497 20995 17555 21001
rect 17497 20961 17509 20995
rect 17543 20961 17555 20995
rect 17497 20955 17555 20961
rect 20070 20952 20076 21004
rect 20128 20992 20134 21004
rect 20128 20964 21036 20992
rect 20128 20952 20134 20964
rect 9398 20924 9404 20936
rect 9359 20896 9404 20924
rect 9398 20884 9404 20896
rect 9456 20884 9462 20936
rect 10137 20927 10195 20933
rect 10137 20893 10149 20927
rect 10183 20924 10195 20927
rect 10410 20924 10416 20936
rect 10183 20896 10416 20924
rect 10183 20893 10195 20896
rect 10137 20887 10195 20893
rect 10410 20884 10416 20896
rect 10468 20884 10474 20936
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20924 10931 20927
rect 11054 20924 11060 20936
rect 10919 20896 11060 20924
rect 10919 20893 10931 20896
rect 10873 20887 10931 20893
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 11514 20924 11520 20936
rect 11475 20896 11520 20924
rect 11514 20884 11520 20896
rect 11572 20884 11578 20936
rect 13354 20884 13360 20936
rect 13412 20924 13418 20936
rect 14553 20927 14611 20933
rect 14553 20924 14565 20927
rect 13412 20896 14565 20924
rect 13412 20884 13418 20896
rect 14553 20893 14565 20896
rect 14599 20893 14611 20927
rect 15654 20924 15660 20936
rect 15615 20896 15660 20924
rect 14553 20887 14611 20893
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 17862 20884 17868 20936
rect 17920 20924 17926 20936
rect 18049 20927 18107 20933
rect 18049 20924 18061 20927
rect 17920 20896 18061 20924
rect 17920 20884 17926 20896
rect 18049 20893 18061 20896
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20924 19303 20927
rect 19426 20924 19432 20936
rect 19291 20896 19432 20924
rect 19291 20893 19303 20896
rect 19245 20887 19303 20893
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 20438 20924 20444 20936
rect 20399 20896 20444 20924
rect 20438 20884 20444 20896
rect 20496 20884 20502 20936
rect 21008 20933 21036 20964
rect 22094 20952 22100 21004
rect 22152 20992 22158 21004
rect 22370 20992 22376 21004
rect 22152 20964 22197 20992
rect 22331 20964 22376 20992
rect 22152 20952 22158 20964
rect 22370 20952 22376 20964
rect 22428 20952 22434 21004
rect 30466 20992 30472 21004
rect 30427 20964 30472 20992
rect 30466 20952 30472 20964
rect 30524 20952 30530 21004
rect 31726 20992 31754 21100
rect 46382 21060 46388 21072
rect 35866 21032 46388 21060
rect 35866 20992 35894 21032
rect 46382 21020 46388 21032
rect 46440 21020 46446 21072
rect 46474 20992 46480 21004
rect 31726 20964 35894 20992
rect 46435 20964 46480 20992
rect 46474 20952 46480 20964
rect 46532 20952 46538 21004
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 20993 20927 21051 20933
rect 20993 20893 21005 20927
rect 21039 20924 21051 20927
rect 21818 20924 21824 20936
rect 21039 20896 21824 20924
rect 21039 20893 21051 20896
rect 20993 20887 21051 20893
rect 21818 20884 21824 20896
rect 21876 20884 21882 20936
rect 25958 20924 25964 20936
rect 25919 20896 25964 20924
rect 25958 20884 25964 20896
rect 26016 20884 26022 20936
rect 30190 20924 30196 20936
rect 30151 20896 30196 20924
rect 30190 20884 30196 20896
rect 30248 20884 30254 20936
rect 33321 20927 33379 20933
rect 33321 20893 33333 20927
rect 33367 20924 33379 20927
rect 33410 20924 33416 20936
rect 33367 20896 33416 20924
rect 33367 20893 33379 20896
rect 33321 20887 33379 20893
rect 33410 20884 33416 20896
rect 33468 20884 33474 20936
rect 43717 20927 43775 20933
rect 43717 20893 43729 20927
rect 43763 20924 43775 20927
rect 45554 20924 45560 20936
rect 43763 20896 45560 20924
rect 43763 20893 43775 20896
rect 43717 20887 43775 20893
rect 45554 20884 45560 20896
rect 45612 20884 45618 20936
rect 46293 20927 46351 20933
rect 46293 20893 46305 20927
rect 46339 20893 46351 20927
rect 46293 20887 46351 20893
rect 72 20828 2774 20856
rect 10965 20859 11023 20865
rect 72 20816 78 20828
rect 10965 20825 10977 20859
rect 11011 20856 11023 20859
rect 11701 20859 11759 20865
rect 11701 20856 11713 20859
rect 11011 20828 11713 20856
rect 11011 20825 11023 20828
rect 10965 20819 11023 20825
rect 11701 20825 11713 20828
rect 11747 20825 11759 20859
rect 23658 20856 23664 20868
rect 23598 20828 23664 20856
rect 11701 20819 11759 20825
rect 23658 20816 23664 20828
rect 23716 20816 23722 20868
rect 31202 20816 31208 20868
rect 31260 20816 31266 20868
rect 46308 20856 46336 20887
rect 47762 20856 47768 20868
rect 46308 20828 47768 20856
rect 47762 20816 47768 20828
rect 47820 20816 47826 20868
rect 14642 20788 14648 20800
rect 14603 20760 14648 20788
rect 14642 20748 14648 20760
rect 14700 20748 14706 20800
rect 19334 20788 19340 20800
rect 19295 20760 19340 20788
rect 19334 20748 19340 20760
rect 19392 20748 19398 20800
rect 22186 20748 22192 20800
rect 22244 20788 22250 20800
rect 23845 20791 23903 20797
rect 23845 20788 23857 20791
rect 22244 20760 23857 20788
rect 22244 20748 22250 20760
rect 23845 20757 23857 20760
rect 23891 20788 23903 20791
rect 23934 20788 23940 20800
rect 23891 20760 23940 20788
rect 23891 20757 23903 20760
rect 23845 20751 23903 20757
rect 23934 20748 23940 20760
rect 23992 20748 23998 20800
rect 31938 20788 31944 20800
rect 31899 20760 31944 20788
rect 31938 20748 31944 20760
rect 31996 20748 32002 20800
rect 33318 20748 33324 20800
rect 33376 20788 33382 20800
rect 33413 20791 33471 20797
rect 33413 20788 33425 20791
rect 33376 20760 33425 20788
rect 33376 20748 33382 20760
rect 33413 20757 33425 20760
rect 33459 20757 33471 20791
rect 43806 20788 43812 20800
rect 43767 20760 43812 20788
rect 33413 20751 33471 20757
rect 43806 20748 43812 20760
rect 43864 20748 43870 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 3970 20544 3976 20596
rect 4028 20584 4034 20596
rect 15381 20587 15439 20593
rect 4028 20556 15332 20584
rect 4028 20544 4034 20556
rect 9398 20516 9404 20528
rect 9311 20488 9404 20516
rect 9324 20457 9352 20488
rect 9398 20476 9404 20488
rect 9456 20516 9462 20528
rect 13078 20516 13084 20528
rect 9456 20488 13084 20516
rect 9456 20476 9462 20488
rect 9309 20451 9367 20457
rect 9309 20417 9321 20451
rect 9355 20417 9367 20451
rect 9309 20411 9367 20417
rect 9953 20451 10011 20457
rect 9953 20417 9965 20451
rect 9999 20448 10011 20451
rect 10410 20448 10416 20460
rect 9999 20420 10416 20448
rect 9999 20417 10011 20420
rect 9953 20411 10011 20417
rect 10410 20408 10416 20420
rect 10468 20408 10474 20460
rect 12360 20457 12388 20488
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 14182 20516 14188 20528
rect 13648 20488 14188 20516
rect 12345 20451 12403 20457
rect 12345 20417 12357 20451
rect 12391 20417 12403 20451
rect 12345 20411 12403 20417
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20448 12955 20451
rect 12986 20448 12992 20460
rect 12943 20420 12992 20448
rect 12943 20417 12955 20420
rect 12897 20411 12955 20417
rect 12986 20408 12992 20420
rect 13044 20448 13050 20460
rect 13648 20448 13676 20488
rect 14182 20476 14188 20488
rect 14240 20476 14246 20528
rect 14642 20476 14648 20528
rect 14700 20476 14706 20528
rect 15304 20516 15332 20556
rect 15381 20553 15393 20587
rect 15427 20584 15439 20587
rect 15654 20584 15660 20596
rect 15427 20556 15660 20584
rect 15427 20553 15439 20556
rect 15381 20547 15439 20553
rect 15654 20544 15660 20556
rect 15712 20544 15718 20596
rect 17770 20544 17776 20596
rect 17828 20584 17834 20596
rect 17828 20556 20287 20584
rect 17828 20544 17834 20556
rect 17954 20516 17960 20528
rect 15304 20488 17960 20516
rect 17954 20476 17960 20488
rect 18012 20476 18018 20528
rect 20162 20516 20168 20528
rect 19826 20488 20168 20516
rect 20162 20476 20168 20488
rect 20220 20476 20226 20528
rect 13044 20420 13676 20448
rect 17037 20451 17095 20457
rect 13044 20408 13050 20420
rect 17037 20417 17049 20451
rect 17083 20448 17095 20451
rect 17218 20448 17224 20460
rect 17083 20420 17224 20448
rect 17083 20417 17095 20420
rect 17037 20411 17095 20417
rect 17218 20408 17224 20420
rect 17276 20448 17282 20460
rect 17862 20448 17868 20460
rect 17276 20420 17868 20448
rect 17276 20408 17282 20420
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 20259 20448 20287 20556
rect 21082 20544 21088 20596
rect 21140 20584 21146 20596
rect 21818 20584 21824 20596
rect 21140 20556 21824 20584
rect 21140 20544 21146 20556
rect 21818 20544 21824 20556
rect 21876 20584 21882 20596
rect 28534 20584 28540 20596
rect 21876 20556 28540 20584
rect 21876 20544 21882 20556
rect 28534 20544 28540 20556
rect 28592 20544 28598 20596
rect 30190 20584 30196 20596
rect 30151 20556 30196 20584
rect 30190 20544 30196 20556
rect 30248 20544 30254 20596
rect 20438 20476 20444 20528
rect 20496 20516 20502 20528
rect 27890 20516 27896 20528
rect 20496 20488 27896 20516
rect 20496 20476 20502 20488
rect 27890 20476 27896 20488
rect 27948 20476 27954 20528
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 20259 20420 21833 20448
rect 21821 20417 21833 20420
rect 21867 20448 21879 20451
rect 22370 20448 22376 20460
rect 21867 20420 22376 20448
rect 21867 20417 21879 20420
rect 21821 20411 21879 20417
rect 22370 20408 22376 20420
rect 22428 20448 22434 20460
rect 23014 20448 23020 20460
rect 22428 20420 23020 20448
rect 22428 20408 22434 20420
rect 23014 20408 23020 20420
rect 23072 20408 23078 20460
rect 23198 20408 23204 20460
rect 23256 20448 23262 20460
rect 24857 20451 24915 20457
rect 24857 20448 24869 20451
rect 23256 20420 24869 20448
rect 23256 20408 23262 20420
rect 24857 20417 24869 20420
rect 24903 20417 24915 20451
rect 26234 20448 26240 20460
rect 26195 20420 26240 20448
rect 24857 20411 24915 20417
rect 26234 20408 26240 20420
rect 26292 20408 26298 20460
rect 27430 20448 27436 20460
rect 27391 20420 27436 20448
rect 27430 20408 27436 20420
rect 27488 20408 27494 20460
rect 27706 20408 27712 20460
rect 27764 20448 27770 20460
rect 28077 20451 28135 20457
rect 28077 20448 28089 20451
rect 27764 20420 28089 20448
rect 27764 20408 27770 20420
rect 28077 20417 28089 20420
rect 28123 20417 28135 20451
rect 28552 20448 28580 20544
rect 33318 20516 33324 20528
rect 33279 20488 33324 20516
rect 33318 20476 33324 20488
rect 33376 20476 33382 20528
rect 43806 20516 43812 20528
rect 43767 20488 43812 20516
rect 43806 20476 43812 20488
rect 43864 20476 43870 20528
rect 30009 20451 30067 20457
rect 30009 20448 30021 20451
rect 28552 20420 30021 20448
rect 28077 20411 28135 20417
rect 30009 20417 30021 20420
rect 30055 20417 30067 20451
rect 30009 20411 30067 20417
rect 31938 20408 31944 20460
rect 31996 20448 32002 20460
rect 33137 20451 33195 20457
rect 33137 20448 33149 20451
rect 31996 20420 33149 20448
rect 31996 20408 32002 20420
rect 33137 20417 33149 20420
rect 33183 20417 33195 20451
rect 46382 20448 46388 20460
rect 46343 20420 46388 20448
rect 33137 20411 33195 20417
rect 46382 20408 46388 20420
rect 46440 20408 46446 20460
rect 46845 20451 46903 20457
rect 46845 20417 46857 20451
rect 46891 20448 46903 20451
rect 46934 20448 46940 20460
rect 46891 20420 46940 20448
rect 46891 20417 46903 20420
rect 46845 20411 46903 20417
rect 46934 20408 46940 20420
rect 46992 20408 46998 20460
rect 47762 20448 47768 20460
rect 47723 20420 47768 20448
rect 47762 20408 47768 20420
rect 47820 20408 47826 20460
rect 12437 20383 12495 20389
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 13633 20383 13691 20389
rect 13633 20380 13645 20383
rect 12483 20352 13645 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 13633 20349 13645 20352
rect 13679 20349 13691 20383
rect 13906 20380 13912 20392
rect 13867 20352 13912 20380
rect 13633 20343 13691 20349
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 17678 20380 17684 20392
rect 17639 20352 17684 20380
rect 17678 20340 17684 20352
rect 17736 20340 17742 20392
rect 18046 20340 18052 20392
rect 18104 20380 18110 20392
rect 18325 20383 18383 20389
rect 18325 20380 18337 20383
rect 18104 20352 18337 20380
rect 18104 20340 18110 20352
rect 18325 20349 18337 20352
rect 18371 20349 18383 20383
rect 18325 20343 18383 20349
rect 18601 20383 18659 20389
rect 18601 20349 18613 20383
rect 18647 20380 18659 20383
rect 19334 20380 19340 20392
rect 18647 20352 19340 20380
rect 18647 20349 18659 20352
rect 18601 20343 18659 20349
rect 19334 20340 19340 20352
rect 19392 20340 19398 20392
rect 25958 20380 25964 20392
rect 19628 20352 25964 20380
rect 3234 20272 3240 20324
rect 3292 20312 3298 20324
rect 3292 20284 13768 20312
rect 3292 20272 3298 20284
rect 8938 20204 8944 20256
rect 8996 20244 9002 20256
rect 9125 20247 9183 20253
rect 9125 20244 9137 20247
rect 8996 20216 9137 20244
rect 8996 20204 9002 20216
rect 9125 20213 9137 20216
rect 9171 20213 9183 20247
rect 9125 20207 9183 20213
rect 9950 20204 9956 20256
rect 10008 20244 10014 20256
rect 10045 20247 10103 20253
rect 10045 20244 10057 20247
rect 10008 20216 10057 20244
rect 10008 20204 10014 20216
rect 10045 20213 10057 20216
rect 10091 20213 10103 20247
rect 13078 20244 13084 20256
rect 13039 20216 13084 20244
rect 10045 20207 10103 20213
rect 13078 20204 13084 20216
rect 13136 20204 13142 20256
rect 13740 20244 13768 20284
rect 14936 20284 17264 20312
rect 14936 20244 14964 20284
rect 13740 20216 14964 20244
rect 17236 20244 17264 20284
rect 19628 20244 19656 20352
rect 25958 20340 25964 20352
rect 26016 20340 26022 20392
rect 34977 20383 35035 20389
rect 34977 20349 34989 20383
rect 35023 20380 35035 20383
rect 35434 20380 35440 20392
rect 35023 20352 35440 20380
rect 35023 20349 35035 20352
rect 34977 20343 35035 20349
rect 35434 20340 35440 20352
rect 35492 20340 35498 20392
rect 43625 20383 43683 20389
rect 43625 20380 43637 20383
rect 35866 20352 43637 20380
rect 19978 20272 19984 20324
rect 20036 20312 20042 20324
rect 24578 20312 24584 20324
rect 20036 20284 24584 20312
rect 20036 20272 20042 20284
rect 24578 20272 24584 20284
rect 24636 20272 24642 20324
rect 25038 20312 25044 20324
rect 24999 20284 25044 20312
rect 25038 20272 25044 20284
rect 25096 20272 25102 20324
rect 26694 20272 26700 20324
rect 26752 20312 26758 20324
rect 28261 20315 28319 20321
rect 28261 20312 28273 20315
rect 26752 20284 28273 20312
rect 26752 20272 26758 20284
rect 28261 20281 28273 20284
rect 28307 20312 28319 20315
rect 35866 20312 35894 20352
rect 43625 20349 43637 20352
rect 43671 20349 43683 20383
rect 45462 20380 45468 20392
rect 45423 20352 45468 20380
rect 43625 20343 43683 20349
rect 45462 20340 45468 20352
rect 45520 20340 45526 20392
rect 45554 20340 45560 20392
rect 45612 20380 45618 20392
rect 46017 20383 46075 20389
rect 46017 20380 46029 20383
rect 45612 20352 46029 20380
rect 45612 20340 45618 20352
rect 46017 20349 46029 20352
rect 46063 20349 46075 20383
rect 46017 20343 46075 20349
rect 46750 20312 46756 20324
rect 28307 20284 35894 20312
rect 46711 20284 46756 20312
rect 28307 20281 28319 20284
rect 28261 20275 28319 20281
rect 46750 20272 46756 20284
rect 46808 20272 46814 20324
rect 20070 20244 20076 20256
rect 17236 20216 19656 20244
rect 20031 20216 20076 20244
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 21910 20244 21916 20256
rect 21871 20216 21916 20244
rect 21910 20204 21916 20216
rect 21968 20204 21974 20256
rect 23014 20204 23020 20256
rect 23072 20244 23078 20256
rect 23382 20244 23388 20256
rect 23072 20216 23388 20244
rect 23072 20204 23078 20216
rect 23382 20204 23388 20216
rect 23440 20204 23446 20256
rect 26329 20247 26387 20253
rect 26329 20213 26341 20247
rect 26375 20244 26387 20247
rect 27338 20244 27344 20256
rect 26375 20216 27344 20244
rect 26375 20213 26387 20216
rect 26329 20207 26387 20213
rect 27338 20204 27344 20216
rect 27396 20204 27402 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 10594 20000 10600 20052
rect 10652 20040 10658 20052
rect 10689 20043 10747 20049
rect 10689 20040 10701 20043
rect 10652 20012 10701 20040
rect 10652 20000 10658 20012
rect 10689 20009 10701 20012
rect 10735 20009 10747 20043
rect 10689 20003 10747 20009
rect 13541 20043 13599 20049
rect 13541 20009 13553 20043
rect 13587 20040 13599 20043
rect 13906 20040 13912 20052
rect 13587 20012 13912 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 14645 20043 14703 20049
rect 14645 20040 14657 20043
rect 14608 20012 14657 20040
rect 14608 20000 14614 20012
rect 14645 20009 14657 20012
rect 14691 20009 14703 20043
rect 14645 20003 14703 20009
rect 20346 20000 20352 20052
rect 20404 20040 20410 20052
rect 20404 20012 23336 20040
rect 20404 20000 20410 20012
rect 13170 19972 13176 19984
rect 12406 19944 13176 19972
rect 8938 19904 8944 19916
rect 8899 19876 8944 19904
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 11514 19864 11520 19916
rect 11572 19904 11578 19916
rect 12406 19904 12434 19944
rect 13170 19932 13176 19944
rect 13228 19972 13234 19984
rect 14093 19975 14151 19981
rect 14093 19972 14105 19975
rect 13228 19944 14105 19972
rect 13228 19932 13234 19944
rect 14093 19941 14105 19944
rect 14139 19941 14151 19975
rect 14093 19935 14151 19941
rect 14182 19932 14188 19984
rect 14240 19972 14246 19984
rect 20070 19972 20076 19984
rect 14240 19944 20076 19972
rect 14240 19932 14246 19944
rect 20070 19932 20076 19944
rect 20128 19932 20134 19984
rect 21450 19932 21456 19984
rect 21508 19972 21514 19984
rect 21508 19944 22232 19972
rect 21508 19932 21514 19944
rect 11572 19876 12434 19904
rect 13265 19907 13323 19913
rect 11572 19864 11578 19876
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 11422 19836 11428 19848
rect 11383 19808 11428 19836
rect 2041 19799 2099 19805
rect 11422 19796 11428 19808
rect 11480 19796 11486 19848
rect 11900 19845 11928 19876
rect 13265 19873 13277 19907
rect 13311 19904 13323 19907
rect 14458 19904 14464 19916
rect 13311 19876 14464 19904
rect 13311 19873 13323 19876
rect 13265 19867 13323 19873
rect 14458 19864 14464 19876
rect 14516 19864 14522 19916
rect 17770 19864 17776 19916
rect 17828 19904 17834 19916
rect 17957 19907 18015 19913
rect 17957 19904 17969 19907
rect 17828 19876 17969 19904
rect 17828 19864 17834 19876
rect 17957 19873 17969 19876
rect 18003 19873 18015 19907
rect 17957 19867 18015 19873
rect 18046 19864 18052 19916
rect 18104 19904 18110 19916
rect 20438 19904 20444 19916
rect 18104 19876 20444 19904
rect 18104 19864 18110 19876
rect 20438 19864 20444 19876
rect 20496 19864 20502 19916
rect 21910 19904 21916 19916
rect 21871 19876 21916 19904
rect 21910 19864 21916 19876
rect 21968 19864 21974 19916
rect 22204 19913 22232 19944
rect 22189 19907 22247 19913
rect 22189 19873 22201 19907
rect 22235 19873 22247 19907
rect 22189 19867 22247 19873
rect 11701 19839 11759 19845
rect 11701 19805 11713 19839
rect 11747 19805 11759 19839
rect 11701 19799 11759 19805
rect 11885 19839 11943 19845
rect 11885 19805 11897 19839
rect 11931 19805 11943 19839
rect 11885 19799 11943 19805
rect 13173 19839 13231 19845
rect 13173 19805 13185 19839
rect 13219 19836 13231 19839
rect 13906 19836 13912 19848
rect 13219 19808 13912 19836
rect 13219 19805 13231 19808
rect 13173 19799 13231 19805
rect 9214 19768 9220 19780
rect 9175 19740 9220 19768
rect 9214 19728 9220 19740
rect 9272 19728 9278 19780
rect 9950 19728 9956 19780
rect 10008 19728 10014 19780
rect 11716 19768 11744 19799
rect 13906 19796 13912 19808
rect 13964 19836 13970 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 13964 19808 14289 19836
rect 13964 19796 13970 19808
rect 14277 19805 14289 19808
rect 14323 19836 14335 19839
rect 15654 19836 15660 19848
rect 14323 19808 15660 19836
rect 14323 19805 14335 19808
rect 14277 19799 14335 19805
rect 15654 19796 15660 19808
rect 15712 19796 15718 19848
rect 16393 19839 16451 19845
rect 16393 19805 16405 19839
rect 16439 19836 16451 19839
rect 17218 19836 17224 19848
rect 16439 19808 17224 19836
rect 16439 19805 16451 19808
rect 16393 19799 16451 19805
rect 17218 19796 17224 19808
rect 17276 19796 17282 19848
rect 19426 19836 19432 19848
rect 19387 19808 19432 19836
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 20809 19839 20867 19845
rect 20809 19805 20821 19839
rect 20855 19836 20867 19839
rect 21729 19839 21787 19845
rect 20855 19808 21680 19836
rect 20855 19805 20867 19808
rect 20809 19799 20867 19805
rect 13722 19768 13728 19780
rect 11716 19740 13728 19768
rect 13722 19728 13728 19740
rect 13780 19728 13786 19780
rect 14182 19728 14188 19780
rect 14240 19768 14246 19780
rect 14461 19771 14519 19777
rect 14461 19768 14473 19771
rect 14240 19740 14473 19768
rect 14240 19728 14246 19740
rect 14461 19737 14473 19740
rect 14507 19737 14519 19771
rect 14461 19731 14519 19737
rect 17678 19728 17684 19780
rect 17736 19768 17742 19780
rect 20346 19768 20352 19780
rect 17736 19740 20352 19768
rect 17736 19728 17742 19740
rect 20346 19728 20352 19740
rect 20404 19728 20410 19780
rect 11238 19700 11244 19712
rect 11199 19672 11244 19700
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 11330 19660 11336 19712
rect 11388 19700 11394 19712
rect 13078 19700 13084 19712
rect 11388 19672 13084 19700
rect 11388 19660 11394 19672
rect 13078 19660 13084 19672
rect 13136 19660 13142 19712
rect 14090 19660 14096 19712
rect 14148 19700 14154 19712
rect 14369 19703 14427 19709
rect 14369 19700 14381 19703
rect 14148 19672 14381 19700
rect 14148 19660 14154 19672
rect 14369 19669 14381 19672
rect 14415 19669 14427 19703
rect 14369 19663 14427 19669
rect 15654 19660 15660 19712
rect 15712 19700 15718 19712
rect 16577 19703 16635 19709
rect 16577 19700 16589 19703
rect 15712 19672 16589 19700
rect 15712 19660 15718 19672
rect 16577 19669 16589 19672
rect 16623 19669 16635 19703
rect 16577 19663 16635 19669
rect 18414 19660 18420 19712
rect 18472 19700 18478 19712
rect 19429 19703 19487 19709
rect 19429 19700 19441 19703
rect 18472 19672 19441 19700
rect 18472 19660 18478 19672
rect 19429 19669 19441 19672
rect 19475 19669 19487 19703
rect 19429 19663 19487 19669
rect 20162 19660 20168 19712
rect 20220 19700 20226 19712
rect 20993 19703 21051 19709
rect 20993 19700 21005 19703
rect 20220 19672 21005 19700
rect 20220 19660 20226 19672
rect 20993 19669 21005 19672
rect 21039 19669 21051 19703
rect 21652 19700 21680 19808
rect 21729 19805 21741 19839
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 21744 19768 21772 19799
rect 22186 19768 22192 19780
rect 21744 19740 22192 19768
rect 22186 19728 22192 19740
rect 22244 19728 22250 19780
rect 23198 19700 23204 19712
rect 21652 19672 23204 19700
rect 20993 19663 21051 19669
rect 23198 19660 23204 19672
rect 23256 19660 23262 19712
rect 23308 19700 23336 20012
rect 23382 20000 23388 20052
rect 23440 20040 23446 20052
rect 26973 20043 27031 20049
rect 23440 20012 26280 20040
rect 23440 20000 23446 20012
rect 24489 19907 24547 19913
rect 24489 19873 24501 19907
rect 24535 19904 24547 19907
rect 24578 19904 24584 19916
rect 24535 19876 24584 19904
rect 24535 19873 24547 19876
rect 24489 19867 24547 19873
rect 24578 19864 24584 19876
rect 24636 19864 24642 19916
rect 25501 19907 25559 19913
rect 25501 19873 25513 19907
rect 25547 19904 25559 19907
rect 26050 19904 26056 19916
rect 25547 19876 26056 19904
rect 25547 19873 25559 19876
rect 25501 19867 25559 19873
rect 26050 19864 26056 19876
rect 26108 19864 26114 19916
rect 26252 19904 26280 20012
rect 26973 20009 26985 20043
rect 27019 20040 27031 20043
rect 27430 20040 27436 20052
rect 27019 20012 27436 20040
rect 27019 20009 27031 20012
rect 26973 20003 27031 20009
rect 27430 20000 27436 20012
rect 27488 20000 27494 20052
rect 41322 20040 41328 20052
rect 27540 20012 41328 20040
rect 26510 19932 26516 19984
rect 26568 19972 26574 19984
rect 27540 19972 27568 20012
rect 41322 20000 41328 20012
rect 41380 20000 41386 20052
rect 46934 20000 46940 20052
rect 46992 20040 46998 20052
rect 47765 20043 47823 20049
rect 47765 20040 47777 20043
rect 46992 20012 47777 20040
rect 46992 20000 46998 20012
rect 47765 20009 47777 20012
rect 47811 20009 47823 20043
rect 47765 20003 47823 20009
rect 27706 19972 27712 19984
rect 26568 19944 27568 19972
rect 27667 19944 27712 19972
rect 26568 19932 26574 19944
rect 27706 19932 27712 19944
rect 27764 19932 27770 19984
rect 45465 19975 45523 19981
rect 45465 19941 45477 19975
rect 45511 19972 45523 19975
rect 46952 19972 46980 20000
rect 45511 19944 46980 19972
rect 45511 19941 45523 19944
rect 45465 19935 45523 19941
rect 29178 19904 29184 19916
rect 26252 19876 29184 19904
rect 29178 19864 29184 19876
rect 29236 19864 29242 19916
rect 44361 19907 44419 19913
rect 44361 19873 44373 19907
rect 44407 19904 44419 19907
rect 45189 19907 45247 19913
rect 45189 19904 45201 19907
rect 44407 19876 45201 19904
rect 44407 19873 44419 19876
rect 44361 19867 44419 19873
rect 45189 19873 45201 19876
rect 45235 19904 45247 19907
rect 45554 19904 45560 19916
rect 45235 19876 45560 19904
rect 45235 19873 45247 19876
rect 45189 19867 45247 19873
rect 45554 19864 45560 19876
rect 45612 19864 45618 19916
rect 45649 19907 45707 19913
rect 45649 19873 45661 19907
rect 45695 19904 45707 19907
rect 46293 19907 46351 19913
rect 46293 19904 46305 19907
rect 45695 19876 46305 19904
rect 45695 19873 45707 19876
rect 45649 19867 45707 19873
rect 46293 19873 46305 19876
rect 46339 19873 46351 19907
rect 46293 19867 46351 19873
rect 46566 19864 46572 19916
rect 46624 19904 46630 19916
rect 47121 19907 47179 19913
rect 47121 19904 47133 19907
rect 46624 19876 47133 19904
rect 46624 19864 46630 19876
rect 47121 19873 47133 19876
rect 47167 19873 47179 19907
rect 47121 19867 47179 19873
rect 47596 19876 47900 19904
rect 25958 19836 25964 19848
rect 25919 19808 25964 19836
rect 25958 19796 25964 19808
rect 26016 19796 26022 19848
rect 26145 19839 26203 19845
rect 26145 19805 26157 19839
rect 26191 19836 26203 19839
rect 26418 19836 26424 19848
rect 26191 19808 26424 19836
rect 26191 19805 26203 19808
rect 26145 19799 26203 19805
rect 26418 19796 26424 19808
rect 26476 19796 26482 19848
rect 26602 19836 26608 19848
rect 26563 19808 26608 19836
rect 26602 19796 26608 19808
rect 26660 19796 26666 19848
rect 26789 19839 26847 19845
rect 26789 19805 26801 19839
rect 26835 19836 26847 19839
rect 27154 19836 27160 19848
rect 26835 19808 27160 19836
rect 26835 19805 26847 19808
rect 26789 19799 26847 19805
rect 27154 19796 27160 19808
rect 27212 19796 27218 19848
rect 27338 19796 27344 19848
rect 27396 19836 27402 19848
rect 27433 19839 27491 19845
rect 27433 19836 27445 19839
rect 27396 19808 27445 19836
rect 27396 19796 27402 19808
rect 27433 19805 27445 19808
rect 27479 19805 27491 19839
rect 27433 19799 27491 19805
rect 27522 19796 27528 19848
rect 27580 19836 27586 19848
rect 27617 19839 27675 19845
rect 27617 19836 27629 19839
rect 27580 19808 27629 19836
rect 27580 19796 27586 19808
rect 27617 19805 27629 19808
rect 27663 19805 27675 19839
rect 28810 19836 28816 19848
rect 28771 19808 28816 19836
rect 27617 19799 27675 19805
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 28994 19796 29000 19848
rect 29052 19836 29058 19848
rect 29549 19839 29607 19845
rect 29549 19836 29561 19839
rect 29052 19808 29561 19836
rect 29052 19796 29058 19808
rect 29549 19805 29561 19808
rect 29595 19805 29607 19839
rect 44266 19836 44272 19848
rect 44227 19808 44272 19836
rect 29549 19799 29607 19805
rect 44266 19796 44272 19808
rect 44324 19796 44330 19848
rect 44453 19839 44511 19845
rect 44453 19805 44465 19839
rect 44499 19805 44511 19839
rect 44453 19799 44511 19805
rect 24581 19771 24639 19777
rect 24581 19737 24593 19771
rect 24627 19737 24639 19771
rect 24581 19731 24639 19737
rect 28905 19771 28963 19777
rect 28905 19737 28917 19771
rect 28951 19768 28963 19771
rect 29733 19771 29791 19777
rect 29733 19768 29745 19771
rect 28951 19740 29745 19768
rect 28951 19737 28963 19740
rect 28905 19731 28963 19737
rect 29733 19737 29745 19740
rect 29779 19737 29791 19771
rect 31386 19768 31392 19780
rect 31347 19740 31392 19768
rect 29733 19731 29791 19737
rect 24596 19700 24624 19731
rect 31386 19728 31392 19740
rect 31444 19728 31450 19780
rect 44468 19768 44496 19799
rect 46014 19796 46020 19848
rect 46072 19836 46078 19848
rect 46382 19836 46388 19848
rect 46072 19808 46388 19836
rect 46072 19796 46078 19808
rect 46382 19796 46388 19808
rect 46440 19796 46446 19848
rect 47596 19836 47624 19876
rect 47872 19845 47900 19876
rect 46584 19808 47624 19836
rect 47673 19839 47731 19845
rect 46584 19780 46612 19808
rect 47673 19805 47685 19839
rect 47719 19805 47731 19839
rect 47673 19799 47731 19805
rect 47857 19839 47915 19845
rect 47857 19805 47869 19839
rect 47903 19805 47915 19839
rect 47857 19799 47915 19805
rect 46566 19768 46572 19780
rect 44468 19740 46572 19768
rect 46566 19728 46572 19740
rect 46624 19728 46630 19780
rect 23308 19672 24624 19700
rect 26145 19703 26203 19709
rect 26145 19669 26157 19703
rect 26191 19700 26203 19703
rect 26234 19700 26240 19712
rect 26191 19672 26240 19700
rect 26191 19669 26203 19672
rect 26145 19663 26203 19669
rect 26234 19660 26240 19672
rect 26292 19700 26298 19712
rect 27338 19700 27344 19712
rect 26292 19672 27344 19700
rect 26292 19660 26298 19672
rect 27338 19660 27344 19672
rect 27396 19660 27402 19712
rect 44266 19660 44272 19712
rect 44324 19700 44330 19712
rect 47688 19700 47716 19799
rect 44324 19672 47716 19700
rect 44324 19660 44330 19672
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 2406 19456 2412 19508
rect 2464 19496 2470 19508
rect 2464 19468 13124 19496
rect 2464 19456 2470 19468
rect 11238 19388 11244 19440
rect 11296 19428 11302 19440
rect 11793 19431 11851 19437
rect 11793 19428 11805 19431
rect 11296 19400 11805 19428
rect 11296 19388 11302 19400
rect 11793 19397 11805 19400
rect 11839 19397 11851 19431
rect 11793 19391 11851 19397
rect 12526 19388 12532 19440
rect 12584 19388 12590 19440
rect 13096 19428 13124 19468
rect 13170 19456 13176 19508
rect 13228 19496 13234 19508
rect 13265 19499 13323 19505
rect 13265 19496 13277 19499
rect 13228 19468 13277 19496
rect 13228 19456 13234 19468
rect 13265 19465 13277 19468
rect 13311 19465 13323 19499
rect 19978 19496 19984 19508
rect 13265 19459 13323 19465
rect 13372 19468 19984 19496
rect 13372 19428 13400 19468
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 21913 19499 21971 19505
rect 21913 19465 21925 19499
rect 21959 19496 21971 19499
rect 22186 19496 22192 19508
rect 21959 19468 22192 19496
rect 21959 19465 21971 19468
rect 21913 19459 21971 19465
rect 22186 19456 22192 19468
rect 22244 19456 22250 19508
rect 26510 19496 26516 19508
rect 26252 19468 26516 19496
rect 13906 19428 13912 19440
rect 13096 19400 13400 19428
rect 13867 19400 13912 19428
rect 13906 19388 13912 19400
rect 13964 19388 13970 19440
rect 14274 19428 14280 19440
rect 14235 19400 14280 19428
rect 14274 19388 14280 19400
rect 14332 19388 14338 19440
rect 16574 19388 16580 19440
rect 16632 19428 16638 19440
rect 17405 19431 17463 19437
rect 17405 19428 17417 19431
rect 16632 19400 17417 19428
rect 16632 19388 16638 19400
rect 17405 19397 17417 19400
rect 17451 19397 17463 19431
rect 20070 19428 20076 19440
rect 19918 19400 20076 19428
rect 17405 19391 17463 19397
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 20346 19388 20352 19440
rect 20404 19428 20410 19440
rect 26252 19428 26280 19468
rect 26510 19456 26516 19468
rect 26568 19456 26574 19508
rect 26602 19456 26608 19508
rect 26660 19496 26666 19508
rect 27249 19499 27307 19505
rect 27249 19496 27261 19499
rect 26660 19468 27261 19496
rect 26660 19456 26666 19468
rect 27249 19465 27261 19468
rect 27295 19465 27307 19499
rect 27249 19459 27307 19465
rect 27338 19456 27344 19508
rect 27396 19496 27402 19508
rect 27396 19468 27441 19496
rect 27396 19456 27402 19468
rect 29362 19456 29368 19508
rect 29420 19456 29426 19508
rect 44821 19499 44879 19505
rect 35866 19468 40264 19496
rect 20404 19400 26280 19428
rect 26329 19431 26387 19437
rect 20404 19388 20410 19400
rect 26329 19397 26341 19431
rect 26375 19428 26387 19431
rect 27522 19428 27528 19440
rect 26375 19400 27528 19428
rect 26375 19397 26387 19400
rect 26329 19391 26387 19397
rect 27522 19388 27528 19400
rect 27580 19388 27586 19440
rect 29380 19428 29408 19456
rect 29549 19431 29607 19437
rect 29549 19428 29561 19431
rect 29380 19400 29561 19428
rect 29549 19397 29561 19400
rect 29595 19397 29607 19431
rect 29549 19391 29607 19397
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 8846 19360 8852 19372
rect 8759 19332 8852 19360
rect 8846 19320 8852 19332
rect 8904 19360 8910 19372
rect 10594 19360 10600 19372
rect 8904 19332 10600 19360
rect 8904 19320 8910 19332
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19360 10931 19363
rect 11330 19360 11336 19372
rect 10919 19332 11336 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 14090 19360 14096 19372
rect 14051 19332 14096 19360
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 14182 19320 14188 19372
rect 14240 19360 14246 19372
rect 17129 19363 17187 19369
rect 14240 19332 14285 19360
rect 14240 19320 14246 19332
rect 17129 19329 17141 19363
rect 17175 19360 17187 19363
rect 17218 19360 17224 19372
rect 17175 19332 17224 19360
rect 17175 19329 17187 19332
rect 17129 19323 17187 19329
rect 17218 19320 17224 19332
rect 17276 19320 17282 19372
rect 18414 19360 18420 19372
rect 18375 19332 18420 19360
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 20717 19363 20775 19369
rect 20717 19329 20729 19363
rect 20763 19360 20775 19363
rect 20806 19360 20812 19372
rect 20763 19332 20812 19360
rect 20763 19329 20775 19332
rect 20717 19323 20775 19329
rect 20806 19320 20812 19332
rect 20864 19320 20870 19372
rect 20901 19363 20959 19369
rect 20901 19329 20913 19363
rect 20947 19360 20959 19363
rect 20990 19360 20996 19372
rect 20947 19332 20996 19360
rect 20947 19329 20959 19332
rect 20901 19323 20959 19329
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 21358 19320 21364 19372
rect 21416 19360 21422 19372
rect 22097 19363 22155 19369
rect 22097 19360 22109 19363
rect 21416 19332 22109 19360
rect 21416 19320 21422 19332
rect 22097 19329 22109 19332
rect 22143 19329 22155 19363
rect 22097 19323 22155 19329
rect 24578 19320 24584 19372
rect 24636 19360 24642 19372
rect 24636 19332 25912 19360
rect 24636 19320 24642 19332
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 8941 19295 8999 19301
rect 8941 19261 8953 19295
rect 8987 19261 8999 19295
rect 9214 19292 9220 19304
rect 9175 19264 9220 19292
rect 8941 19255 8999 19261
rect 8956 19224 8984 19255
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 10965 19295 11023 19301
rect 10965 19261 10977 19295
rect 11011 19292 11023 19295
rect 11517 19295 11575 19301
rect 11517 19292 11529 19295
rect 11011 19264 11529 19292
rect 11011 19261 11023 19264
rect 10965 19255 11023 19261
rect 11517 19261 11529 19264
rect 11563 19261 11575 19295
rect 11517 19255 11575 19261
rect 13722 19252 13728 19304
rect 13780 19292 13786 19304
rect 14461 19295 14519 19301
rect 14461 19292 14473 19295
rect 13780 19264 14473 19292
rect 13780 19252 13786 19264
rect 14461 19261 14473 19264
rect 14507 19261 14519 19295
rect 18690 19292 18696 19304
rect 18651 19264 18696 19292
rect 14461 19255 14519 19261
rect 18690 19252 18696 19264
rect 18748 19252 18754 19304
rect 18782 19252 18788 19304
rect 18840 19292 18846 19304
rect 19058 19292 19064 19304
rect 18840 19264 19064 19292
rect 18840 19252 18846 19264
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 19242 19252 19248 19304
rect 19300 19292 19306 19304
rect 24026 19292 24032 19304
rect 19300 19264 24032 19292
rect 19300 19252 19306 19264
rect 24026 19252 24032 19264
rect 24084 19252 24090 19304
rect 25884 19292 25912 19332
rect 25958 19320 25964 19372
rect 26016 19360 26022 19372
rect 26237 19363 26295 19369
rect 26237 19360 26249 19363
rect 26016 19332 26249 19360
rect 26016 19320 26022 19332
rect 26237 19329 26249 19332
rect 26283 19329 26295 19363
rect 26237 19323 26295 19329
rect 26418 19320 26424 19372
rect 26476 19360 26482 19372
rect 26970 19360 26976 19372
rect 26476 19332 26976 19360
rect 26476 19320 26482 19332
rect 26970 19320 26976 19332
rect 27028 19320 27034 19372
rect 27154 19360 27160 19372
rect 27115 19332 27160 19360
rect 27154 19320 27160 19332
rect 27212 19320 27218 19372
rect 27264 19332 29316 19360
rect 27264 19292 27292 19332
rect 25884 19264 27292 19292
rect 29288 19292 29316 19332
rect 29457 19295 29515 19301
rect 29457 19292 29469 19295
rect 29288 19264 29469 19292
rect 29457 19261 29469 19264
rect 29503 19261 29515 19295
rect 29457 19255 29515 19261
rect 30469 19295 30527 19301
rect 30469 19261 30481 19295
rect 30515 19292 30527 19295
rect 35866 19292 35894 19468
rect 39298 19428 39304 19440
rect 39259 19400 39304 19428
rect 39298 19388 39304 19400
rect 39356 19388 39362 19440
rect 40236 19437 40264 19468
rect 44821 19465 44833 19499
rect 44867 19496 44879 19499
rect 46842 19496 46848 19508
rect 44867 19468 46848 19496
rect 44867 19465 44879 19468
rect 44821 19459 44879 19465
rect 46842 19456 46848 19468
rect 46900 19456 46906 19508
rect 40221 19431 40279 19437
rect 40221 19397 40233 19431
rect 40267 19397 40279 19431
rect 47210 19428 47216 19440
rect 40221 19391 40279 19397
rect 45204 19400 47216 19428
rect 42794 19360 42800 19372
rect 40052 19332 42800 19360
rect 30515 19264 35894 19292
rect 39209 19295 39267 19301
rect 30515 19261 30527 19264
rect 30469 19255 30527 19261
rect 39209 19261 39221 19295
rect 39255 19292 39267 19295
rect 40052 19292 40080 19332
rect 42794 19320 42800 19332
rect 42852 19320 42858 19372
rect 45204 19369 45232 19400
rect 47210 19388 47216 19400
rect 47268 19388 47274 19440
rect 45189 19363 45247 19369
rect 45189 19329 45201 19363
rect 45235 19329 45247 19363
rect 45189 19323 45247 19329
rect 45281 19363 45339 19369
rect 45281 19329 45293 19363
rect 45327 19329 45339 19363
rect 46934 19360 46940 19372
rect 46690 19332 46940 19360
rect 45281 19323 45339 19329
rect 39255 19264 40080 19292
rect 39255 19261 39267 19264
rect 39209 19255 39267 19261
rect 11422 19224 11428 19236
rect 8956 19196 11428 19224
rect 11422 19184 11428 19196
rect 11480 19184 11486 19236
rect 18414 19224 18420 19236
rect 15764 19196 18420 19224
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 15764 19156 15792 19196
rect 18414 19184 18420 19196
rect 18472 19184 18478 19236
rect 21082 19224 21088 19236
rect 20180 19196 21088 19224
rect 7616 19128 15792 19156
rect 7616 19116 7622 19128
rect 17310 19116 17316 19168
rect 17368 19156 17374 19168
rect 20180 19165 20208 19196
rect 21082 19184 21088 19196
rect 21140 19184 21146 19236
rect 26973 19227 27031 19233
rect 26973 19193 26985 19227
rect 27019 19224 27031 19227
rect 29362 19224 29368 19236
rect 27019 19196 29368 19224
rect 27019 19193 27031 19196
rect 26973 19187 27031 19193
rect 29362 19184 29368 19196
rect 29420 19184 29426 19236
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 17368 19128 20177 19156
rect 17368 19116 17374 19128
rect 20165 19125 20177 19128
rect 20211 19125 20223 19159
rect 20806 19156 20812 19168
rect 20767 19128 20812 19156
rect 20165 19119 20223 19125
rect 20806 19116 20812 19128
rect 20864 19116 20870 19168
rect 26878 19116 26884 19168
rect 26936 19156 26942 19168
rect 30484 19156 30512 19255
rect 30558 19184 30564 19236
rect 30616 19224 30622 19236
rect 45296 19224 45324 19323
rect 46934 19320 46940 19332
rect 46992 19320 46998 19372
rect 47486 19320 47492 19372
rect 47544 19360 47550 19372
rect 47581 19363 47639 19369
rect 47581 19360 47593 19363
rect 47544 19332 47593 19360
rect 47544 19320 47550 19332
rect 47581 19329 47593 19332
rect 47627 19360 47639 19363
rect 47762 19360 47768 19372
rect 47627 19332 47768 19360
rect 47627 19329 47639 19332
rect 47581 19323 47639 19329
rect 47762 19320 47768 19332
rect 47820 19320 47826 19372
rect 45465 19295 45523 19301
rect 45465 19261 45477 19295
rect 45511 19292 45523 19295
rect 46014 19292 46020 19304
rect 45511 19264 46020 19292
rect 45511 19261 45523 19264
rect 45465 19255 45523 19261
rect 46014 19252 46020 19264
rect 46072 19252 46078 19304
rect 46201 19295 46259 19301
rect 46201 19261 46213 19295
rect 46247 19261 46259 19295
rect 47026 19292 47032 19304
rect 46987 19264 47032 19292
rect 46201 19255 46259 19261
rect 46216 19224 46244 19255
rect 47026 19252 47032 19264
rect 47084 19252 47090 19304
rect 30616 19196 46244 19224
rect 30616 19184 30622 19196
rect 47670 19156 47676 19168
rect 26936 19128 30512 19156
rect 47631 19128 47676 19156
rect 26936 19116 26942 19128
rect 47670 19116 47676 19128
rect 47728 19116 47734 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 2225 18915 2283 18921
rect 4890 18912 4896 18964
rect 4948 18912 4954 18964
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 12621 18955 12679 18961
rect 12621 18952 12633 18955
rect 12584 18924 12633 18952
rect 12584 18912 12590 18924
rect 12621 18921 12633 18924
rect 12667 18921 12679 18955
rect 12621 18915 12679 18921
rect 14182 18912 14188 18964
rect 14240 18952 14246 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 14240 18924 14289 18952
rect 14240 18912 14246 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 14458 18952 14464 18964
rect 14419 18924 14464 18952
rect 14277 18915 14335 18921
rect 14458 18912 14464 18924
rect 14516 18912 14522 18964
rect 15194 18912 15200 18964
rect 15252 18952 15258 18964
rect 17865 18955 17923 18961
rect 17865 18952 17877 18955
rect 15252 18924 17877 18952
rect 15252 18912 15258 18924
rect 17865 18921 17877 18924
rect 17911 18921 17923 18955
rect 17865 18915 17923 18921
rect 18509 18955 18567 18961
rect 18509 18921 18521 18955
rect 18555 18952 18567 18955
rect 18690 18952 18696 18964
rect 18555 18924 18696 18952
rect 18555 18921 18567 18924
rect 18509 18915 18567 18921
rect 18690 18912 18696 18924
rect 18748 18912 18754 18964
rect 26421 18955 26479 18961
rect 20916 18924 22094 18952
rect 4908 18884 4936 18912
rect 20916 18884 20944 18924
rect 4908 18856 20944 18884
rect 4890 18776 4896 18828
rect 4948 18816 4954 18828
rect 9401 18819 9459 18825
rect 9401 18816 9413 18819
rect 4948 18788 9413 18816
rect 4948 18776 4954 18788
rect 9401 18785 9413 18788
rect 9447 18785 9459 18819
rect 13354 18816 13360 18828
rect 9401 18779 9459 18785
rect 12544 18788 13360 18816
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 8202 18748 8208 18760
rect 8163 18720 8208 18748
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 8846 18708 8852 18760
rect 8904 18748 8910 18760
rect 12544 18757 12572 18788
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 15194 18776 15200 18828
rect 15252 18816 15258 18828
rect 19242 18816 19248 18828
rect 15252 18788 15516 18816
rect 15252 18776 15258 18788
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8904 18720 8953 18748
rect 8904 18708 8910 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 12529 18751 12587 18757
rect 12529 18717 12541 18751
rect 12575 18717 12587 18751
rect 12529 18711 12587 18717
rect 13078 18708 13084 18760
rect 13136 18748 13142 18760
rect 13173 18751 13231 18757
rect 13173 18748 13185 18751
rect 13136 18720 13185 18748
rect 13136 18708 13142 18720
rect 13173 18717 13185 18720
rect 13219 18717 13231 18751
rect 15378 18748 15384 18760
rect 15339 18720 15384 18748
rect 13173 18711 13231 18717
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 15488 18757 15516 18788
rect 17512 18788 19248 18816
rect 17512 18757 17540 18788
rect 19242 18776 19248 18788
rect 19300 18776 19306 18828
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 19978 18816 19984 18828
rect 19484 18788 19984 18816
rect 19484 18776 19490 18788
rect 19978 18776 19984 18788
rect 20036 18776 20042 18828
rect 20714 18816 20720 18828
rect 20675 18788 20720 18816
rect 20714 18776 20720 18788
rect 20772 18776 20778 18828
rect 20993 18819 21051 18825
rect 20993 18785 21005 18819
rect 21039 18816 21051 18819
rect 21082 18816 21088 18828
rect 21039 18788 21088 18816
rect 21039 18785 21051 18788
rect 20993 18779 21051 18785
rect 21082 18776 21088 18788
rect 21140 18776 21146 18828
rect 22066 18816 22094 18924
rect 26421 18921 26433 18955
rect 26467 18952 26479 18955
rect 27154 18952 27160 18964
rect 26467 18924 27160 18952
rect 26467 18921 26479 18924
rect 26421 18915 26479 18921
rect 27154 18912 27160 18924
rect 27212 18912 27218 18964
rect 26252 18856 27108 18884
rect 26252 18825 26280 18856
rect 26237 18819 26295 18825
rect 26237 18816 26249 18819
rect 22066 18788 26249 18816
rect 26237 18785 26249 18788
rect 26283 18785 26295 18819
rect 26237 18779 26295 18785
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18717 18751 18751
rect 18693 18711 18751 18717
rect 8297 18683 8355 18689
rect 8297 18649 8309 18683
rect 8343 18680 8355 18683
rect 9125 18683 9183 18689
rect 9125 18680 9137 18683
rect 8343 18652 9137 18680
rect 8343 18649 8355 18652
rect 8297 18643 8355 18649
rect 9125 18649 9137 18652
rect 9171 18649 9183 18683
rect 14090 18680 14096 18692
rect 14003 18652 14096 18680
rect 9125 18643 9183 18649
rect 14090 18640 14096 18652
rect 14148 18680 14154 18692
rect 14642 18680 14648 18692
rect 14148 18652 14648 18680
rect 14148 18640 14154 18652
rect 14642 18640 14648 18652
rect 14700 18640 14706 18692
rect 17310 18680 17316 18692
rect 17271 18652 17316 18680
rect 17310 18640 17316 18652
rect 17368 18640 17374 18692
rect 17589 18683 17647 18689
rect 17589 18649 17601 18683
rect 17635 18680 17647 18683
rect 18230 18680 18236 18692
rect 17635 18652 18236 18680
rect 17635 18649 17647 18652
rect 17589 18643 17647 18649
rect 18230 18640 18236 18652
rect 18288 18640 18294 18692
rect 18708 18680 18736 18711
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 19392 18720 19533 18748
rect 19392 18708 19398 18720
rect 19521 18717 19533 18720
rect 19567 18748 19579 18751
rect 20809 18751 20867 18757
rect 20809 18748 20821 18751
rect 19567 18720 20821 18748
rect 19567 18717 19579 18720
rect 19521 18711 19579 18717
rect 20809 18717 20821 18720
rect 20855 18717 20867 18751
rect 20809 18711 20867 18717
rect 19426 18680 19432 18692
rect 18708 18652 19432 18680
rect 19426 18640 19432 18652
rect 19484 18640 19490 18692
rect 12894 18572 12900 18624
rect 12952 18612 12958 18624
rect 13265 18615 13323 18621
rect 13265 18612 13277 18615
rect 12952 18584 13277 18612
rect 12952 18572 12958 18584
rect 13265 18581 13277 18584
rect 13311 18581 13323 18615
rect 13265 18575 13323 18581
rect 14274 18572 14280 18624
rect 14332 18621 14338 18624
rect 14332 18615 14361 18621
rect 14349 18612 14361 18615
rect 15657 18615 15715 18621
rect 15657 18612 15669 18615
rect 14349 18584 15669 18612
rect 14349 18581 14361 18584
rect 14332 18575 14361 18581
rect 15657 18581 15669 18584
rect 15703 18581 15715 18615
rect 15657 18575 15715 18581
rect 14332 18572 14338 18575
rect 17678 18572 17684 18624
rect 17736 18612 17742 18624
rect 20530 18612 20536 18624
rect 17736 18584 17781 18612
rect 20491 18584 20536 18612
rect 17736 18572 17742 18584
rect 20530 18572 20536 18584
rect 20588 18572 20594 18624
rect 20824 18612 20852 18711
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 20956 18720 21001 18748
rect 20956 18708 20962 18720
rect 22002 18708 22008 18760
rect 22060 18750 22066 18760
rect 22281 18751 22339 18757
rect 22060 18748 22094 18750
rect 22281 18748 22293 18751
rect 22060 18720 22293 18748
rect 22060 18708 22066 18720
rect 22281 18717 22293 18720
rect 22327 18748 22339 18751
rect 22833 18751 22891 18757
rect 22833 18748 22845 18751
rect 22327 18720 22845 18748
rect 22327 18717 22339 18720
rect 22281 18711 22339 18717
rect 22833 18717 22845 18720
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18748 23719 18751
rect 24397 18751 24455 18757
rect 24397 18748 24409 18751
rect 23707 18720 24409 18748
rect 23707 18717 23719 18720
rect 23661 18711 23719 18717
rect 24397 18717 24409 18720
rect 24443 18748 24455 18751
rect 25038 18748 25044 18760
rect 24443 18720 25044 18748
rect 24443 18717 24455 18720
rect 24397 18711 24455 18717
rect 25038 18708 25044 18720
rect 25096 18708 25102 18760
rect 25961 18751 26019 18757
rect 25961 18717 25973 18751
rect 26007 18717 26019 18751
rect 25961 18711 26019 18717
rect 25976 18680 26004 18711
rect 26050 18708 26056 18760
rect 26108 18748 26114 18760
rect 26329 18751 26387 18757
rect 26108 18720 26153 18748
rect 26108 18708 26114 18720
rect 26329 18717 26341 18751
rect 26375 18748 26387 18751
rect 26878 18748 26884 18760
rect 26375 18720 26884 18748
rect 26375 18717 26387 18720
rect 26329 18711 26387 18717
rect 26878 18708 26884 18720
rect 26936 18708 26942 18760
rect 27080 18757 27108 18856
rect 46477 18819 46535 18825
rect 46477 18785 46489 18819
rect 46523 18816 46535 18819
rect 47670 18816 47676 18828
rect 46523 18788 47676 18816
rect 46523 18785 46535 18788
rect 46477 18779 46535 18785
rect 47670 18776 47676 18788
rect 47728 18776 47734 18828
rect 48130 18816 48136 18828
rect 48091 18788 48136 18816
rect 48130 18776 48136 18788
rect 48188 18776 48194 18828
rect 27065 18751 27123 18757
rect 27065 18717 27077 18751
rect 27111 18748 27123 18751
rect 27154 18748 27160 18760
rect 27111 18720 27160 18748
rect 27111 18717 27123 18720
rect 27065 18711 27123 18717
rect 27154 18708 27160 18720
rect 27212 18708 27218 18760
rect 27614 18708 27620 18760
rect 27672 18748 27678 18760
rect 45833 18751 45891 18757
rect 27672 18720 28488 18748
rect 27672 18708 27678 18720
rect 27249 18683 27307 18689
rect 25976 18652 26280 18680
rect 26252 18624 26280 18652
rect 27249 18649 27261 18683
rect 27295 18680 27307 18683
rect 27798 18680 27804 18692
rect 27295 18652 27804 18680
rect 27295 18649 27307 18652
rect 27249 18643 27307 18649
rect 27798 18640 27804 18652
rect 27856 18640 27862 18692
rect 28074 18680 28080 18692
rect 28035 18652 28080 18680
rect 28074 18640 28080 18652
rect 28132 18640 28138 18692
rect 28460 18689 28488 18720
rect 45833 18717 45845 18751
rect 45879 18748 45891 18751
rect 46293 18751 46351 18757
rect 46293 18748 46305 18751
rect 45879 18720 46305 18748
rect 45879 18717 45891 18720
rect 45833 18711 45891 18717
rect 46293 18717 46305 18720
rect 46339 18717 46351 18751
rect 46293 18711 46351 18717
rect 28445 18683 28503 18689
rect 28445 18649 28457 18683
rect 28491 18680 28503 18683
rect 29546 18680 29552 18692
rect 28491 18652 29552 18680
rect 28491 18649 28503 18652
rect 28445 18643 28503 18649
rect 29546 18640 29552 18652
rect 29604 18640 29610 18692
rect 20990 18612 20996 18624
rect 20824 18584 20996 18612
rect 20990 18572 20996 18584
rect 21048 18572 21054 18624
rect 22278 18612 22284 18624
rect 22239 18584 22284 18612
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 22462 18572 22468 18624
rect 22520 18612 22526 18624
rect 23017 18615 23075 18621
rect 23017 18612 23029 18615
rect 22520 18584 23029 18612
rect 22520 18572 22526 18584
rect 23017 18581 23029 18584
rect 23063 18581 23075 18615
rect 23017 18575 23075 18581
rect 23566 18572 23572 18624
rect 23624 18612 23630 18624
rect 23753 18615 23811 18621
rect 23753 18612 23765 18615
rect 23624 18584 23765 18612
rect 23624 18572 23630 18584
rect 23753 18581 23765 18584
rect 23799 18581 23811 18615
rect 24486 18612 24492 18624
rect 24447 18584 24492 18612
rect 23753 18575 23811 18581
rect 24486 18572 24492 18584
rect 24544 18572 24550 18624
rect 26234 18572 26240 18624
rect 26292 18572 26298 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1949 18411 2007 18417
rect 1949 18377 1961 18411
rect 1995 18408 2007 18411
rect 7558 18408 7564 18420
rect 1995 18380 7564 18408
rect 1995 18377 2007 18380
rect 1949 18371 2007 18377
rect 7558 18368 7564 18380
rect 7616 18368 7622 18420
rect 12406 18380 28028 18408
rect 2130 18300 2136 18352
rect 2188 18340 2194 18352
rect 6638 18340 6644 18352
rect 2188 18312 6644 18340
rect 2188 18300 2194 18312
rect 6638 18300 6644 18312
rect 6696 18340 6702 18352
rect 12406 18340 12434 18380
rect 6696 18312 12434 18340
rect 6696 18300 6702 18312
rect 13906 18300 13912 18352
rect 13964 18300 13970 18352
rect 14458 18300 14464 18352
rect 14516 18340 14522 18352
rect 16025 18343 16083 18349
rect 14516 18312 15332 18340
rect 14516 18300 14522 18312
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 12894 18272 12900 18284
rect 12855 18244 12900 18272
rect 12894 18232 12900 18244
rect 12952 18232 12958 18284
rect 15102 18272 15108 18284
rect 15063 18244 15108 18272
rect 15102 18232 15108 18244
rect 15160 18232 15166 18284
rect 15304 18281 15332 18312
rect 16025 18309 16037 18343
rect 16071 18340 16083 18343
rect 16853 18343 16911 18349
rect 16853 18340 16865 18343
rect 16071 18312 16865 18340
rect 16071 18309 16083 18312
rect 16025 18303 16083 18309
rect 16853 18309 16865 18312
rect 16899 18309 16911 18343
rect 16853 18303 16911 18309
rect 17310 18300 17316 18352
rect 17368 18340 17374 18352
rect 18969 18343 19027 18349
rect 18969 18340 18981 18343
rect 17368 18312 18981 18340
rect 17368 18300 17374 18312
rect 18969 18309 18981 18312
rect 19015 18309 19027 18343
rect 19334 18340 19340 18352
rect 19295 18312 19340 18340
rect 18969 18303 19027 18309
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 20070 18340 20076 18352
rect 20031 18312 20076 18340
rect 20070 18300 20076 18312
rect 20128 18300 20134 18352
rect 24486 18340 24492 18352
rect 23966 18312 24492 18340
rect 24486 18300 24492 18312
rect 24544 18300 24550 18352
rect 26145 18343 26203 18349
rect 26145 18340 26157 18343
rect 25608 18312 26157 18340
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18241 15347 18275
rect 15289 18235 15347 18241
rect 15654 18232 15660 18284
rect 15712 18272 15718 18284
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15712 18244 15945 18272
rect 15712 18232 15718 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 16114 18232 16120 18284
rect 16172 18272 16178 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16172 18244 16681 18272
rect 16172 18232 16178 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19153 18275 19211 18281
rect 19153 18272 19165 18275
rect 19116 18244 19165 18272
rect 19116 18232 19122 18244
rect 19153 18241 19165 18244
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 13173 18207 13231 18213
rect 13173 18173 13185 18207
rect 13219 18204 13231 18207
rect 18509 18207 18567 18213
rect 13219 18176 15148 18204
rect 13219 18173 13231 18176
rect 13173 18167 13231 18173
rect 15120 18145 15148 18176
rect 18509 18173 18521 18207
rect 18555 18204 18567 18207
rect 18782 18204 18788 18216
rect 18555 18176 18788 18204
rect 18555 18173 18567 18176
rect 18509 18167 18567 18173
rect 18782 18164 18788 18176
rect 18840 18164 18846 18216
rect 19168 18204 19196 18235
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 19981 18275 20039 18281
rect 19300 18244 19345 18272
rect 19300 18232 19306 18244
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 20162 18272 20168 18284
rect 20027 18244 20168 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20898 18272 20904 18284
rect 20272 18244 20904 18272
rect 20272 18204 20300 18244
rect 20898 18232 20904 18244
rect 20956 18232 20962 18284
rect 22462 18272 22468 18284
rect 22423 18244 22468 18272
rect 22462 18232 22468 18244
rect 22520 18232 22526 18284
rect 25608 18281 25636 18312
rect 26145 18309 26157 18312
rect 26191 18340 26203 18343
rect 26602 18340 26608 18352
rect 26191 18312 26608 18340
rect 26191 18309 26203 18312
rect 26145 18303 26203 18309
rect 26602 18300 26608 18312
rect 26660 18300 26666 18352
rect 26878 18300 26884 18352
rect 26936 18340 26942 18352
rect 26973 18343 27031 18349
rect 26973 18340 26985 18343
rect 26936 18312 26985 18340
rect 26936 18300 26942 18312
rect 26973 18309 26985 18312
rect 27019 18309 27031 18343
rect 27154 18340 27160 18352
rect 27115 18312 27160 18340
rect 26973 18303 27031 18309
rect 27154 18300 27160 18312
rect 27212 18300 27218 18352
rect 28000 18340 28028 18380
rect 28074 18368 28080 18420
rect 28132 18408 28138 18420
rect 28169 18411 28227 18417
rect 28169 18408 28181 18411
rect 28132 18380 28181 18408
rect 28132 18368 28138 18380
rect 28169 18377 28181 18380
rect 28215 18377 28227 18411
rect 46934 18408 46940 18420
rect 46895 18380 46940 18408
rect 28169 18371 28227 18377
rect 46934 18368 46940 18380
rect 46992 18368 46998 18420
rect 47949 18343 48007 18349
rect 47949 18340 47961 18343
rect 28000 18312 28672 18340
rect 25409 18275 25467 18281
rect 25409 18241 25421 18275
rect 25455 18241 25467 18275
rect 25409 18235 25467 18241
rect 25593 18275 25651 18281
rect 25593 18241 25605 18275
rect 25639 18241 25651 18275
rect 26050 18272 26056 18284
rect 26011 18244 26056 18272
rect 25593 18235 25651 18241
rect 20806 18204 20812 18216
rect 19168 18176 20300 18204
rect 20767 18176 20812 18204
rect 20806 18164 20812 18176
rect 20864 18164 20870 18216
rect 15105 18139 15163 18145
rect 15105 18105 15117 18139
rect 15151 18105 15163 18139
rect 15105 18099 15163 18105
rect 14642 18068 14648 18080
rect 14603 18040 14648 18068
rect 14642 18028 14648 18040
rect 14700 18028 14706 18080
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 18138 18068 18144 18080
rect 15436 18040 18144 18068
rect 15436 18028 15442 18040
rect 18138 18028 18144 18040
rect 18196 18068 18202 18080
rect 19334 18068 19340 18080
rect 18196 18040 19340 18068
rect 18196 18028 18202 18040
rect 19334 18028 19340 18040
rect 19392 18028 19398 18080
rect 19518 18068 19524 18080
rect 19479 18040 19524 18068
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 20916 18068 20944 18232
rect 22741 18207 22799 18213
rect 22741 18204 22753 18207
rect 22572 18176 22753 18204
rect 21269 18139 21327 18145
rect 21269 18105 21281 18139
rect 21315 18136 21327 18139
rect 22572 18136 22600 18176
rect 22741 18173 22753 18176
rect 22787 18173 22799 18207
rect 22741 18167 22799 18173
rect 24489 18207 24547 18213
rect 24489 18173 24501 18207
rect 24535 18204 24547 18207
rect 25424 18204 25452 18235
rect 26050 18232 26056 18244
rect 26108 18232 26114 18284
rect 26234 18272 26240 18284
rect 26195 18244 26240 18272
rect 26234 18232 26240 18244
rect 26292 18232 26298 18284
rect 28644 18281 28672 18312
rect 46860 18312 47961 18340
rect 46860 18284 46888 18312
rect 47949 18309 47961 18312
rect 47995 18309 48007 18343
rect 47949 18303 48007 18309
rect 27341 18275 27399 18281
rect 27341 18241 27353 18275
rect 27387 18272 27399 18275
rect 27985 18275 28043 18281
rect 27985 18272 27997 18275
rect 27387 18244 27997 18272
rect 27387 18241 27399 18244
rect 27341 18235 27399 18241
rect 27985 18241 27997 18244
rect 28031 18241 28043 18275
rect 27985 18235 28043 18241
rect 28629 18275 28687 18281
rect 28629 18241 28641 18275
rect 28675 18272 28687 18275
rect 32766 18272 32772 18284
rect 28675 18244 32772 18272
rect 28675 18241 28687 18244
rect 28629 18235 28687 18241
rect 32766 18232 32772 18244
rect 32824 18232 32830 18284
rect 46842 18272 46848 18284
rect 46803 18244 46848 18272
rect 46842 18232 46848 18244
rect 46900 18232 46906 18284
rect 47029 18275 47087 18281
rect 47029 18241 47041 18275
rect 47075 18272 47087 18275
rect 47210 18272 47216 18284
rect 47075 18244 47216 18272
rect 47075 18241 47087 18244
rect 47029 18235 47087 18241
rect 47210 18232 47216 18244
rect 47268 18232 47274 18284
rect 47486 18232 47492 18284
rect 47544 18272 47550 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 47544 18244 47593 18272
rect 47544 18232 47550 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47762 18272 47768 18284
rect 47723 18244 47768 18272
rect 47581 18235 47639 18241
rect 47762 18232 47768 18244
rect 47820 18232 47826 18284
rect 26418 18204 26424 18216
rect 24535 18176 25360 18204
rect 25424 18176 26424 18204
rect 24535 18173 24547 18176
rect 24489 18167 24547 18173
rect 21315 18108 22600 18136
rect 21315 18105 21327 18108
rect 21269 18099 21327 18105
rect 24504 18068 24532 18167
rect 20916 18040 24532 18068
rect 25332 18068 25360 18176
rect 26418 18164 26424 18176
rect 26476 18164 26482 18216
rect 27798 18204 27804 18216
rect 27711 18176 27804 18204
rect 27798 18164 27804 18176
rect 27856 18204 27862 18216
rect 28074 18204 28080 18216
rect 27856 18176 28080 18204
rect 27856 18164 27862 18176
rect 28074 18164 28080 18176
rect 28132 18164 28138 18216
rect 25501 18139 25559 18145
rect 25501 18105 25513 18139
rect 25547 18136 25559 18139
rect 27430 18136 27436 18148
rect 25547 18108 27436 18136
rect 25547 18105 25559 18108
rect 25501 18099 25559 18105
rect 27430 18096 27436 18108
rect 27488 18096 27494 18148
rect 28994 18136 29000 18148
rect 27540 18108 29000 18136
rect 27540 18068 27568 18108
rect 28994 18096 29000 18108
rect 29052 18096 29058 18148
rect 28718 18068 28724 18080
rect 25332 18040 27568 18068
rect 28679 18040 28724 18068
rect 28718 18028 28724 18040
rect 28776 18028 28782 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 14093 17867 14151 17873
rect 14093 17833 14105 17867
rect 14139 17864 14151 17867
rect 15102 17864 15108 17876
rect 14139 17836 15108 17864
rect 14139 17833 14151 17836
rect 14093 17827 14151 17833
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 19426 17824 19432 17876
rect 19484 17864 19490 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 19484 17836 19717 17864
rect 19484 17824 19490 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 21358 17864 21364 17876
rect 21319 17836 21364 17864
rect 19705 17827 19763 17833
rect 21358 17824 21364 17836
rect 21416 17824 21422 17876
rect 23753 17867 23811 17873
rect 23753 17833 23765 17867
rect 23799 17864 23811 17867
rect 24026 17864 24032 17876
rect 23799 17836 24032 17864
rect 23799 17833 23811 17836
rect 23753 17827 23811 17833
rect 24026 17824 24032 17836
rect 24084 17824 24090 17876
rect 26418 17864 26424 17876
rect 26379 17836 26424 17864
rect 26418 17824 26424 17836
rect 26476 17824 26482 17876
rect 47210 17824 47216 17876
rect 47268 17864 47274 17876
rect 47489 17867 47547 17873
rect 47489 17864 47501 17867
rect 47268 17836 47501 17864
rect 47268 17824 47274 17836
rect 47489 17833 47501 17836
rect 47535 17833 47547 17867
rect 47489 17827 47547 17833
rect 19613 17799 19671 17805
rect 19613 17765 19625 17799
rect 19659 17796 19671 17799
rect 20530 17796 20536 17808
rect 19659 17768 20536 17796
rect 19659 17765 19671 17768
rect 19613 17759 19671 17765
rect 20530 17756 20536 17768
rect 20588 17756 20594 17808
rect 46753 17799 46811 17805
rect 46753 17765 46765 17799
rect 46799 17796 46811 17799
rect 46799 17768 47624 17796
rect 46799 17765 46811 17768
rect 46753 17759 46811 17765
rect 3970 17688 3976 17740
rect 4028 17728 4034 17740
rect 11885 17731 11943 17737
rect 11885 17728 11897 17731
rect 4028 17700 11897 17728
rect 4028 17688 4034 17700
rect 11885 17697 11897 17700
rect 11931 17697 11943 17731
rect 14642 17728 14648 17740
rect 11885 17691 11943 17697
rect 14108 17700 14648 17728
rect 14108 17669 14136 17700
rect 14642 17688 14648 17700
rect 14700 17728 14706 17740
rect 15381 17731 15439 17737
rect 15381 17728 15393 17731
rect 14700 17700 15393 17728
rect 14700 17688 14706 17700
rect 15381 17697 15393 17700
rect 15427 17697 15439 17731
rect 15381 17691 15439 17697
rect 17862 17688 17868 17740
rect 17920 17728 17926 17740
rect 18417 17731 18475 17737
rect 18417 17728 18429 17731
rect 17920 17700 18429 17728
rect 17920 17688 17926 17700
rect 18417 17697 18429 17700
rect 18463 17697 18475 17731
rect 18417 17691 18475 17697
rect 19245 17731 19303 17737
rect 19245 17697 19257 17731
rect 19291 17728 19303 17731
rect 19334 17728 19340 17740
rect 19291 17700 19340 17728
rect 19291 17697 19303 17700
rect 19245 17691 19303 17697
rect 19334 17688 19340 17700
rect 19392 17728 19398 17740
rect 19518 17728 19524 17740
rect 19392 17700 19524 17728
rect 19392 17688 19398 17700
rect 19518 17688 19524 17700
rect 19576 17688 19582 17740
rect 20806 17688 20812 17740
rect 20864 17728 20870 17740
rect 20993 17731 21051 17737
rect 20993 17728 21005 17731
rect 20864 17700 21005 17728
rect 20864 17688 20870 17700
rect 20993 17697 21005 17700
rect 21039 17697 21051 17731
rect 20993 17691 21051 17697
rect 22005 17731 22063 17737
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22278 17728 22284 17740
rect 22051 17700 22284 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 22278 17688 22284 17700
rect 22336 17688 22342 17740
rect 11425 17663 11483 17669
rect 11425 17629 11437 17663
rect 11471 17629 11483 17663
rect 11425 17623 11483 17629
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17629 14151 17663
rect 14366 17660 14372 17672
rect 14327 17632 14372 17660
rect 14093 17623 14151 17629
rect 11440 17524 11468 17623
rect 14366 17620 14372 17632
rect 14424 17620 14430 17672
rect 18230 17660 18236 17672
rect 18191 17632 18236 17660
rect 18230 17620 18236 17632
rect 18288 17620 18294 17672
rect 20349 17663 20407 17669
rect 20349 17660 20361 17663
rect 19260 17632 20361 17660
rect 19260 17604 19288 17632
rect 20349 17629 20361 17632
rect 20395 17629 20407 17663
rect 20349 17623 20407 17629
rect 21177 17663 21235 17669
rect 21177 17629 21189 17663
rect 21223 17629 21235 17663
rect 21177 17623 21235 17629
rect 11609 17595 11667 17601
rect 11609 17561 11621 17595
rect 11655 17592 11667 17595
rect 11698 17592 11704 17604
rect 11655 17564 11704 17592
rect 11655 17561 11667 17564
rect 11609 17555 11667 17561
rect 11698 17552 11704 17564
rect 11756 17552 11762 17604
rect 15194 17552 15200 17604
rect 15252 17592 15258 17604
rect 15565 17595 15623 17601
rect 15565 17592 15577 17595
rect 15252 17564 15577 17592
rect 15252 17552 15258 17564
rect 15565 17561 15577 17564
rect 15611 17561 15623 17595
rect 17218 17592 17224 17604
rect 17179 17564 17224 17592
rect 15565 17555 15623 17561
rect 17218 17552 17224 17564
rect 17276 17552 17282 17604
rect 17770 17552 17776 17604
rect 17828 17592 17834 17604
rect 17865 17595 17923 17601
rect 17865 17592 17877 17595
rect 17828 17564 17877 17592
rect 17828 17552 17834 17564
rect 17865 17561 17877 17564
rect 17911 17561 17923 17595
rect 17865 17555 17923 17561
rect 18049 17595 18107 17601
rect 18049 17561 18061 17595
rect 18095 17592 18107 17595
rect 19242 17592 19248 17604
rect 18095 17564 19248 17592
rect 18095 17561 18107 17564
rect 18049 17555 18107 17561
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 20165 17595 20223 17601
rect 20165 17561 20177 17595
rect 20211 17561 20223 17595
rect 20165 17555 20223 17561
rect 20533 17595 20591 17601
rect 20533 17561 20545 17595
rect 20579 17592 20591 17595
rect 21192 17592 21220 17623
rect 27430 17620 27436 17672
rect 27488 17660 27494 17672
rect 27617 17663 27675 17669
rect 27617 17660 27629 17663
rect 27488 17632 27629 17660
rect 27488 17620 27494 17632
rect 27617 17629 27629 17632
rect 27663 17629 27675 17663
rect 28074 17660 28080 17672
rect 28035 17632 28080 17660
rect 27617 17623 27675 17629
rect 28074 17620 28080 17632
rect 28132 17620 28138 17672
rect 46937 17663 46995 17669
rect 46937 17629 46949 17663
rect 46983 17660 46995 17663
rect 47026 17660 47032 17672
rect 46983 17632 47032 17660
rect 46983 17629 46995 17632
rect 46937 17623 46995 17629
rect 47026 17620 47032 17632
rect 47084 17620 47090 17672
rect 47596 17669 47624 17768
rect 47397 17663 47455 17669
rect 47397 17629 47409 17663
rect 47443 17629 47455 17663
rect 47397 17623 47455 17629
rect 47581 17663 47639 17669
rect 47581 17629 47593 17663
rect 47627 17660 47639 17663
rect 47762 17660 47768 17672
rect 47627 17632 47768 17660
rect 47627 17629 47639 17632
rect 47581 17623 47639 17629
rect 20579 17564 21220 17592
rect 20579 17561 20591 17564
rect 20533 17555 20591 17561
rect 11974 17524 11980 17536
rect 11440 17496 11980 17524
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 14182 17484 14188 17536
rect 14240 17524 14246 17536
rect 14277 17527 14335 17533
rect 14277 17524 14289 17527
rect 14240 17496 14289 17524
rect 14240 17484 14246 17496
rect 14277 17493 14289 17496
rect 14323 17493 14335 17527
rect 18138 17524 18144 17536
rect 18099 17496 18144 17524
rect 14277 17487 14335 17493
rect 18138 17484 18144 17496
rect 18196 17524 18202 17536
rect 20180 17524 20208 17555
rect 22186 17552 22192 17604
rect 22244 17592 22250 17604
rect 22281 17595 22339 17601
rect 22281 17592 22293 17595
rect 22244 17564 22293 17592
rect 22244 17552 22250 17564
rect 22281 17561 22293 17564
rect 22327 17561 22339 17595
rect 23566 17592 23572 17604
rect 23506 17564 23572 17592
rect 22281 17555 22339 17561
rect 23566 17552 23572 17564
rect 23624 17552 23630 17604
rect 25682 17552 25688 17604
rect 25740 17592 25746 17604
rect 26050 17592 26056 17604
rect 25740 17564 26056 17592
rect 25740 17552 25746 17564
rect 26050 17552 26056 17564
rect 26108 17552 26114 17604
rect 26234 17592 26240 17604
rect 26195 17564 26240 17592
rect 26234 17552 26240 17564
rect 26292 17552 26298 17604
rect 27706 17552 27712 17604
rect 27764 17592 27770 17604
rect 47412 17592 47440 17623
rect 47762 17620 47768 17632
rect 47820 17620 47826 17672
rect 47486 17592 47492 17604
rect 27764 17564 27922 17592
rect 47399 17564 47492 17592
rect 27764 17552 27770 17564
rect 47486 17552 47492 17564
rect 47544 17592 47550 17604
rect 48038 17592 48044 17604
rect 47544 17564 48044 17592
rect 47544 17552 47550 17564
rect 48038 17552 48044 17564
rect 48096 17552 48102 17604
rect 18196 17496 20208 17524
rect 18196 17484 18202 17496
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 11698 17320 11704 17332
rect 11659 17292 11704 17320
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 13906 17280 13912 17332
rect 13964 17320 13970 17332
rect 14001 17323 14059 17329
rect 14001 17320 14013 17323
rect 13964 17292 14013 17320
rect 13964 17280 13970 17292
rect 14001 17289 14013 17292
rect 14047 17289 14059 17323
rect 15194 17320 15200 17332
rect 15155 17292 15200 17320
rect 14001 17283 14059 17289
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 18443 17323 18501 17329
rect 18443 17289 18455 17323
rect 18489 17320 18501 17323
rect 19058 17320 19064 17332
rect 18489 17292 19064 17320
rect 18489 17289 18501 17292
rect 18443 17283 18501 17289
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 19978 17280 19984 17332
rect 20036 17320 20042 17332
rect 22002 17320 22008 17332
rect 20036 17292 22008 17320
rect 20036 17280 20042 17292
rect 22002 17280 22008 17292
rect 22060 17280 22066 17332
rect 8021 17255 8079 17261
rect 8021 17221 8033 17255
rect 8067 17252 8079 17255
rect 8757 17255 8815 17261
rect 8757 17252 8769 17255
rect 8067 17224 8769 17252
rect 8067 17221 8079 17224
rect 8021 17215 8079 17221
rect 8757 17221 8769 17224
rect 8803 17221 8815 17255
rect 17310 17252 17316 17264
rect 8757 17215 8815 17221
rect 10244 17224 17316 17252
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17184 7987 17187
rect 8202 17184 8208 17196
rect 7975 17156 8208 17184
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 8202 17144 8208 17156
rect 8260 17144 8266 17196
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 10244 17116 10272 17224
rect 17310 17212 17316 17224
rect 17368 17252 17374 17264
rect 17770 17252 17776 17264
rect 17368 17224 17776 17252
rect 17368 17212 17374 17224
rect 17770 17212 17776 17224
rect 17828 17212 17834 17264
rect 18138 17212 18144 17264
rect 18196 17252 18202 17264
rect 18233 17255 18291 17261
rect 18233 17252 18245 17255
rect 18196 17224 18245 17252
rect 18196 17212 18202 17224
rect 18233 17221 18245 17224
rect 18279 17221 18291 17255
rect 18233 17215 18291 17221
rect 27893 17255 27951 17261
rect 27893 17221 27905 17255
rect 27939 17252 27951 17255
rect 28718 17252 28724 17264
rect 27939 17224 28724 17252
rect 27939 17221 27951 17224
rect 27893 17215 27951 17221
rect 28718 17212 28724 17224
rect 28776 17212 28782 17264
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 11606 17184 11612 17196
rect 11112 17156 11612 17184
rect 11112 17144 11118 17156
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 12406 17156 12572 17184
rect 10410 17116 10416 17128
rect 8619 17088 10272 17116
rect 10371 17088 10416 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 10410 17076 10416 17088
rect 10468 17076 10474 17128
rect 8202 17008 8208 17060
rect 8260 17048 8266 17060
rect 12406 17048 12434 17156
rect 12544 17116 12572 17156
rect 13354 17144 13360 17196
rect 13412 17184 13418 17196
rect 13909 17187 13967 17193
rect 13909 17184 13921 17187
rect 13412 17156 13921 17184
rect 13412 17144 13418 17156
rect 13909 17153 13921 17156
rect 13955 17184 13967 17187
rect 14826 17184 14832 17196
rect 13955 17156 14832 17184
rect 13955 17153 13967 17156
rect 13909 17147 13967 17153
rect 14826 17144 14832 17156
rect 14884 17144 14890 17196
rect 15105 17187 15163 17193
rect 15105 17184 15117 17187
rect 14936 17156 15117 17184
rect 14936 17116 14964 17156
rect 15105 17153 15117 17156
rect 15151 17184 15163 17187
rect 15151 17156 15516 17184
rect 15151 17153 15163 17156
rect 15105 17147 15163 17153
rect 12544 17088 14964 17116
rect 15488 17116 15516 17156
rect 15654 17144 15660 17196
rect 15712 17184 15718 17196
rect 15749 17187 15807 17193
rect 15749 17184 15761 17187
rect 15712 17156 15761 17184
rect 15712 17144 15718 17156
rect 15749 17153 15761 17156
rect 15795 17153 15807 17187
rect 15749 17147 15807 17153
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17184 19855 17187
rect 19978 17184 19984 17196
rect 19843 17156 19984 17184
rect 19843 17153 19855 17156
rect 19797 17147 19855 17153
rect 19978 17144 19984 17156
rect 20036 17144 20042 17196
rect 21818 17184 21824 17196
rect 21779 17156 21824 17184
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 47578 17184 47584 17196
rect 47539 17156 47584 17184
rect 47578 17144 47584 17156
rect 47636 17144 47642 17196
rect 16574 17116 16580 17128
rect 15488 17088 16580 17116
rect 16574 17076 16580 17088
rect 16632 17076 16638 17128
rect 27706 17116 27712 17128
rect 27667 17088 27712 17116
rect 27706 17076 27712 17088
rect 27764 17076 27770 17128
rect 28166 17116 28172 17128
rect 28127 17088 28172 17116
rect 28166 17076 28172 17088
rect 28224 17076 28230 17128
rect 8260 17020 12434 17048
rect 8260 17008 8266 17020
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 18601 17051 18659 17057
rect 18601 17048 18613 17051
rect 18288 17020 18613 17048
rect 18288 17008 18294 17020
rect 18601 17017 18613 17020
rect 18647 17017 18659 17051
rect 18601 17011 18659 17017
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 1452 16952 2053 16980
rect 1452 16940 1458 16952
rect 2041 16949 2053 16952
rect 2087 16949 2099 16983
rect 2041 16943 2099 16949
rect 11606 16940 11612 16992
rect 11664 16980 11670 16992
rect 15654 16980 15660 16992
rect 11664 16952 15660 16980
rect 11664 16940 11670 16952
rect 15654 16940 15660 16952
rect 15712 16940 15718 16992
rect 15746 16940 15752 16992
rect 15804 16980 15810 16992
rect 15841 16983 15899 16989
rect 15841 16980 15853 16983
rect 15804 16952 15853 16980
rect 15804 16940 15810 16952
rect 15841 16949 15853 16952
rect 15887 16949 15899 16983
rect 15841 16943 15899 16949
rect 18417 16983 18475 16989
rect 18417 16949 18429 16983
rect 18463 16980 18475 16983
rect 18506 16980 18512 16992
rect 18463 16952 18512 16980
rect 18463 16949 18475 16952
rect 18417 16943 18475 16949
rect 18506 16940 18512 16952
rect 18564 16940 18570 16992
rect 19426 16940 19432 16992
rect 19484 16980 19490 16992
rect 19613 16983 19671 16989
rect 19613 16980 19625 16983
rect 19484 16952 19625 16980
rect 19484 16940 19490 16952
rect 19613 16949 19625 16952
rect 19659 16949 19671 16983
rect 19613 16943 19671 16949
rect 46290 16940 46296 16992
rect 46348 16980 46354 16992
rect 47029 16983 47087 16989
rect 47029 16980 47041 16983
rect 46348 16952 47041 16980
rect 46348 16940 46354 16952
rect 47029 16949 47041 16952
rect 47075 16949 47087 16983
rect 47670 16980 47676 16992
rect 47631 16952 47676 16980
rect 47029 16943 47087 16949
rect 47670 16940 47676 16952
rect 47728 16940 47734 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 28166 16776 28172 16788
rect 3384 16748 28172 16776
rect 3384 16736 3390 16748
rect 28166 16736 28172 16748
rect 28224 16736 28230 16788
rect 18046 16668 18052 16720
rect 18104 16708 18110 16720
rect 18322 16708 18328 16720
rect 18104 16680 18328 16708
rect 18104 16668 18110 16680
rect 18322 16668 18328 16680
rect 18380 16668 18386 16720
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 15746 16640 15752 16652
rect 15707 16612 15752 16640
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 19334 16640 19340 16652
rect 18432 16612 19340 16640
rect 15102 16532 15108 16584
rect 15160 16572 15166 16584
rect 15565 16575 15623 16581
rect 15565 16572 15577 16575
rect 15160 16544 15577 16572
rect 15160 16532 15166 16544
rect 15565 16541 15577 16544
rect 15611 16541 15623 16575
rect 15565 16535 15623 16541
rect 17218 16532 17224 16584
rect 17276 16572 17282 16584
rect 18432 16581 18460 16612
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16640 19855 16643
rect 19978 16640 19984 16652
rect 19843 16612 19984 16640
rect 19843 16609 19855 16612
rect 19797 16603 19855 16609
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 46290 16640 46296 16652
rect 46251 16612 46296 16640
rect 46290 16600 46296 16612
rect 46348 16600 46354 16652
rect 48130 16640 48136 16652
rect 48091 16612 48136 16640
rect 48130 16600 48136 16612
rect 48188 16600 48194 16652
rect 18417 16575 18475 16581
rect 17276 16544 18368 16572
rect 17276 16532 17282 16544
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 2130 16504 2136 16516
rect 1627 16476 2136 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 17405 16507 17463 16513
rect 17405 16473 17417 16507
rect 17451 16504 17463 16507
rect 17494 16504 17500 16516
rect 17451 16476 17500 16504
rect 17451 16473 17463 16476
rect 17405 16467 17463 16473
rect 17494 16464 17500 16476
rect 17552 16464 17558 16516
rect 18138 16504 18144 16516
rect 18099 16476 18144 16504
rect 18138 16464 18144 16476
rect 18196 16464 18202 16516
rect 18340 16504 18368 16544
rect 18417 16541 18429 16575
rect 18463 16541 18475 16575
rect 18417 16535 18475 16541
rect 18506 16532 18512 16584
rect 18564 16572 18570 16584
rect 19242 16572 19248 16584
rect 18564 16544 19248 16572
rect 18564 16532 18570 16544
rect 19242 16532 19248 16544
rect 19300 16572 19306 16584
rect 19429 16575 19487 16581
rect 19429 16572 19441 16575
rect 19300 16544 19441 16572
rect 19300 16532 19306 16544
rect 19429 16541 19441 16544
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 20272 16544 22094 16572
rect 20272 16504 20300 16544
rect 18340 16476 20300 16504
rect 20349 16507 20407 16513
rect 20349 16473 20361 16507
rect 20395 16504 20407 16507
rect 21818 16504 21824 16516
rect 20395 16476 21824 16504
rect 20395 16473 20407 16476
rect 20349 16467 20407 16473
rect 21818 16464 21824 16476
rect 21876 16464 21882 16516
rect 17954 16396 17960 16448
rect 18012 16436 18018 16448
rect 18239 16439 18297 16445
rect 18239 16436 18251 16439
rect 18012 16408 18251 16436
rect 18012 16396 18018 16408
rect 18239 16405 18251 16408
rect 18285 16405 18297 16439
rect 18239 16399 18297 16405
rect 18325 16439 18383 16445
rect 18325 16405 18337 16439
rect 18371 16436 18383 16439
rect 18506 16436 18512 16448
rect 18371 16408 18512 16436
rect 18371 16405 18383 16408
rect 18325 16399 18383 16405
rect 18506 16396 18512 16408
rect 18564 16396 18570 16448
rect 20438 16436 20444 16448
rect 20399 16408 20444 16436
rect 20438 16396 20444 16408
rect 20496 16396 20502 16448
rect 22066 16436 22094 16544
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 47670 16504 47676 16516
rect 46523 16476 47676 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 47670 16464 47676 16476
rect 47728 16464 47734 16516
rect 45554 16436 45560 16448
rect 22066 16408 45560 16436
rect 45554 16396 45560 16408
rect 45612 16396 45618 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 14182 16232 14188 16244
rect 12728 16204 14188 16232
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16096 2102 16108
rect 12728 16105 12756 16204
rect 14182 16192 14188 16204
rect 14240 16232 14246 16244
rect 15102 16232 15108 16244
rect 14240 16204 15108 16232
rect 14240 16192 14246 16204
rect 15102 16192 15108 16204
rect 15160 16232 15166 16244
rect 15289 16235 15347 16241
rect 15289 16232 15301 16235
rect 15160 16204 15301 16232
rect 15160 16192 15166 16204
rect 15289 16201 15301 16204
rect 15335 16201 15347 16235
rect 15289 16195 15347 16201
rect 18138 16192 18144 16244
rect 18196 16232 18202 16244
rect 18969 16235 19027 16241
rect 18969 16232 18981 16235
rect 18196 16204 18981 16232
rect 18196 16192 18202 16204
rect 18969 16201 18981 16204
rect 19015 16201 19027 16235
rect 18969 16195 19027 16201
rect 19242 16192 19248 16244
rect 19300 16232 19306 16244
rect 21177 16235 21235 16241
rect 21177 16232 21189 16235
rect 19300 16204 21189 16232
rect 19300 16192 19306 16204
rect 21177 16201 21189 16204
rect 21223 16201 21235 16235
rect 21177 16195 21235 16201
rect 19705 16167 19763 16173
rect 19705 16133 19717 16167
rect 19751 16164 19763 16167
rect 19978 16164 19984 16176
rect 19751 16136 19984 16164
rect 19751 16133 19763 16136
rect 19705 16127 19763 16133
rect 19978 16124 19984 16136
rect 20036 16124 20042 16176
rect 12713 16099 12771 16105
rect 2096 16068 2774 16096
rect 2096 16056 2102 16068
rect 2746 15892 2774 16068
rect 12713 16065 12725 16099
rect 12759 16065 12771 16099
rect 12713 16059 12771 16065
rect 14918 16056 14924 16108
rect 14976 16056 14982 16108
rect 18598 16056 18604 16108
rect 18656 16056 18662 16108
rect 19426 16096 19432 16108
rect 19387 16068 19432 16096
rect 19426 16056 19432 16068
rect 19484 16056 19490 16108
rect 20806 16056 20812 16108
rect 20864 16056 20870 16108
rect 47118 16056 47124 16108
rect 47176 16096 47182 16108
rect 47581 16099 47639 16105
rect 47581 16096 47593 16099
rect 47176 16068 47593 16096
rect 47176 16056 47182 16068
rect 47581 16065 47593 16068
rect 47627 16065 47639 16099
rect 47581 16059 47639 16065
rect 12805 16031 12863 16037
rect 12805 15997 12817 16031
rect 12851 15997 12863 16031
rect 13538 16028 13544 16040
rect 13499 16000 13544 16028
rect 12805 15991 12863 15997
rect 12710 15892 12716 15904
rect 2746 15864 12716 15892
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 12820 15892 12848 15991
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 13817 16031 13875 16037
rect 13817 16028 13829 16031
rect 13648 16000 13829 16028
rect 13081 15963 13139 15969
rect 13081 15929 13093 15963
rect 13127 15960 13139 15963
rect 13648 15960 13676 16000
rect 13817 15997 13829 16000
rect 13863 15997 13875 16031
rect 17218 16028 17224 16040
rect 17179 16000 17224 16028
rect 13817 15991 13875 15997
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 17497 16031 17555 16037
rect 17497 15997 17509 16031
rect 17543 16028 17555 16031
rect 18046 16028 18052 16040
rect 17543 16000 18052 16028
rect 17543 15997 17555 16000
rect 17497 15991 17555 15997
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 18966 15988 18972 16040
rect 19024 16028 19030 16040
rect 28810 16028 28816 16040
rect 19024 16000 28816 16028
rect 19024 15988 19030 16000
rect 28810 15988 28816 16000
rect 28868 15988 28874 16040
rect 13127 15932 13676 15960
rect 13127 15929 13139 15932
rect 13081 15923 13139 15929
rect 14366 15892 14372 15904
rect 12820 15864 14372 15892
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 46290 15852 46296 15904
rect 46348 15892 46354 15904
rect 47029 15895 47087 15901
rect 47029 15892 47041 15895
rect 46348 15864 47041 15892
rect 46348 15852 46354 15864
rect 47029 15861 47041 15864
rect 47075 15861 47087 15895
rect 47670 15892 47676 15904
rect 47631 15864 47676 15892
rect 47029 15855 47087 15861
rect 47670 15852 47676 15864
rect 47728 15852 47734 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 13538 15648 13544 15700
rect 13596 15688 13602 15700
rect 14093 15691 14151 15697
rect 14093 15688 14105 15691
rect 13596 15660 14105 15688
rect 13596 15648 13602 15660
rect 14093 15657 14105 15660
rect 14139 15657 14151 15691
rect 14918 15688 14924 15700
rect 14879 15660 14924 15688
rect 14093 15651 14151 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 18598 15648 18604 15700
rect 18656 15688 18662 15700
rect 19337 15691 19395 15697
rect 19337 15688 19349 15691
rect 18656 15660 19349 15688
rect 18656 15648 18662 15660
rect 19337 15657 19349 15660
rect 19383 15657 19395 15691
rect 19337 15651 19395 15657
rect 20625 15691 20683 15697
rect 20625 15657 20637 15691
rect 20671 15688 20683 15691
rect 20806 15688 20812 15700
rect 20671 15660 20812 15688
rect 20671 15657 20683 15660
rect 20625 15651 20683 15657
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 12710 15580 12716 15632
rect 12768 15620 12774 15632
rect 18874 15620 18880 15632
rect 12768 15592 18880 15620
rect 12768 15580 12774 15592
rect 18874 15580 18880 15592
rect 18932 15580 18938 15632
rect 16393 15555 16451 15561
rect 16393 15521 16405 15555
rect 16439 15552 16451 15555
rect 18138 15552 18144 15564
rect 16439 15524 18144 15552
rect 16439 15521 16451 15524
rect 16393 15515 16451 15521
rect 18138 15512 18144 15524
rect 18196 15512 18202 15564
rect 46290 15552 46296 15564
rect 46251 15524 46296 15552
rect 46290 15512 46296 15524
rect 46348 15512 46354 15564
rect 46477 15555 46535 15561
rect 46477 15521 46489 15555
rect 46523 15552 46535 15555
rect 47670 15552 47676 15564
rect 46523 15524 47676 15552
rect 46523 15521 46535 15524
rect 46477 15515 46535 15521
rect 47670 15512 47676 15524
rect 47728 15512 47734 15564
rect 48130 15552 48136 15564
rect 48091 15524 48136 15552
rect 48130 15512 48136 15524
rect 48188 15512 48194 15564
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 14274 15484 14280 15496
rect 14235 15456 14280 15484
rect 2041 15447 2099 15453
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 14826 15484 14832 15496
rect 14787 15456 14832 15484
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15453 15807 15487
rect 19242 15484 19248 15496
rect 19155 15456 19248 15484
rect 15749 15447 15807 15453
rect 15764 15348 15792 15447
rect 19242 15444 19248 15456
rect 19300 15484 19306 15496
rect 20162 15484 20168 15496
rect 19300 15456 20168 15484
rect 19300 15444 19306 15456
rect 20162 15444 20168 15456
rect 20220 15484 20226 15496
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 20220 15456 20545 15484
rect 20220 15444 20226 15456
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 15841 15419 15899 15425
rect 15841 15385 15853 15419
rect 15887 15416 15899 15419
rect 16577 15419 16635 15425
rect 16577 15416 16589 15419
rect 15887 15388 16589 15416
rect 15887 15385 15899 15388
rect 15841 15379 15899 15385
rect 16577 15385 16589 15388
rect 16623 15385 16635 15419
rect 16577 15379 16635 15385
rect 18138 15376 18144 15428
rect 18196 15416 18202 15428
rect 18233 15419 18291 15425
rect 18233 15416 18245 15419
rect 18196 15388 18245 15416
rect 18196 15376 18202 15388
rect 18233 15385 18245 15388
rect 18279 15385 18291 15419
rect 18233 15379 18291 15385
rect 16298 15348 16304 15360
rect 15764 15320 16304 15348
rect 16298 15308 16304 15320
rect 16356 15348 16362 15360
rect 18966 15348 18972 15360
rect 16356 15320 18972 15348
rect 16356 15308 16362 15320
rect 18966 15308 18972 15320
rect 19024 15308 19030 15360
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 17218 15104 17224 15156
rect 17276 15144 17282 15156
rect 17405 15147 17463 15153
rect 17405 15144 17417 15147
rect 17276 15116 17417 15144
rect 17276 15104 17282 15116
rect 17405 15113 17417 15116
rect 17451 15113 17463 15147
rect 18046 15144 18052 15156
rect 18007 15116 18052 15144
rect 17405 15107 17463 15113
rect 18046 15104 18052 15116
rect 18104 15104 18110 15156
rect 17862 15036 17868 15088
rect 17920 15076 17926 15088
rect 17920 15048 18184 15076
rect 17920 15036 17926 15048
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 14826 15008 14832 15020
rect 14787 14980 14832 15008
rect 14826 14968 14832 14980
rect 14884 14968 14890 15020
rect 17405 15011 17463 15017
rect 17405 14977 17417 15011
rect 17451 15008 17463 15011
rect 17770 15008 17776 15020
rect 17451 14980 17776 15008
rect 17451 14977 17463 14980
rect 17405 14971 17463 14977
rect 17770 14968 17776 14980
rect 17828 14968 17834 15020
rect 17954 15008 17960 15020
rect 17915 14980 17960 15008
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 18156 15017 18184 15048
rect 18141 15011 18199 15017
rect 18141 14977 18153 15011
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 2832 14912 2877 14940
rect 2832 14900 2838 14912
rect 14921 14807 14979 14813
rect 14921 14773 14933 14807
rect 14967 14804 14979 14807
rect 15010 14804 15016 14816
rect 14967 14776 15016 14804
rect 14967 14773 14979 14776
rect 14921 14767 14979 14773
rect 15010 14764 15016 14776
rect 15068 14764 15074 14816
rect 17218 14764 17224 14816
rect 17276 14804 17282 14816
rect 17586 14804 17592 14816
rect 17276 14776 17592 14804
rect 17276 14764 17282 14776
rect 17586 14764 17592 14776
rect 17644 14764 17650 14816
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 17310 14560 17316 14612
rect 17368 14600 17374 14612
rect 17405 14603 17463 14609
rect 17405 14600 17417 14603
rect 17368 14572 17417 14600
rect 17368 14560 17374 14572
rect 17405 14569 17417 14572
rect 17451 14569 17463 14603
rect 17405 14563 17463 14569
rect 17218 14532 17224 14544
rect 2746 14504 17224 14532
rect 2746 14408 2774 14504
rect 17218 14492 17224 14504
rect 17276 14492 17282 14544
rect 17589 14535 17647 14541
rect 17589 14501 17601 14535
rect 17635 14501 17647 14535
rect 17589 14495 17647 14501
rect 17604 14464 17632 14495
rect 15672 14436 17632 14464
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2682 14396 2688 14408
rect 2179 14368 2688 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2682 14356 2688 14368
rect 2740 14368 2774 14408
rect 14274 14396 14280 14408
rect 14187 14368 14280 14396
rect 2740 14356 2746 14368
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 15672 14405 15700 14436
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 20438 14464 20444 14476
rect 17828 14436 20444 14464
rect 17828 14424 17834 14436
rect 15381 14399 15439 14405
rect 15381 14396 15393 14399
rect 14424 14368 15393 14396
rect 14424 14356 14430 14368
rect 15381 14365 15393 14368
rect 15427 14365 15439 14399
rect 15381 14359 15439 14365
rect 15657 14399 15715 14405
rect 15657 14365 15669 14399
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14396 15899 14399
rect 16022 14396 16028 14408
rect 15887 14368 16028 14396
rect 15887 14365 15899 14368
rect 15841 14359 15899 14365
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16298 14396 16304 14408
rect 16259 14368 16304 14396
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 17788 14396 17816 14424
rect 18248 14405 18276 14436
rect 20438 14424 20444 14436
rect 20496 14424 20502 14476
rect 16408 14368 17816 14396
rect 18233 14399 18291 14405
rect 14292 14328 14320 14356
rect 16408 14328 16436 14368
rect 18233 14365 18245 14399
rect 18279 14365 18291 14399
rect 19242 14396 19248 14408
rect 19203 14368 19248 14396
rect 18233 14359 18291 14365
rect 19242 14356 19248 14368
rect 19300 14356 19306 14408
rect 17218 14328 17224 14340
rect 14292 14300 16436 14328
rect 17179 14300 17224 14328
rect 17218 14288 17224 14300
rect 17276 14288 17282 14340
rect 17437 14331 17495 14337
rect 17437 14297 17449 14331
rect 17483 14328 17495 14331
rect 17862 14328 17868 14340
rect 17483 14300 17868 14328
rect 17483 14297 17495 14300
rect 17437 14291 17495 14297
rect 17862 14288 17868 14300
rect 17920 14288 17926 14340
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 14461 14263 14519 14269
rect 14461 14260 14473 14263
rect 14332 14232 14473 14260
rect 14332 14220 14338 14232
rect 14461 14229 14473 14232
rect 14507 14229 14519 14263
rect 15194 14260 15200 14272
rect 15155 14232 15200 14260
rect 14461 14223 14519 14229
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 15838 14220 15844 14272
rect 15896 14260 15902 14272
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 15896 14232 16405 14260
rect 15896 14220 15902 14232
rect 16393 14229 16405 14232
rect 16439 14229 16451 14263
rect 16393 14223 16451 14229
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 18233 14263 18291 14269
rect 18233 14260 18245 14263
rect 18012 14232 18245 14260
rect 18012 14220 18018 14232
rect 18233 14229 18245 14232
rect 18279 14229 18291 14263
rect 18233 14223 18291 14229
rect 19337 14263 19395 14269
rect 19337 14229 19349 14263
rect 19383 14260 19395 14263
rect 19426 14260 19432 14272
rect 19383 14232 19432 14260
rect 19383 14229 19395 14232
rect 19337 14223 19395 14229
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 16022 14056 16028 14068
rect 15935 14028 16028 14056
rect 16022 14016 16028 14028
rect 16080 14016 16086 14068
rect 17405 14059 17463 14065
rect 17405 14025 17417 14059
rect 17451 14056 17463 14059
rect 17678 14056 17684 14068
rect 17451 14028 17684 14056
rect 17451 14025 17463 14028
rect 17405 14019 17463 14025
rect 17678 14016 17684 14028
rect 17736 14016 17742 14068
rect 20809 14059 20867 14065
rect 20809 14056 20821 14059
rect 18248 14028 20821 14056
rect 15010 13948 15016 14000
rect 15068 13948 15074 14000
rect 16040 13988 16068 14016
rect 17310 13997 17316 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 16040 13960 17049 13988
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17253 13991 17316 13997
rect 17253 13988 17265 13991
rect 17223 13960 17265 13988
rect 17037 13951 17095 13957
rect 17253 13957 17265 13960
rect 17299 13957 17316 13991
rect 17253 13951 17316 13957
rect 17310 13948 17316 13951
rect 17368 13988 17374 14000
rect 18248 13988 18276 14028
rect 20809 14025 20821 14028
rect 20855 14025 20867 14059
rect 20809 14019 20867 14025
rect 19337 13991 19395 13997
rect 19337 13988 19349 13991
rect 17368 13960 18276 13988
rect 17368 13948 17374 13960
rect 14274 13920 14280 13932
rect 14235 13892 14280 13920
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 18248 13929 18276 13960
rect 18984 13960 19349 13988
rect 18233 13923 18291 13929
rect 18233 13889 18245 13923
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 18141 13855 18199 13861
rect 18141 13852 18153 13855
rect 17920 13824 18153 13852
rect 17920 13812 17926 13824
rect 18141 13821 18153 13824
rect 18187 13821 18199 13855
rect 18141 13815 18199 13821
rect 18601 13855 18659 13861
rect 18601 13821 18613 13855
rect 18647 13852 18659 13855
rect 18984 13852 19012 13960
rect 19337 13957 19349 13960
rect 19383 13957 19395 13991
rect 19337 13951 19395 13957
rect 20070 13948 20076 14000
rect 20128 13948 20134 14000
rect 47118 13880 47124 13932
rect 47176 13920 47182 13932
rect 47581 13923 47639 13929
rect 47581 13920 47593 13923
rect 47176 13892 47593 13920
rect 47176 13880 47182 13892
rect 47581 13889 47593 13892
rect 47627 13889 47639 13923
rect 47581 13883 47639 13889
rect 18647 13824 19012 13852
rect 19061 13855 19119 13861
rect 18647 13821 18659 13824
rect 18601 13815 18659 13821
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 19334 13852 19340 13864
rect 19107 13824 19340 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4614 13716 4620 13728
rect 4028 13688 4620 13716
rect 4028 13676 4034 13688
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 14540 13719 14598 13725
rect 14540 13685 14552 13719
rect 14586 13716 14598 13719
rect 15194 13716 15200 13728
rect 14586 13688 15200 13716
rect 14586 13685 14598 13688
rect 14540 13679 14598 13685
rect 15194 13676 15200 13688
rect 15252 13676 15258 13728
rect 17218 13716 17224 13728
rect 17179 13688 17224 13716
rect 17218 13676 17224 13688
rect 17276 13676 17282 13728
rect 47670 13716 47676 13728
rect 47631 13688 47676 13716
rect 47670 13676 47676 13688
rect 47728 13676 47734 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12492 13484 16160 13512
rect 12492 13472 12498 13484
rect 16022 13444 16028 13456
rect 15672 13416 16028 13444
rect 15672 13385 15700 13416
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13345 15715 13379
rect 15838 13376 15844 13388
rect 15799 13348 15844 13376
rect 15657 13339 15715 13345
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 16132 13385 16160 13484
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19392 13484 19441 13512
rect 19392 13472 19398 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 19429 13475 19487 13481
rect 20070 13472 20076 13524
rect 20128 13512 20134 13524
rect 20165 13515 20223 13521
rect 20165 13512 20177 13515
rect 20128 13484 20177 13512
rect 20128 13472 20134 13484
rect 20165 13481 20177 13484
rect 20211 13481 20223 13515
rect 20165 13475 20223 13481
rect 19242 13404 19248 13456
rect 19300 13404 19306 13456
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 17402 13336 17408 13388
rect 17460 13376 17466 13388
rect 18049 13379 18107 13385
rect 18049 13376 18061 13379
rect 17460 13348 18061 13376
rect 17460 13336 17466 13348
rect 18049 13345 18061 13348
rect 18095 13345 18107 13379
rect 19260 13376 19288 13404
rect 46477 13379 46535 13385
rect 19260 13348 20116 13376
rect 18049 13339 18107 13345
rect 17218 13268 17224 13320
rect 17276 13308 17282 13320
rect 18141 13311 18199 13317
rect 18141 13308 18153 13311
rect 17276 13280 18153 13308
rect 17276 13268 17282 13280
rect 18141 13277 18153 13280
rect 18187 13308 18199 13311
rect 18230 13308 18236 13320
rect 18187 13280 18236 13308
rect 18187 13277 18199 13280
rect 18141 13271 18199 13277
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 20088 13317 20116 13348
rect 46477 13345 46489 13379
rect 46523 13376 46535 13379
rect 47670 13376 47676 13388
rect 46523 13348 47676 13376
rect 46523 13345 46535 13348
rect 46477 13339 46535 13345
rect 47670 13336 47676 13348
rect 47728 13336 47734 13388
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 20073 13311 20131 13317
rect 20073 13277 20085 13311
rect 20119 13277 20131 13311
rect 46290 13308 46296 13320
rect 46251 13280 46296 13308
rect 20073 13271 20131 13277
rect 16850 13200 16856 13252
rect 16908 13240 16914 13252
rect 17236 13240 17264 13268
rect 16908 13212 17264 13240
rect 19444 13240 19472 13271
rect 46290 13268 46296 13280
rect 46348 13268 46354 13320
rect 20438 13240 20444 13252
rect 19444 13212 20444 13240
rect 16908 13200 16914 13212
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 48130 13240 48136 13252
rect 48091 13212 48136 13240
rect 48130 13200 48136 13212
rect 48188 13200 48194 13252
rect 18138 13132 18144 13184
rect 18196 13172 18202 13184
rect 18509 13175 18567 13181
rect 18509 13172 18521 13175
rect 18196 13144 18521 13172
rect 18196 13132 18202 13144
rect 18509 13141 18521 13144
rect 18555 13141 18567 13175
rect 18509 13135 18567 13141
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 17402 12968 17408 12980
rect 1627 12940 2774 12968
rect 17363 12940 17408 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 2746 12696 2774 12940
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 17862 12928 17868 12980
rect 17920 12928 17926 12980
rect 18230 12928 18236 12980
rect 18288 12968 18294 12980
rect 19613 12971 19671 12977
rect 19613 12968 19625 12971
rect 18288 12940 19625 12968
rect 18288 12928 18294 12940
rect 19613 12937 19625 12940
rect 19659 12937 19671 12971
rect 19613 12931 19671 12937
rect 17880 12900 17908 12928
rect 18138 12900 18144 12912
rect 17236 12872 17908 12900
rect 18099 12872 18144 12900
rect 17236 12841 17264 12872
rect 18138 12860 18144 12872
rect 18196 12860 18202 12912
rect 19426 12900 19432 12912
rect 19366 12872 19432 12900
rect 19426 12860 19432 12872
rect 19484 12860 19490 12912
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 17368 12804 17417 12832
rect 17368 12792 17374 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17862 12832 17868 12844
rect 17823 12804 17868 12832
rect 17405 12795 17463 12801
rect 17862 12792 17868 12804
rect 17920 12792 17926 12844
rect 46290 12792 46296 12844
rect 46348 12832 46354 12844
rect 47765 12835 47823 12841
rect 47765 12832 47777 12835
rect 46348 12804 47777 12832
rect 46348 12792 46354 12804
rect 47765 12801 47777 12804
rect 47811 12801 47823 12835
rect 47765 12795 47823 12801
rect 25590 12764 25596 12776
rect 17972 12736 25596 12764
rect 17972 12696 18000 12736
rect 25590 12724 25596 12736
rect 25648 12724 25654 12776
rect 2746 12668 18000 12696
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 41598 12180 41604 12232
rect 41656 12220 41662 12232
rect 46753 12223 46811 12229
rect 46753 12220 46765 12223
rect 41656 12192 46765 12220
rect 41656 12180 41662 12192
rect 46753 12189 46765 12192
rect 46799 12189 46811 12223
rect 46753 12183 46811 12189
rect 46474 12044 46480 12096
rect 46532 12084 46538 12096
rect 46845 12087 46903 12093
rect 46845 12084 46857 12087
rect 46532 12056 46857 12084
rect 46532 12044 46538 12056
rect 46845 12053 46857 12056
rect 46891 12053 46903 12087
rect 46845 12047 46903 12053
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 20622 11880 20628 11892
rect 18012 11852 20628 11880
rect 18012 11840 18018 11852
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 16574 11772 16580 11824
rect 16632 11812 16638 11824
rect 18877 11815 18935 11821
rect 16632 11784 18828 11812
rect 16632 11772 16638 11784
rect 17773 11747 17831 11753
rect 17773 11713 17785 11747
rect 17819 11744 17831 11747
rect 17954 11744 17960 11756
rect 17819 11716 17960 11744
rect 17819 11713 17831 11716
rect 17773 11707 17831 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 18800 11753 18828 11784
rect 18877 11781 18889 11815
rect 18923 11812 18935 11815
rect 19613 11815 19671 11821
rect 19613 11812 19625 11815
rect 18923 11784 19625 11812
rect 18923 11781 18935 11784
rect 18877 11775 18935 11781
rect 19613 11781 19625 11784
rect 19659 11781 19671 11815
rect 19613 11775 19671 11781
rect 18785 11747 18843 11753
rect 18785 11713 18797 11747
rect 18831 11713 18843 11747
rect 18785 11707 18843 11713
rect 17310 11636 17316 11688
rect 17368 11676 17374 11688
rect 19429 11679 19487 11685
rect 19429 11676 19441 11679
rect 17368 11648 19441 11676
rect 17368 11636 17374 11648
rect 19429 11645 19441 11648
rect 19475 11645 19487 11679
rect 19429 11639 19487 11645
rect 21269 11679 21327 11685
rect 21269 11645 21281 11679
rect 21315 11676 21327 11679
rect 27614 11676 27620 11688
rect 21315 11648 27620 11676
rect 21315 11645 21327 11648
rect 21269 11639 21327 11645
rect 27614 11636 27620 11648
rect 27672 11636 27678 11688
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 17865 11543 17923 11549
rect 17865 11540 17877 11543
rect 17092 11512 17877 11540
rect 17092 11500 17098 11512
rect 17865 11509 17877 11512
rect 17911 11509 17923 11543
rect 17865 11503 17923 11509
rect 46290 11500 46296 11552
rect 46348 11540 46354 11552
rect 47765 11543 47823 11549
rect 47765 11540 47777 11543
rect 46348 11512 47777 11540
rect 46348 11500 46354 11512
rect 47765 11509 47777 11512
rect 47811 11509 47823 11543
rect 47765 11503 47823 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 14826 11228 14832 11280
rect 14884 11268 14890 11280
rect 14884 11240 17356 11268
rect 14884 11228 14890 11240
rect 16850 11200 16856 11212
rect 16811 11172 16856 11200
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 17034 11200 17040 11212
rect 16995 11172 17040 11200
rect 17034 11160 17040 11172
rect 17092 11160 17098 11212
rect 17328 11209 17356 11240
rect 17313 11203 17371 11209
rect 17313 11169 17325 11203
rect 17359 11169 17371 11203
rect 46290 11200 46296 11212
rect 46251 11172 46296 11200
rect 17313 11163 17371 11169
rect 46290 11160 46296 11172
rect 46348 11160 46354 11212
rect 46474 11200 46480 11212
rect 46435 11172 46480 11200
rect 46474 11160 46480 11172
rect 46532 11160 46538 11212
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 4890 10996 4896 11008
rect 2832 10968 4896 10996
rect 2832 10956 2838 10968
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 18506 10724 18512 10736
rect 17880 10696 18512 10724
rect 17880 10665 17908 10696
rect 18506 10684 18512 10696
rect 18564 10684 18570 10736
rect 46106 10724 46112 10736
rect 46067 10696 46112 10724
rect 46106 10684 46112 10696
rect 46164 10684 46170 10736
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18138 10588 18144 10600
rect 18095 10560 18144 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 18325 10591 18383 10597
rect 18325 10557 18337 10591
rect 18371 10557 18383 10591
rect 46014 10588 46020 10600
rect 45975 10560 46020 10588
rect 18325 10551 18383 10557
rect 3510 10480 3516 10532
rect 3568 10520 3574 10532
rect 18340 10520 18368 10551
rect 46014 10548 46020 10560
rect 46072 10548 46078 10600
rect 46293 10591 46351 10597
rect 46293 10557 46305 10591
rect 46339 10557 46351 10591
rect 46293 10551 46351 10557
rect 3568 10492 18368 10520
rect 3568 10480 3574 10492
rect 45922 10480 45928 10532
rect 45980 10520 45986 10532
rect 46308 10520 46336 10551
rect 45980 10492 46336 10520
rect 45980 10480 45986 10492
rect 46290 10412 46296 10464
rect 46348 10452 46354 10464
rect 47765 10455 47823 10461
rect 47765 10452 47777 10455
rect 46348 10424 47777 10452
rect 46348 10412 46354 10424
rect 47765 10421 47777 10424
rect 47811 10421 47823 10455
rect 47765 10415 47823 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 18138 10248 18144 10260
rect 18099 10220 18144 10248
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 17954 10004 17960 10056
rect 18012 10044 18018 10056
rect 18049 10047 18107 10053
rect 18049 10044 18061 10047
rect 18012 10016 18061 10044
rect 18012 10004 18018 10016
rect 18049 10013 18061 10016
rect 18095 10013 18107 10047
rect 18049 10007 18107 10013
rect 46477 9979 46535 9985
rect 46477 9945 46489 9979
rect 46523 9976 46535 9979
rect 47670 9976 47676 9988
rect 46523 9948 47676 9976
rect 46523 9945 46535 9948
rect 46477 9939 46535 9945
rect 47670 9936 47676 9948
rect 47728 9936 47734 9988
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 46106 9664 46112 9716
rect 46164 9704 46170 9716
rect 46845 9707 46903 9713
rect 46845 9704 46857 9707
rect 46164 9676 46857 9704
rect 46164 9664 46170 9676
rect 46845 9673 46857 9676
rect 46891 9673 46903 9707
rect 46845 9667 46903 9673
rect 47670 9636 47676 9648
rect 47631 9608 47676 9636
rect 47670 9596 47676 9608
rect 47728 9596 47734 9648
rect 46842 9528 46848 9580
rect 46900 9568 46906 9580
rect 47029 9571 47087 9577
rect 47029 9568 47041 9571
rect 46900 9540 47041 9568
rect 46900 9528 46906 9540
rect 47029 9537 47041 9540
rect 47075 9537 47087 9571
rect 47029 9531 47087 9537
rect 47486 9528 47492 9580
rect 47544 9568 47550 9580
rect 47581 9571 47639 9577
rect 47581 9568 47593 9571
rect 47544 9540 47593 9568
rect 47544 9528 47550 9540
rect 47581 9537 47593 9540
rect 47627 9537 47639 9571
rect 47581 9531 47639 9537
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 47302 8956 47308 8968
rect 47263 8928 47308 8956
rect 47302 8916 47308 8928
rect 47360 8916 47366 8968
rect 47394 8916 47400 8968
rect 47452 8956 47458 8968
rect 47581 8959 47639 8965
rect 47581 8956 47593 8959
rect 47452 8928 47593 8956
rect 47452 8916 47458 8928
rect 47581 8925 47593 8928
rect 47627 8925 47639 8959
rect 47581 8919 47639 8925
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 47670 8480 47676 8492
rect 47631 8452 47676 8480
rect 47670 8440 47676 8452
rect 47728 8440 47734 8492
rect 24946 8372 24952 8424
rect 25004 8412 25010 8424
rect 47857 8415 47915 8421
rect 47857 8412 47869 8415
rect 25004 8384 47869 8412
rect 25004 8372 25010 8384
rect 47857 8381 47869 8384
rect 47903 8381 47915 8415
rect 47857 8375 47915 8381
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 12434 8276 12440 8288
rect 3476 8248 12440 8276
rect 3476 8236 3482 8248
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 17494 8236 17500 8288
rect 17552 8276 17558 8288
rect 45554 8276 45560 8288
rect 17552 8248 45560 8276
rect 17552 8236 17558 8248
rect 45554 8236 45560 8248
rect 45612 8236 45618 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 47854 8004 47860 8016
rect 46308 7976 47860 8004
rect 46308 7945 46336 7976
rect 47854 7964 47860 7976
rect 47912 7964 47918 8016
rect 46293 7939 46351 7945
rect 46293 7905 46305 7939
rect 46339 7905 46351 7939
rect 46293 7899 46351 7905
rect 46477 7939 46535 7945
rect 46477 7905 46489 7939
rect 46523 7936 46535 7939
rect 47394 7936 47400 7948
rect 46523 7908 47400 7936
rect 46523 7905 46535 7908
rect 46477 7899 46535 7905
rect 47394 7896 47400 7908
rect 47452 7896 47458 7948
rect 47670 7936 47676 7948
rect 47631 7908 47676 7936
rect 47670 7896 47676 7908
rect 47728 7896 47734 7948
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 48130 7392 48136 7404
rect 48091 7364 48136 7392
rect 48130 7352 48136 7364
rect 48188 7352 48194 7404
rect 47026 7148 47032 7200
rect 47084 7188 47090 7200
rect 47949 7191 48007 7197
rect 47949 7188 47961 7191
rect 47084 7160 47961 7188
rect 47084 7148 47090 7160
rect 47949 7157 47961 7160
rect 47995 7157 48007 7191
rect 47949 7151 48007 7157
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 18138 6848 18144 6860
rect 3568 6820 18144 6848
rect 3568 6808 3574 6820
rect 18138 6808 18144 6820
rect 18196 6808 18202 6860
rect 47026 6848 47032 6860
rect 46987 6820 47032 6848
rect 47026 6808 47032 6820
rect 47084 6808 47090 6860
rect 48038 6848 48044 6860
rect 47999 6820 48044 6848
rect 48038 6808 48044 6820
rect 48096 6808 48102 6860
rect 1670 6672 1676 6724
rect 1728 6712 1734 6724
rect 47121 6715 47179 6721
rect 1728 6684 22094 6712
rect 1728 6672 1734 6684
rect 22066 6644 22094 6684
rect 47121 6681 47133 6715
rect 47167 6681 47179 6715
rect 47121 6675 47179 6681
rect 47136 6644 47164 6675
rect 22066 6616 47164 6644
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 46477 6307 46535 6313
rect 46477 6273 46489 6307
rect 46523 6304 46535 6307
rect 46566 6304 46572 6316
rect 46523 6276 46572 6304
rect 46523 6273 46535 6276
rect 46477 6267 46535 6273
rect 46566 6264 46572 6276
rect 46624 6264 46630 6316
rect 48130 6304 48136 6316
rect 48091 6276 48136 6304
rect 48130 6264 48136 6276
rect 48188 6264 48194 6316
rect 46198 6236 46204 6248
rect 46159 6208 46204 6236
rect 46198 6196 46204 6208
rect 46256 6196 46262 6248
rect 47946 6100 47952 6112
rect 47907 6072 47952 6100
rect 47946 6060 47952 6072
rect 48004 6060 48010 6112
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 44358 5720 44364 5772
rect 44416 5760 44422 5772
rect 47670 5760 47676 5772
rect 44416 5732 47676 5760
rect 44416 5720 44422 5732
rect 47670 5720 47676 5732
rect 47728 5720 47734 5772
rect 27706 5652 27712 5704
rect 27764 5692 27770 5704
rect 46293 5695 46351 5701
rect 46293 5692 46305 5695
rect 27764 5664 46305 5692
rect 27764 5652 27770 5664
rect 46293 5661 46305 5664
rect 46339 5661 46351 5695
rect 46293 5655 46351 5661
rect 46474 5624 46480 5636
rect 46435 5596 46480 5624
rect 46474 5584 46480 5596
rect 46532 5584 46538 5636
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 46014 5284 46020 5296
rect 45975 5256 46020 5284
rect 46014 5244 46020 5256
rect 46072 5244 46078 5296
rect 46109 5287 46167 5293
rect 46109 5253 46121 5287
rect 46155 5284 46167 5287
rect 47946 5284 47952 5296
rect 46155 5256 47952 5284
rect 46155 5253 46167 5256
rect 46109 5247 46167 5253
rect 47946 5244 47952 5256
rect 48004 5244 48010 5296
rect 47581 5219 47639 5225
rect 47581 5185 47593 5219
rect 47627 5216 47639 5219
rect 47762 5216 47768 5228
rect 47627 5188 47768 5216
rect 47627 5185 47639 5188
rect 47581 5179 47639 5185
rect 47762 5176 47768 5188
rect 47820 5176 47826 5228
rect 46845 5151 46903 5157
rect 46845 5117 46857 5151
rect 46891 5148 46903 5151
rect 48038 5148 48044 5160
rect 46891 5120 48044 5148
rect 46891 5117 46903 5120
rect 46845 5111 46903 5117
rect 48038 5108 48044 5120
rect 48096 5108 48102 5160
rect 47670 5012 47676 5024
rect 47631 4984 47676 5012
rect 47670 4972 47676 4984
rect 47728 4972 47734 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 43530 4632 43536 4684
rect 43588 4672 43594 4684
rect 46014 4672 46020 4684
rect 43588 4644 46020 4672
rect 43588 4632 43594 4644
rect 46014 4632 46020 4644
rect 46072 4672 46078 4684
rect 46109 4675 46167 4681
rect 46109 4672 46121 4675
rect 46072 4644 46121 4672
rect 46072 4632 46078 4644
rect 46109 4641 46121 4644
rect 46155 4641 46167 4675
rect 46566 4672 46572 4684
rect 46527 4644 46572 4672
rect 46109 4635 46167 4641
rect 46566 4632 46572 4644
rect 46624 4632 46630 4684
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 7708 4576 7849 4604
rect 7708 4564 7714 4576
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 7837 4567 7895 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 20254 4604 20260 4616
rect 19751 4576 20260 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 20349 4607 20407 4613
rect 20349 4573 20361 4607
rect 20395 4604 20407 4607
rect 20806 4604 20812 4616
rect 20395 4576 20812 4604
rect 20395 4573 20407 4576
rect 20349 4567 20407 4573
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 20990 4604 20996 4616
rect 20951 4576 20996 4604
rect 20990 4564 20996 4576
rect 21048 4564 21054 4616
rect 21637 4607 21695 4613
rect 21637 4573 21649 4607
rect 21683 4573 21695 4607
rect 21637 4567 21695 4573
rect 21729 4607 21787 4613
rect 21729 4573 21741 4607
rect 21775 4604 21787 4607
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 21775 4576 22293 4604
rect 21775 4573 21787 4576
rect 21729 4567 21787 4573
rect 22281 4573 22293 4576
rect 22327 4573 22339 4607
rect 22281 4567 22339 4573
rect 22925 4607 22983 4613
rect 22925 4573 22937 4607
rect 22971 4604 22983 4607
rect 23566 4604 23572 4616
rect 22971 4576 23572 4604
rect 22971 4573 22983 4576
rect 22925 4567 22983 4573
rect 19797 4539 19855 4545
rect 19797 4505 19809 4539
rect 19843 4536 19855 4539
rect 20898 4536 20904 4548
rect 19843 4508 20904 4536
rect 19843 4505 19855 4508
rect 19797 4499 19855 4505
rect 20898 4496 20904 4508
rect 20956 4496 20962 4548
rect 21652 4536 21680 4567
rect 23566 4564 23572 4576
rect 23624 4564 23630 4616
rect 42886 4604 42892 4616
rect 42847 4576 42892 4604
rect 42886 4564 42892 4576
rect 42944 4564 42950 4616
rect 45646 4604 45652 4616
rect 45607 4576 45652 4604
rect 45646 4564 45652 4576
rect 45704 4564 45710 4616
rect 22738 4536 22744 4548
rect 21652 4508 22744 4536
rect 22738 4496 22744 4508
rect 22796 4496 22802 4548
rect 46290 4536 46296 4548
rect 46251 4508 46296 4536
rect 46290 4496 46296 4508
rect 46348 4496 46354 4548
rect 18601 4471 18659 4477
rect 18601 4437 18613 4471
rect 18647 4468 18659 4471
rect 19426 4468 19432 4480
rect 18647 4440 19432 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 20441 4471 20499 4477
rect 20441 4437 20453 4471
rect 20487 4468 20499 4471
rect 20714 4468 20720 4480
rect 20487 4440 20720 4468
rect 20487 4437 20499 4440
rect 20441 4431 20499 4437
rect 20714 4428 20720 4440
rect 20772 4428 20778 4480
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21358 4468 21364 4480
rect 21131 4440 21364 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21358 4428 21364 4440
rect 21416 4428 21422 4480
rect 22373 4471 22431 4477
rect 22373 4437 22385 4471
rect 22419 4468 22431 4471
rect 22830 4468 22836 4480
rect 22419 4440 22836 4468
rect 22419 4437 22431 4440
rect 22373 4431 22431 4437
rect 22830 4428 22836 4440
rect 22888 4428 22894 4480
rect 23014 4468 23020 4480
rect 22975 4440 23020 4468
rect 23014 4428 23020 4440
rect 23072 4428 23078 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 20254 4224 20260 4276
rect 20312 4264 20318 4276
rect 20441 4267 20499 4273
rect 20441 4264 20453 4267
rect 20312 4236 20453 4264
rect 20312 4224 20318 4236
rect 20441 4233 20453 4236
rect 20487 4233 20499 4267
rect 20441 4227 20499 4233
rect 45738 4196 45744 4208
rect 20824 4168 21128 4196
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 6638 4128 6644 4140
rect 6599 4100 6644 4128
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 8202 4128 8208 4140
rect 8163 4100 8208 4128
rect 7377 4091 7435 4097
rect 7392 4060 7420 4091
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 18141 4131 18199 4137
rect 18141 4097 18153 4131
rect 18187 4128 18199 4131
rect 18966 4128 18972 4140
rect 18187 4100 18972 4128
rect 18187 4097 18199 4100
rect 18141 4091 18199 4097
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4128 19119 4131
rect 19518 4128 19524 4140
rect 19107 4100 19524 4128
rect 19107 4097 19119 4100
rect 19061 4091 19119 4097
rect 19518 4088 19524 4100
rect 19576 4088 19582 4140
rect 19702 4128 19708 4140
rect 19663 4100 19708 4128
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 19797 4131 19855 4137
rect 19797 4097 19809 4131
rect 19843 4128 19855 4131
rect 20349 4131 20407 4137
rect 20349 4128 20361 4131
rect 19843 4100 20361 4128
rect 19843 4097 19855 4100
rect 19797 4091 19855 4097
rect 20349 4097 20361 4100
rect 20395 4097 20407 4131
rect 20824 4128 20852 4168
rect 20349 4091 20407 4097
rect 20456 4100 20852 4128
rect 14090 4060 14096 4072
rect 7392 4032 14096 4060
rect 14090 4020 14096 4032
rect 14148 4020 14154 4072
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 20456 4060 20484 4100
rect 20898 4088 20904 4140
rect 20956 4128 20962 4140
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 20956 4100 21005 4128
rect 20956 4088 20962 4100
rect 20993 4097 21005 4100
rect 21039 4097 21051 4131
rect 21100 4128 21128 4168
rect 23308 4168 24440 4196
rect 22189 4131 22247 4137
rect 21100 4100 21220 4128
rect 20993 4091 21051 4097
rect 18472 4032 20484 4060
rect 18472 4020 18478 4032
rect 20806 4020 20812 4072
rect 20864 4060 20870 4072
rect 21085 4063 21143 4069
rect 21085 4060 21097 4063
rect 20864 4032 21097 4060
rect 20864 4020 20870 4032
rect 21085 4029 21097 4032
rect 21131 4029 21143 4063
rect 21192 4060 21220 4100
rect 22189 4097 22201 4131
rect 22235 4128 22247 4131
rect 22370 4128 22376 4140
rect 22235 4100 22376 4128
rect 22235 4097 22247 4100
rect 22189 4091 22247 4097
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 22830 4128 22836 4140
rect 22791 4100 22836 4128
rect 22830 4088 22836 4100
rect 22888 4088 22894 4140
rect 23308 4128 23336 4168
rect 23474 4128 23480 4140
rect 22940 4100 23336 4128
rect 23435 4100 23480 4128
rect 22462 4060 22468 4072
rect 21192 4032 22468 4060
rect 21085 4023 21143 4029
rect 22462 4020 22468 4032
rect 22520 4020 22526 4072
rect 22554 4020 22560 4072
rect 22612 4060 22618 4072
rect 22940 4060 22968 4100
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 23566 4088 23572 4140
rect 23624 4128 23630 4140
rect 24305 4131 24363 4137
rect 23624 4100 23669 4128
rect 23624 4088 23630 4100
rect 24305 4097 24317 4131
rect 24351 4097 24363 4131
rect 24412 4128 24440 4168
rect 38626 4168 45744 4196
rect 26234 4128 26240 4140
rect 24412 4100 26240 4128
rect 24305 4091 24363 4097
rect 22612 4032 22968 4060
rect 22612 4020 22618 4032
rect 23198 4020 23204 4072
rect 23256 4060 23262 4072
rect 24320 4060 24348 4091
rect 26234 4088 26240 4100
rect 26292 4088 26298 4140
rect 23256 4032 24348 4060
rect 23256 4020 23262 4032
rect 24394 4020 24400 4072
rect 24452 4060 24458 4072
rect 28534 4060 28540 4072
rect 24452 4032 28540 4060
rect 24452 4020 24458 4032
rect 28534 4020 28540 4032
rect 28592 4020 28598 4072
rect 29454 4060 29460 4072
rect 29415 4032 29460 4060
rect 29454 4020 29460 4032
rect 29512 4020 29518 4072
rect 29641 4063 29699 4069
rect 29641 4029 29653 4063
rect 29687 4060 29699 4063
rect 30006 4060 30012 4072
rect 29687 4032 30012 4060
rect 29687 4029 29699 4032
rect 29641 4023 29699 4029
rect 30006 4020 30012 4032
rect 30064 4020 30070 4072
rect 31297 4063 31355 4069
rect 31297 4029 31309 4063
rect 31343 4060 31355 4063
rect 38626 4060 38654 4168
rect 45738 4156 45744 4168
rect 45796 4196 45802 4208
rect 46566 4196 46572 4208
rect 45796 4168 46572 4196
rect 45796 4156 45802 4168
rect 46566 4156 46572 4168
rect 46624 4156 46630 4208
rect 47762 4196 47768 4208
rect 47723 4168 47768 4196
rect 47762 4156 47768 4168
rect 47820 4156 47826 4208
rect 39206 4088 39212 4140
rect 39264 4128 39270 4140
rect 39945 4131 40003 4137
rect 39945 4128 39957 4131
rect 39264 4100 39957 4128
rect 39264 4088 39270 4100
rect 39945 4097 39957 4100
rect 39991 4097 40003 4131
rect 39945 4091 40003 4097
rect 42797 4131 42855 4137
rect 42797 4097 42809 4131
rect 42843 4128 42855 4131
rect 43438 4128 43444 4140
rect 42843 4100 43444 4128
rect 42843 4097 42855 4100
rect 42797 4091 42855 4097
rect 43438 4088 43444 4100
rect 43496 4088 43502 4140
rect 46474 4128 46480 4140
rect 46435 4100 46480 4128
rect 46474 4088 46480 4100
rect 46532 4088 46538 4140
rect 31343 4032 38654 4060
rect 31343 4029 31355 4032
rect 31297 4023 31355 4029
rect 41322 4020 41328 4072
rect 41380 4060 41386 4072
rect 43530 4060 43536 4072
rect 41380 4032 43536 4060
rect 41380 4020 41386 4032
rect 43530 4020 43536 4032
rect 43588 4020 43594 4072
rect 43714 4060 43720 4072
rect 43675 4032 43720 4060
rect 43714 4020 43720 4032
rect 43772 4020 43778 4072
rect 43806 4020 43812 4072
rect 43864 4060 43870 4072
rect 43993 4063 44051 4069
rect 43993 4060 44005 4063
rect 43864 4032 44005 4060
rect 43864 4020 43870 4032
rect 43993 4029 44005 4032
rect 44039 4029 44051 4063
rect 43993 4023 44051 4029
rect 46201 4063 46259 4069
rect 46201 4029 46213 4063
rect 46247 4060 46259 4063
rect 48314 4060 48320 4072
rect 46247 4032 48320 4060
rect 46247 4029 46259 4032
rect 46201 4023 46259 4029
rect 48314 4020 48320 4032
rect 48372 4020 48378 4072
rect 19978 3952 19984 4004
rect 20036 3992 20042 4004
rect 22925 3995 22983 4001
rect 22925 3992 22937 3995
rect 20036 3964 22937 3992
rect 20036 3952 20042 3964
rect 22925 3961 22937 3964
rect 22971 3961 22983 3995
rect 22925 3955 22983 3961
rect 23106 3952 23112 4004
rect 23164 3992 23170 4004
rect 23164 3964 24808 3992
rect 23164 3952 23170 3964
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1636 3896 2145 3924
rect 1636 3884 1642 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2133 3887 2191 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2832 3896 2881 3924
rect 2832 3884 2838 3896
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 6730 3924 6736 3936
rect 6691 3896 6736 3924
rect 2869 3887 2927 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7466 3924 7472 3936
rect 7427 3896 7472 3924
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 7834 3884 7840 3936
rect 7892 3924 7898 3936
rect 8297 3927 8355 3933
rect 8297 3924 8309 3927
rect 7892 3896 8309 3924
rect 7892 3884 7898 3896
rect 8297 3893 8309 3896
rect 8343 3893 8355 3927
rect 8297 3887 8355 3893
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 9272 3896 9413 3924
rect 9272 3884 9278 3896
rect 9401 3893 9413 3896
rect 9447 3893 9459 3927
rect 9401 3887 9459 3893
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11572 3896 11713 3924
rect 11572 3884 11578 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 18233 3927 18291 3933
rect 18233 3893 18245 3927
rect 18279 3924 18291 3927
rect 19058 3924 19064 3936
rect 18279 3896 19064 3924
rect 18279 3893 18291 3896
rect 18233 3887 18291 3893
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 19153 3927 19211 3933
rect 19153 3893 19165 3927
rect 19199 3924 19211 3927
rect 20254 3924 20260 3936
rect 19199 3896 20260 3924
rect 19199 3893 19211 3896
rect 19153 3887 19211 3893
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 21726 3924 21732 3936
rect 20588 3896 21732 3924
rect 20588 3884 20594 3896
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 22281 3927 22339 3933
rect 22281 3893 22293 3927
rect 22327 3924 22339 3927
rect 22370 3924 22376 3936
rect 22327 3896 22376 3924
rect 22327 3893 22339 3896
rect 22281 3887 22339 3893
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 24121 3927 24179 3933
rect 24121 3893 24133 3927
rect 24167 3924 24179 3927
rect 24670 3924 24676 3936
rect 24167 3896 24676 3924
rect 24167 3893 24179 3896
rect 24121 3887 24179 3893
rect 24670 3884 24676 3896
rect 24728 3884 24734 3936
rect 24780 3924 24808 3964
rect 26878 3952 26884 4004
rect 26936 3992 26942 4004
rect 33962 3992 33968 4004
rect 26936 3964 33968 3992
rect 26936 3952 26942 3964
rect 33962 3952 33968 3964
rect 34020 3952 34026 4004
rect 47949 3995 48007 4001
rect 47949 3992 47961 3995
rect 34072 3964 47961 3992
rect 34072 3924 34100 3964
rect 47949 3961 47961 3964
rect 47995 3961 48007 3995
rect 47949 3955 48007 3961
rect 40034 3924 40040 3936
rect 24780 3896 34100 3924
rect 39995 3896 40040 3924
rect 40034 3884 40040 3896
rect 40092 3884 40098 3936
rect 42794 3884 42800 3936
rect 42852 3924 42858 3936
rect 42889 3927 42947 3933
rect 42889 3924 42901 3927
rect 42852 3896 42901 3924
rect 42852 3884 42858 3896
rect 42889 3893 42901 3896
rect 42935 3893 42947 3927
rect 42889 3887 42947 3893
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 6914 3680 6920 3732
rect 6972 3720 6978 3732
rect 15286 3720 15292 3732
rect 6972 3692 15292 3720
rect 6972 3680 6978 3692
rect 15286 3680 15292 3692
rect 15344 3680 15350 3732
rect 19518 3720 19524 3732
rect 19479 3692 19524 3720
rect 19518 3680 19524 3692
rect 19576 3680 19582 3732
rect 19702 3680 19708 3732
rect 19760 3720 19766 3732
rect 20165 3723 20223 3729
rect 20165 3720 20177 3723
rect 19760 3692 20177 3720
rect 19760 3680 19766 3692
rect 20165 3689 20177 3692
rect 20211 3689 20223 3723
rect 20165 3683 20223 3689
rect 20809 3723 20867 3729
rect 20809 3689 20821 3723
rect 20855 3720 20867 3723
rect 20990 3720 20996 3732
rect 20855 3692 20996 3720
rect 20855 3689 20867 3692
rect 20809 3683 20867 3689
rect 20990 3680 20996 3692
rect 21048 3680 21054 3732
rect 22554 3720 22560 3732
rect 22066 3692 22560 3720
rect 9030 3612 9036 3664
rect 9088 3652 9094 3664
rect 9088 3624 9720 3652
rect 9088 3612 9094 3624
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 1820 3556 3985 3584
rect 1820 3544 1826 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 6730 3584 6736 3596
rect 6691 3556 6736 3584
rect 3973 3547 4031 3553
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 7098 3584 7104 3596
rect 7059 3556 7104 3584
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 9214 3584 9220 3596
rect 9175 3556 9220 3584
rect 9214 3544 9220 3556
rect 9272 3544 9278 3596
rect 9692 3593 9720 3624
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 19886 3652 19892 3664
rect 10008 3624 19892 3652
rect 10008 3612 10014 3624
rect 19886 3612 19892 3624
rect 19944 3612 19950 3664
rect 22066 3652 22094 3692
rect 22554 3680 22560 3692
rect 22612 3680 22618 3732
rect 22738 3680 22744 3732
rect 22796 3720 22802 3732
rect 22925 3723 22983 3729
rect 22925 3720 22937 3723
rect 22796 3692 22937 3720
rect 22796 3680 22802 3692
rect 22925 3689 22937 3692
rect 22971 3689 22983 3723
rect 22925 3683 22983 3689
rect 23382 3680 23388 3732
rect 23440 3720 23446 3732
rect 23440 3692 28488 3720
rect 23440 3680 23446 3692
rect 19996 3624 22094 3652
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3553 9735 3587
rect 19242 3584 19248 3596
rect 9677 3547 9735 3553
rect 12084 3556 19248 3584
rect 2682 3516 2688 3528
rect 2643 3488 2688 3516
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 12084 3525 12112 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3516 6147 3519
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6135 3488 6561 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 12069 3519 12127 3525
rect 12069 3485 12081 3519
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13814 3516 13820 3528
rect 13587 3488 13820 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 14090 3516 14096 3528
rect 14051 3488 14096 3516
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3516 17739 3519
rect 17954 3516 17960 3528
rect 17727 3488 17960 3516
rect 17727 3485 17739 3488
rect 17681 3479 17739 3485
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 18598 3516 18604 3528
rect 18371 3488 18604 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 19426 3516 19432 3528
rect 19387 3488 19432 3516
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 19996 3516 20024 3624
rect 22186 3612 22192 3664
rect 22244 3652 22250 3664
rect 28460 3652 28488 3692
rect 28534 3680 28540 3732
rect 28592 3720 28598 3732
rect 28592 3692 33916 3720
rect 28592 3680 28598 3692
rect 33042 3652 33048 3664
rect 22244 3624 28396 3652
rect 28460 3624 33048 3652
rect 22244 3612 22250 3624
rect 20162 3544 20168 3596
rect 20220 3584 20226 3596
rect 21450 3584 21456 3596
rect 20220 3556 21456 3584
rect 20220 3544 20226 3556
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 21542 3544 21548 3596
rect 21600 3584 21606 3596
rect 21600 3556 24716 3584
rect 21600 3544 21606 3556
rect 19536 3488 20024 3516
rect 20073 3519 20131 3525
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 1857 3451 1915 3457
rect 1857 3448 1869 3451
rect 1360 3420 1869 3448
rect 1360 3408 1366 3420
rect 1857 3417 1869 3420
rect 1903 3417 1915 3451
rect 1857 3411 1915 3417
rect 2225 3451 2283 3457
rect 2225 3417 2237 3451
rect 2271 3448 2283 3451
rect 9401 3451 9459 3457
rect 2271 3420 6914 3448
rect 2271 3417 2283 3420
rect 2225 3411 2283 3417
rect 1946 3340 1952 3392
rect 2004 3380 2010 3392
rect 2777 3383 2835 3389
rect 2777 3380 2789 3383
rect 2004 3352 2789 3380
rect 2004 3340 2010 3352
rect 2777 3349 2789 3352
rect 2823 3349 2835 3383
rect 6886 3380 6914 3420
rect 9401 3417 9413 3451
rect 9447 3448 9459 3451
rect 10042 3448 10048 3460
rect 9447 3420 10048 3448
rect 9447 3417 9459 3420
rect 9401 3411 9459 3417
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 15470 3448 15476 3460
rect 11348 3420 14320 3448
rect 15431 3420 15476 3448
rect 11348 3380 11376 3420
rect 6886 3352 11376 3380
rect 2777 3343 2835 3349
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 12161 3383 12219 3389
rect 12161 3380 12173 3383
rect 11756 3352 12173 3380
rect 11756 3340 11762 3352
rect 12161 3349 12173 3352
rect 12207 3349 12219 3383
rect 12161 3343 12219 3349
rect 13998 3340 14004 3392
rect 14056 3380 14062 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 14056 3352 14197 3380
rect 14056 3340 14062 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14292 3380 14320 3420
rect 15470 3408 15476 3420
rect 15528 3408 15534 3460
rect 17126 3448 17132 3460
rect 17087 3420 17132 3448
rect 17126 3408 17132 3420
rect 17184 3408 17190 3460
rect 19536 3448 19564 3488
rect 20073 3485 20085 3519
rect 20119 3516 20131 3519
rect 20254 3516 20260 3528
rect 20119 3488 20260 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 20714 3516 20720 3528
rect 20675 3488 20720 3516
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 21358 3516 21364 3528
rect 21319 3488 21364 3516
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 22094 3476 22100 3528
rect 22152 3516 22158 3528
rect 22373 3519 22431 3525
rect 22373 3516 22385 3519
rect 22152 3488 22385 3516
rect 22152 3476 22158 3488
rect 22373 3485 22385 3488
rect 22419 3485 22431 3519
rect 22830 3516 22836 3528
rect 22791 3488 22836 3516
rect 22373 3479 22431 3485
rect 22830 3476 22836 3488
rect 22888 3476 22894 3528
rect 24688 3525 24716 3556
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3485 23535 3519
rect 23477 3479 23535 3485
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3485 24731 3519
rect 24673 3479 24731 3485
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3485 25559 3519
rect 25501 3479 25559 3485
rect 17696 3420 19564 3448
rect 17696 3380 17724 3420
rect 20162 3408 20168 3460
rect 20220 3448 20226 3460
rect 23492 3448 23520 3479
rect 20220 3420 23520 3448
rect 20220 3408 20226 3420
rect 24578 3408 24584 3460
rect 24636 3448 24642 3460
rect 25516 3448 25544 3479
rect 24636 3420 25544 3448
rect 28368 3448 28396 3624
rect 33042 3612 33048 3624
rect 33100 3612 33106 3664
rect 33888 3652 33916 3692
rect 33962 3680 33968 3732
rect 34020 3720 34026 3732
rect 34020 3692 43392 3720
rect 34020 3680 34026 3692
rect 33888 3624 35388 3652
rect 29546 3584 29552 3596
rect 29507 3556 29552 3584
rect 29546 3544 29552 3556
rect 29604 3544 29610 3596
rect 29733 3587 29791 3593
rect 29733 3553 29745 3587
rect 29779 3584 29791 3587
rect 29779 3556 31708 3584
rect 29779 3553 29791 3556
rect 29733 3547 29791 3553
rect 31680 3516 31708 3556
rect 32876 3556 34192 3584
rect 32876 3516 32904 3556
rect 33042 3516 33048 3528
rect 31680 3488 32904 3516
rect 33003 3488 33048 3516
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33873 3519 33931 3525
rect 33873 3485 33885 3519
rect 33919 3485 33931 3519
rect 33873 3479 33931 3485
rect 31389 3451 31447 3457
rect 31389 3448 31401 3451
rect 28368 3420 31401 3448
rect 24636 3408 24642 3420
rect 31389 3417 31401 3420
rect 31435 3448 31447 3451
rect 31435 3420 31754 3448
rect 31435 3417 31447 3420
rect 31389 3411 31447 3417
rect 14292 3352 17724 3380
rect 17773 3383 17831 3389
rect 14185 3343 14243 3349
rect 17773 3349 17785 3383
rect 17819 3380 17831 3383
rect 18322 3380 18328 3392
rect 17819 3352 18328 3380
rect 17819 3349 17831 3352
rect 17773 3343 17831 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 18417 3383 18475 3389
rect 18417 3349 18429 3383
rect 18463 3380 18475 3383
rect 19150 3380 19156 3392
rect 18463 3352 19156 3380
rect 18463 3349 18475 3352
rect 18417 3343 18475 3349
rect 19150 3340 19156 3352
rect 19208 3340 19214 3392
rect 19242 3340 19248 3392
rect 19300 3380 19306 3392
rect 20530 3380 20536 3392
rect 19300 3352 20536 3380
rect 19300 3340 19306 3352
rect 20530 3340 20536 3352
rect 20588 3340 20594 3392
rect 20622 3340 20628 3392
rect 20680 3380 20686 3392
rect 21453 3383 21511 3389
rect 21453 3380 21465 3383
rect 20680 3352 21465 3380
rect 20680 3340 20686 3352
rect 21453 3349 21465 3352
rect 21499 3349 21511 3383
rect 21453 3343 21511 3349
rect 21726 3340 21732 3392
rect 21784 3380 21790 3392
rect 23382 3380 23388 3392
rect 21784 3352 23388 3380
rect 21784 3340 21790 3352
rect 23382 3340 23388 3352
rect 23440 3340 23446 3392
rect 23569 3383 23627 3389
rect 23569 3349 23581 3383
rect 23615 3380 23627 3383
rect 23658 3380 23664 3392
rect 23615 3352 23664 3380
rect 23615 3349 23627 3352
rect 23569 3343 23627 3349
rect 23658 3340 23664 3352
rect 23716 3340 23722 3392
rect 24762 3380 24768 3392
rect 24723 3352 24768 3380
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 24854 3340 24860 3392
rect 24912 3380 24918 3392
rect 31294 3380 31300 3392
rect 24912 3352 31300 3380
rect 24912 3340 24918 3352
rect 31294 3340 31300 3352
rect 31352 3340 31358 3392
rect 31726 3380 31754 3420
rect 32950 3408 32956 3460
rect 33008 3448 33014 3460
rect 33888 3448 33916 3479
rect 33008 3420 33916 3448
rect 33008 3408 33014 3420
rect 32858 3380 32864 3392
rect 31726 3352 32864 3380
rect 32858 3340 32864 3352
rect 32916 3340 32922 3392
rect 33134 3380 33140 3392
rect 33095 3352 33140 3380
rect 33134 3340 33140 3352
rect 33192 3340 33198 3392
rect 34164 3380 34192 3556
rect 35360 3516 35388 3624
rect 35434 3612 35440 3664
rect 35492 3652 35498 3664
rect 42518 3652 42524 3664
rect 35492 3624 42524 3652
rect 35492 3612 35498 3624
rect 42518 3612 42524 3624
rect 42576 3612 42582 3664
rect 42886 3652 42892 3664
rect 42628 3624 42892 3652
rect 42628 3593 42656 3624
rect 42886 3612 42892 3624
rect 42944 3612 42950 3664
rect 43364 3652 43392 3692
rect 43438 3680 43444 3732
rect 43496 3720 43502 3732
rect 46658 3720 46664 3732
rect 43496 3692 46664 3720
rect 43496 3680 43502 3692
rect 46658 3680 46664 3692
rect 46716 3680 46722 3732
rect 47210 3652 47216 3664
rect 43364 3624 47216 3652
rect 47210 3612 47216 3624
rect 47268 3612 47274 3664
rect 37737 3587 37795 3593
rect 37737 3553 37749 3587
rect 37783 3584 37795 3587
rect 42613 3587 42671 3593
rect 37783 3556 42564 3584
rect 37783 3553 37795 3556
rect 37737 3547 37795 3553
rect 35894 3516 35900 3528
rect 35360 3488 35900 3516
rect 35894 3476 35900 3488
rect 35952 3476 35958 3528
rect 39114 3516 39120 3528
rect 39075 3488 39120 3516
rect 39114 3476 39120 3488
rect 39172 3476 39178 3528
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 40000 3488 40049 3516
rect 40000 3476 40006 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 40313 3519 40371 3525
rect 40313 3485 40325 3519
rect 40359 3485 40371 3519
rect 41322 3516 41328 3528
rect 41283 3488 41328 3516
rect 40313 3479 40371 3485
rect 36081 3451 36139 3457
rect 36081 3417 36093 3451
rect 36127 3448 36139 3451
rect 36170 3448 36176 3460
rect 36127 3420 36176 3448
rect 36127 3417 36139 3420
rect 36081 3411 36139 3417
rect 36170 3408 36176 3420
rect 36228 3408 36234 3460
rect 36280 3420 39344 3448
rect 36280 3380 36308 3420
rect 34164 3352 36308 3380
rect 37918 3340 37924 3392
rect 37976 3380 37982 3392
rect 39209 3383 39267 3389
rect 39209 3380 39221 3383
rect 37976 3352 39221 3380
rect 37976 3340 37982 3352
rect 39209 3349 39221 3352
rect 39255 3349 39267 3383
rect 39316 3380 39344 3420
rect 39850 3408 39856 3460
rect 39908 3448 39914 3460
rect 40328 3448 40356 3479
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41506 3516 41512 3528
rect 41467 3488 41512 3516
rect 41506 3476 41512 3488
rect 41564 3476 41570 3528
rect 39908 3420 40356 3448
rect 42536 3448 42564 3556
rect 42613 3553 42625 3587
rect 42659 3553 42671 3587
rect 42794 3584 42800 3596
rect 42755 3556 42800 3584
rect 42613 3547 42671 3553
rect 42794 3544 42800 3556
rect 42852 3544 42858 3596
rect 43162 3584 43168 3596
rect 43123 3556 43168 3584
rect 43162 3544 43168 3556
rect 43220 3544 43226 3596
rect 45189 3587 45247 3593
rect 45189 3553 45201 3587
rect 45235 3584 45247 3587
rect 46293 3587 46351 3593
rect 46293 3584 46305 3587
rect 45235 3556 46305 3584
rect 45235 3553 45247 3556
rect 45189 3547 45247 3553
rect 46293 3553 46305 3556
rect 46339 3553 46351 3587
rect 46293 3547 46351 3553
rect 46477 3587 46535 3593
rect 46477 3553 46489 3587
rect 46523 3584 46535 3587
rect 47670 3584 47676 3596
rect 46523 3556 47676 3584
rect 46523 3553 46535 3556
rect 46477 3547 46535 3553
rect 47670 3544 47676 3556
rect 47728 3544 47734 3596
rect 45649 3519 45707 3525
rect 45649 3485 45661 3519
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 44266 3448 44272 3460
rect 42536 3420 44272 3448
rect 39908 3408 39914 3420
rect 44266 3408 44272 3420
rect 44324 3408 44330 3460
rect 45664 3448 45692 3479
rect 47486 3448 47492 3460
rect 45664 3420 47492 3448
rect 47486 3408 47492 3420
rect 47544 3408 47550 3460
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 40126 3380 40132 3392
rect 39316 3352 40132 3380
rect 39209 3343 39267 3349
rect 40126 3340 40132 3352
rect 40184 3340 40190 3392
rect 41969 3383 42027 3389
rect 41969 3349 41981 3383
rect 42015 3380 42027 3383
rect 42426 3380 42432 3392
rect 42015 3352 42432 3380
rect 42015 3349 42027 3352
rect 41969 3343 42027 3349
rect 42426 3340 42432 3352
rect 42484 3340 42490 3392
rect 45370 3340 45376 3392
rect 45428 3380 45434 3392
rect 45741 3383 45799 3389
rect 45741 3380 45753 3383
rect 45428 3352 45753 3380
rect 45428 3340 45434 3352
rect 45741 3349 45753 3352
rect 45787 3349 45799 3383
rect 45741 3343 45799 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 17954 3176 17960 3188
rect 3936 3148 16574 3176
rect 17915 3148 17960 3176
rect 3936 3136 3942 3148
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 7834 3108 7840 3120
rect 7795 3080 7840 3108
rect 7834 3068 7840 3080
rect 7892 3068 7898 3120
rect 10042 3108 10048 3120
rect 10003 3080 10048 3108
rect 10042 3068 10048 3080
rect 10100 3068 10106 3120
rect 11698 3108 11704 3120
rect 11659 3080 11704 3108
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 13998 3108 14004 3120
rect 13959 3080 14004 3108
rect 13998 3068 14004 3080
rect 14056 3068 14062 3120
rect 16546 3108 16574 3148
rect 17954 3136 17960 3148
rect 18012 3136 18018 3188
rect 18598 3176 18604 3188
rect 18559 3148 18604 3176
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 18966 3136 18972 3188
rect 19024 3176 19030 3188
rect 19245 3179 19303 3185
rect 19245 3176 19257 3179
rect 19024 3148 19257 3176
rect 19024 3136 19030 3148
rect 19245 3145 19257 3148
rect 19291 3145 19303 3179
rect 19245 3139 19303 3145
rect 20073 3179 20131 3185
rect 20073 3145 20085 3179
rect 20119 3176 20131 3179
rect 20162 3176 20168 3188
rect 20119 3148 20168 3176
rect 20119 3145 20131 3148
rect 20073 3139 20131 3145
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 20714 3176 20720 3188
rect 20675 3148 20720 3176
rect 20714 3136 20720 3148
rect 20772 3136 20778 3188
rect 36170 3176 36176 3188
rect 21744 3148 33272 3176
rect 36131 3148 36176 3176
rect 21744 3108 21772 3148
rect 16546 3080 21772 3108
rect 22281 3111 22339 3117
rect 22281 3077 22293 3111
rect 22327 3108 22339 3111
rect 22370 3108 22376 3120
rect 22327 3080 22376 3108
rect 22327 3077 22339 3080
rect 22281 3071 22339 3077
rect 22370 3068 22376 3080
rect 22428 3068 22434 3120
rect 22462 3068 22468 3120
rect 22520 3108 22526 3120
rect 24762 3108 24768 3120
rect 22520 3080 23520 3108
rect 24723 3080 24768 3108
rect 22520 3068 22526 3080
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 7650 3040 7656 3052
rect 7611 3012 7656 3040
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 9950 3040 9956 3052
rect 9911 3012 9956 3040
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 13814 3040 13820 3052
rect 13775 3012 13820 3040
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 17310 3040 17316 3052
rect 17083 3012 17316 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 17865 3043 17923 3049
rect 17865 3040 17877 3043
rect 17420 3012 17877 3040
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 716 2944 2237 2972
rect 716 2932 722 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 8113 2975 8171 2981
rect 8113 2972 8125 2975
rect 2225 2935 2283 2941
rect 7760 2944 8125 2972
rect 7760 2916 7788 2944
rect 8113 2941 8125 2944
rect 8159 2941 8171 2975
rect 8113 2935 8171 2941
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11020 2944 11989 2972
rect 11020 2932 11026 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14240 2944 14289 2972
rect 14240 2932 14246 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 15194 2932 15200 2984
rect 15252 2972 15258 2984
rect 17420 2981 17448 3012
rect 17865 3009 17877 3012
rect 17911 3009 17923 3043
rect 17865 3003 17923 3009
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 18380 3012 18521 3040
rect 18380 3000 18386 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 19150 3040 19156 3052
rect 19111 3012 19156 3040
rect 18509 3003 18567 3009
rect 19150 3000 19156 3012
rect 19208 3000 19214 3052
rect 19978 3040 19984 3052
rect 19939 3012 19984 3040
rect 19978 3000 19984 3012
rect 20036 3000 20042 3052
rect 20622 3040 20628 3052
rect 20583 3012 20628 3040
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 16945 2975 17003 2981
rect 16945 2972 16957 2975
rect 15252 2944 16957 2972
rect 15252 2932 15258 2944
rect 16945 2941 16957 2944
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 17678 2932 17684 2984
rect 17736 2972 17742 2984
rect 21542 2972 21548 2984
rect 17736 2944 21548 2972
rect 17736 2932 17742 2944
rect 21542 2932 21548 2944
rect 21600 2932 21606 2984
rect 22094 2932 22100 2984
rect 22152 2981 22158 2984
rect 22152 2972 22160 2981
rect 22925 2975 22983 2981
rect 22152 2944 22197 2972
rect 22152 2935 22160 2944
rect 22925 2941 22937 2975
rect 22971 2941 22983 2975
rect 22925 2935 22983 2941
rect 22152 2932 22158 2935
rect 7742 2864 7748 2916
rect 7800 2864 7806 2916
rect 14090 2864 14096 2916
rect 14148 2904 14154 2916
rect 22462 2904 22468 2916
rect 14148 2876 22468 2904
rect 14148 2864 14154 2876
rect 22462 2864 22468 2876
rect 22520 2864 22526 2916
rect 22554 2864 22560 2916
rect 22612 2904 22618 2916
rect 22940 2904 22968 2935
rect 22612 2876 22968 2904
rect 23492 2904 23520 3080
rect 24762 3068 24768 3080
rect 24820 3068 24826 3120
rect 27617 3111 27675 3117
rect 27617 3077 27629 3111
rect 27663 3108 27675 3111
rect 27982 3108 27988 3120
rect 27663 3080 27988 3108
rect 27663 3077 27675 3080
rect 27617 3071 27675 3077
rect 27982 3068 27988 3080
rect 28040 3068 28046 3120
rect 33134 3108 33140 3120
rect 33095 3080 33140 3108
rect 33134 3068 33140 3080
rect 33192 3068 33198 3120
rect 33244 3108 33272 3148
rect 36170 3136 36176 3148
rect 36228 3136 36234 3188
rect 38562 3136 38568 3188
rect 38620 3176 38626 3188
rect 41230 3176 41236 3188
rect 38620 3148 41236 3176
rect 38620 3136 38626 3148
rect 41230 3136 41236 3148
rect 41288 3136 41294 3188
rect 45278 3176 45284 3188
rect 41386 3148 45284 3176
rect 41386 3108 41414 3148
rect 45278 3136 45284 3148
rect 45336 3136 45342 3188
rect 33244 3080 41414 3108
rect 41506 3068 41512 3120
rect 41564 3108 41570 3120
rect 42613 3111 42671 3117
rect 42613 3108 42625 3111
rect 41564 3080 42625 3108
rect 41564 3068 41570 3080
rect 42613 3077 42625 3080
rect 42659 3077 42671 3111
rect 42613 3071 42671 3077
rect 44269 3111 44327 3117
rect 44269 3077 44281 3111
rect 44315 3108 44327 3111
rect 44358 3108 44364 3120
rect 44315 3080 44364 3108
rect 44315 3077 44327 3080
rect 44269 3071 44327 3077
rect 24578 3040 24584 3052
rect 24539 3012 24584 3040
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 27062 3000 27068 3052
rect 27120 3040 27126 3052
rect 27433 3043 27491 3049
rect 27433 3040 27445 3043
rect 27120 3012 27445 3040
rect 27120 3000 27126 3012
rect 27433 3009 27445 3012
rect 27479 3009 27491 3043
rect 32214 3040 32220 3052
rect 27433 3003 27491 3009
rect 31726 3012 32220 3040
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 31726 2972 31754 3012
rect 32214 3000 32220 3012
rect 32272 3000 32278 3052
rect 32950 3040 32956 3052
rect 32911 3012 32956 3040
rect 32950 3000 32956 3012
rect 33008 3000 33014 3052
rect 36078 3000 36084 3052
rect 36136 3040 36142 3052
rect 36357 3043 36415 3049
rect 36357 3040 36369 3043
rect 36136 3012 36369 3040
rect 36136 3000 36142 3012
rect 36357 3009 36369 3012
rect 36403 3009 36415 3043
rect 37918 3040 37924 3052
rect 37879 3012 37924 3040
rect 36357 3003 36415 3009
rect 37918 3000 37924 3012
rect 37976 3000 37982 3052
rect 38013 3043 38071 3049
rect 38013 3009 38025 3043
rect 38059 3040 38071 3043
rect 39669 3043 39727 3049
rect 39669 3040 39681 3043
rect 38059 3012 39681 3040
rect 38059 3009 38071 3012
rect 38013 3003 38071 3009
rect 39669 3009 39681 3012
rect 39715 3009 39727 3043
rect 42426 3040 42432 3052
rect 42387 3012 42432 3040
rect 39669 3003 39727 3009
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 33502 2972 33508 2984
rect 25240 2944 31754 2972
rect 33463 2944 33508 2972
rect 25240 2904 25268 2944
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 35894 2932 35900 2984
rect 35952 2972 35958 2984
rect 38562 2972 38568 2984
rect 35952 2944 38568 2972
rect 35952 2932 35958 2944
rect 38562 2932 38568 2944
rect 38620 2932 38626 2984
rect 38749 2975 38807 2981
rect 38749 2941 38761 2975
rect 38795 2972 38807 2975
rect 39850 2972 39856 2984
rect 38795 2944 39856 2972
rect 38795 2941 38807 2944
rect 38749 2935 38807 2941
rect 39850 2932 39856 2944
rect 39908 2932 39914 2984
rect 41509 2975 41567 2981
rect 41509 2972 41521 2975
rect 39960 2944 41521 2972
rect 23492 2876 25268 2904
rect 22612 2864 22618 2876
rect 29086 2864 29092 2916
rect 29144 2904 29150 2916
rect 39022 2904 39028 2916
rect 29144 2876 39028 2904
rect 29144 2864 29150 2876
rect 39022 2864 39028 2876
rect 39080 2864 39086 2916
rect 39206 2904 39212 2916
rect 39167 2876 39212 2904
rect 39206 2864 39212 2876
rect 39264 2864 39270 2916
rect 6822 2836 6828 2848
rect 6783 2808 6828 2836
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 19886 2836 19892 2848
rect 17460 2808 19892 2836
rect 17460 2796 17466 2808
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 21174 2836 21180 2848
rect 20036 2808 21180 2836
rect 20036 2796 20042 2808
rect 21174 2796 21180 2808
rect 21232 2796 21238 2848
rect 21266 2796 21272 2848
rect 21324 2836 21330 2848
rect 26878 2836 26884 2848
rect 21324 2808 26884 2836
rect 21324 2796 21330 2808
rect 26878 2796 26884 2808
rect 26936 2796 26942 2848
rect 27614 2796 27620 2848
rect 27672 2836 27678 2848
rect 30926 2836 30932 2848
rect 27672 2808 30932 2836
rect 27672 2796 27678 2808
rect 30926 2796 30932 2808
rect 30984 2796 30990 2848
rect 32858 2796 32864 2848
rect 32916 2836 32922 2848
rect 39960 2836 39988 2944
rect 41509 2941 41521 2944
rect 41555 2972 41567 2975
rect 44284 2972 44312 3071
rect 44358 3068 44364 3080
rect 44416 3068 44422 3120
rect 45370 3108 45376 3120
rect 45331 3080 45376 3108
rect 45370 3068 45376 3080
rect 45428 3068 45434 3120
rect 47762 3040 47768 3052
rect 47723 3012 47768 3040
rect 47762 3000 47768 3012
rect 47820 3000 47826 3052
rect 41555 2944 44312 2972
rect 45189 2975 45247 2981
rect 41555 2941 41567 2944
rect 41509 2935 41567 2941
rect 45189 2941 45201 2975
rect 45235 2972 45247 2975
rect 45646 2972 45652 2984
rect 45235 2944 45652 2972
rect 45235 2941 45247 2944
rect 45189 2935 45247 2941
rect 45646 2932 45652 2944
rect 45704 2932 45710 2984
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 32916 2808 39988 2836
rect 32916 2796 32922 2808
rect 40126 2796 40132 2848
rect 40184 2836 40190 2848
rect 44358 2836 44364 2848
rect 40184 2808 44364 2836
rect 40184 2796 40190 2808
rect 44358 2796 44364 2808
rect 44416 2796 44422 2848
rect 47854 2836 47860 2848
rect 47815 2808 47860 2836
rect 47854 2796 47860 2808
rect 47912 2796 47918 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 3234 2592 3240 2644
rect 3292 2632 3298 2644
rect 10410 2632 10416 2644
rect 3292 2604 10416 2632
rect 3292 2592 3298 2604
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 15470 2592 15476 2644
rect 15528 2632 15534 2644
rect 15565 2635 15623 2641
rect 15565 2632 15577 2635
rect 15528 2604 15577 2632
rect 15528 2592 15534 2604
rect 15565 2601 15577 2604
rect 15611 2601 15623 2635
rect 15565 2595 15623 2601
rect 16942 2592 16948 2644
rect 17000 2632 17006 2644
rect 17221 2635 17279 2641
rect 17221 2632 17233 2635
rect 17000 2604 17233 2632
rect 17000 2592 17006 2604
rect 17221 2601 17233 2604
rect 17267 2601 17279 2635
rect 17221 2595 17279 2601
rect 17865 2635 17923 2641
rect 17865 2601 17877 2635
rect 17911 2632 17923 2635
rect 18506 2632 18512 2644
rect 17911 2604 18512 2632
rect 17911 2601 17923 2604
rect 17865 2595 17923 2601
rect 18506 2592 18512 2604
rect 18564 2592 18570 2644
rect 19886 2592 19892 2644
rect 19944 2632 19950 2644
rect 21266 2632 21272 2644
rect 19944 2604 21272 2632
rect 19944 2592 19950 2604
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 23474 2592 23480 2644
rect 23532 2632 23538 2644
rect 23753 2635 23811 2641
rect 23753 2632 23765 2635
rect 23532 2604 23765 2632
rect 23532 2592 23538 2604
rect 23753 2601 23765 2604
rect 23799 2601 23811 2635
rect 23753 2595 23811 2601
rect 23842 2592 23848 2644
rect 23900 2632 23906 2644
rect 28626 2632 28632 2644
rect 23900 2604 28488 2632
rect 28587 2604 28632 2632
rect 23900 2592 23906 2604
rect 2774 2564 2780 2576
rect 1412 2536 2780 2564
rect 1412 2505 1440 2536
rect 2774 2524 2780 2536
rect 2832 2524 2838 2576
rect 15194 2564 15200 2576
rect 5276 2536 15200 2564
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1397 2459 1455 2465
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2866 2496 2872 2508
rect 2827 2468 2872 2496
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 5276 2505 5304 2536
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 20533 2567 20591 2573
rect 20533 2533 20545 2567
rect 20579 2564 20591 2567
rect 22646 2564 22652 2576
rect 20579 2536 22652 2564
rect 20579 2533 20591 2536
rect 20533 2527 20591 2533
rect 22646 2524 22652 2536
rect 22704 2524 22710 2576
rect 22925 2567 22983 2573
rect 22925 2533 22937 2567
rect 22971 2564 22983 2567
rect 24394 2564 24400 2576
rect 22971 2536 24400 2564
rect 22971 2533 22983 2536
rect 22925 2527 22983 2533
rect 24394 2524 24400 2536
rect 24452 2524 24458 2576
rect 25406 2564 25412 2576
rect 24504 2536 25412 2564
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2465 5319 2499
rect 5261 2459 5319 2465
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 6822 2496 6828 2508
rect 6595 2468 6828 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 6972 2468 7021 2496
rect 6972 2456 6978 2468
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 18509 2499 18567 2505
rect 18509 2496 18521 2499
rect 7009 2459 7067 2465
rect 17788 2468 18521 2496
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 2792 2400 3801 2428
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 2792 2360 2820 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5166 2428 5172 2440
rect 5031 2400 5172 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 17788 2437 17816 2468
rect 18509 2465 18521 2468
rect 18555 2465 18567 2499
rect 18509 2459 18567 2465
rect 21634 2456 21640 2508
rect 21692 2496 21698 2508
rect 24504 2496 24532 2536
rect 25406 2524 25412 2536
rect 25464 2524 25470 2576
rect 28460 2564 28488 2604
rect 28626 2592 28632 2604
rect 28684 2592 28690 2644
rect 38286 2632 38292 2644
rect 38247 2604 38292 2632
rect 38286 2592 38292 2604
rect 38344 2592 38350 2644
rect 39114 2592 39120 2644
rect 39172 2632 39178 2644
rect 39209 2635 39267 2641
rect 39209 2632 39221 2635
rect 39172 2604 39221 2632
rect 39172 2592 39178 2604
rect 39209 2601 39221 2604
rect 39255 2601 39267 2635
rect 39209 2595 39267 2601
rect 39298 2592 39304 2644
rect 39356 2632 39362 2644
rect 40405 2635 40463 2641
rect 40405 2632 40417 2635
rect 39356 2604 40417 2632
rect 39356 2592 39362 2604
rect 40405 2601 40417 2604
rect 40451 2601 40463 2635
rect 40405 2595 40463 2601
rect 43533 2635 43591 2641
rect 43533 2601 43545 2635
rect 43579 2632 43591 2635
rect 43714 2632 43720 2644
rect 43579 2604 43720 2632
rect 43579 2601 43591 2604
rect 43533 2595 43591 2601
rect 43714 2592 43720 2604
rect 43772 2592 43778 2644
rect 44358 2632 44364 2644
rect 44319 2604 44364 2632
rect 44358 2592 44364 2604
rect 44416 2592 44422 2644
rect 45557 2567 45615 2573
rect 45557 2564 45569 2567
rect 25516 2536 28396 2564
rect 28460 2536 45569 2564
rect 24670 2496 24676 2508
rect 21692 2468 24532 2496
rect 24631 2468 24676 2496
rect 21692 2456 21698 2468
rect 24670 2456 24676 2468
rect 24728 2456 24734 2508
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15528 2400 15761 2428
rect 15528 2388 15534 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2397 17831 2431
rect 17773 2391 17831 2397
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 2648 2332 2820 2360
rect 6733 2363 6791 2369
rect 2648 2320 2654 2332
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 7466 2360 7472 2372
rect 6779 2332 7472 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 7466 2320 7472 2332
rect 7524 2320 7530 2372
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 8444 2332 9413 2360
rect 8444 2320 8450 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9401 2323 9459 2329
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16172 2332 17141 2360
rect 16172 2320 16178 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 18432 2360 18460 2391
rect 19058 2388 19064 2440
rect 19116 2428 19122 2440
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 19116 2400 19257 2428
rect 19116 2388 19122 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 21913 2431 21971 2437
rect 21913 2428 21925 2431
rect 21315 2400 21925 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 21913 2397 21925 2400
rect 21959 2397 21971 2431
rect 23014 2428 23020 2440
rect 22975 2400 23020 2428
rect 21913 2391 21971 2397
rect 23014 2388 23020 2400
rect 23072 2388 23078 2440
rect 23658 2428 23664 2440
rect 23619 2400 23664 2428
rect 23658 2388 23664 2400
rect 23716 2388 23722 2440
rect 19337 2363 19395 2369
rect 19337 2360 19349 2363
rect 18432 2332 19349 2360
rect 17129 2323 17187 2329
rect 19337 2329 19349 2332
rect 19383 2329 19395 2363
rect 19337 2323 19395 2329
rect 20349 2363 20407 2369
rect 20349 2329 20361 2363
rect 20395 2360 20407 2363
rect 20622 2360 20628 2372
rect 20395 2332 20628 2360
rect 20395 2329 20407 2332
rect 20349 2323 20407 2329
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 21085 2363 21143 2369
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 24765 2363 24823 2369
rect 21131 2332 21956 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 21928 2304 21956 2332
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 25516 2360 25544 2536
rect 25682 2496 25688 2508
rect 25643 2468 25688 2496
rect 25682 2456 25688 2468
rect 25740 2456 25746 2508
rect 27154 2456 27160 2508
rect 27212 2496 27218 2508
rect 27249 2499 27307 2505
rect 27249 2496 27261 2499
rect 27212 2468 27261 2496
rect 27212 2456 27218 2468
rect 27249 2465 27261 2468
rect 27295 2465 27307 2499
rect 28368 2496 28396 2536
rect 45557 2533 45569 2536
rect 45603 2533 45615 2567
rect 45557 2527 45615 2533
rect 30006 2496 30012 2508
rect 28368 2468 29868 2496
rect 29967 2468 30012 2496
rect 27249 2459 27307 2465
rect 25590 2388 25596 2440
rect 25648 2428 25654 2440
rect 25648 2400 26372 2428
rect 25648 2388 25654 2400
rect 24811 2332 25544 2360
rect 26237 2363 26295 2369
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 26237 2329 26249 2363
rect 26283 2329 26295 2363
rect 26237 2323 26295 2329
rect 3970 2292 3976 2304
rect 3931 2264 3976 2292
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 9674 2292 9680 2304
rect 9635 2264 9680 2292
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 21910 2252 21916 2304
rect 21968 2252 21974 2304
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 26252 2292 26280 2323
rect 26344 2301 26372 2400
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26476 2400 26985 2428
rect 26476 2388 26482 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29840 2428 29868 2468
rect 30006 2456 30012 2468
rect 30064 2456 30070 2508
rect 35805 2499 35863 2505
rect 35805 2496 35817 2499
rect 30116 2468 35817 2496
rect 30116 2428 30144 2468
rect 35805 2465 35817 2468
rect 35851 2465 35863 2499
rect 35805 2459 35863 2465
rect 41325 2499 41383 2505
rect 41325 2465 41337 2499
rect 41371 2496 41383 2499
rect 41506 2496 41512 2508
rect 41371 2468 41512 2496
rect 41371 2465 41383 2468
rect 41325 2459 41383 2465
rect 41506 2456 41512 2468
rect 41564 2456 41570 2508
rect 43073 2499 43131 2505
rect 43073 2465 43085 2499
rect 43119 2496 43131 2499
rect 46106 2496 46112 2508
rect 43119 2468 46112 2496
rect 43119 2465 43131 2468
rect 43073 2459 43131 2465
rect 46106 2456 46112 2468
rect 46164 2456 46170 2508
rect 46201 2499 46259 2505
rect 46201 2465 46213 2499
rect 46247 2496 46259 2499
rect 47026 2496 47032 2508
rect 46247 2468 47032 2496
rect 46247 2465 46259 2468
rect 46201 2459 46259 2465
rect 47026 2456 47032 2468
rect 47084 2456 47090 2508
rect 29840 2400 30144 2428
rect 29733 2391 29791 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35492 2400 35541 2428
rect 35492 2388 35498 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 38010 2388 38016 2440
rect 38068 2428 38074 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 38068 2400 38117 2428
rect 38068 2388 38074 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 39117 2431 39175 2437
rect 39117 2397 39129 2431
rect 39163 2428 39175 2431
rect 40034 2428 40040 2440
rect 39163 2400 40040 2428
rect 39163 2397 39175 2400
rect 39117 2391 39175 2397
rect 40034 2388 40040 2400
rect 40092 2388 40098 2440
rect 41049 2431 41107 2437
rect 41049 2397 41061 2431
rect 41095 2428 41107 2431
rect 41230 2428 41236 2440
rect 41095 2400 41236 2428
rect 41095 2397 41107 2400
rect 41049 2391 41107 2397
rect 41230 2388 41236 2400
rect 41288 2388 41294 2440
rect 43717 2431 43775 2437
rect 43717 2397 43729 2431
rect 43763 2428 43775 2431
rect 43806 2428 43812 2440
rect 43763 2400 43812 2428
rect 43763 2397 43775 2400
rect 43717 2391 43775 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 44174 2428 44180 2440
rect 44135 2400 44180 2428
rect 44174 2388 44180 2400
rect 44232 2388 44238 2440
rect 46290 2388 46296 2440
rect 46348 2428 46354 2440
rect 46477 2431 46535 2437
rect 46477 2428 46489 2431
rect 46348 2400 46489 2428
rect 46348 2388 46354 2400
rect 46477 2397 46489 2400
rect 46523 2397 46535 2431
rect 46477 2391 46535 2397
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28537 2363 28595 2369
rect 28537 2360 28549 2363
rect 28408 2332 28549 2360
rect 28408 2320 28414 2332
rect 28537 2329 28549 2332
rect 28583 2329 28595 2363
rect 28537 2323 28595 2329
rect 39298 2320 39304 2372
rect 39356 2360 39362 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39356 2332 40325 2360
rect 39356 2320 39362 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 42889 2363 42947 2369
rect 42889 2360 42901 2363
rect 40644 2332 42901 2360
rect 40644 2320 40650 2332
rect 42889 2329 42901 2332
rect 42935 2329 42947 2363
rect 45373 2363 45431 2369
rect 42889 2323 42947 2329
rect 42996 2332 44496 2360
rect 24544 2264 26280 2292
rect 26329 2295 26387 2301
rect 24544 2252 24550 2264
rect 26329 2261 26341 2295
rect 26375 2261 26387 2295
rect 26329 2255 26387 2261
rect 31570 2252 31576 2304
rect 31628 2292 31634 2304
rect 42996 2292 43024 2332
rect 31628 2264 43024 2292
rect 44468 2292 44496 2332
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46382 2360 46388 2372
rect 45419 2332 46388 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46382 2320 46388 2332
rect 46440 2320 46446 2372
rect 47765 2363 47823 2369
rect 47765 2329 47777 2363
rect 47811 2360 47823 2363
rect 47946 2360 47952 2372
rect 47811 2332 47952 2360
rect 47811 2329 47823 2332
rect 47765 2323 47823 2329
rect 47946 2320 47952 2332
rect 48004 2320 48010 2372
rect 47857 2295 47915 2301
rect 47857 2292 47869 2295
rect 44468 2264 47869 2292
rect 31628 2252 31634 2264
rect 47857 2261 47869 2264
rect 47903 2261 47915 2295
rect 47857 2255 47915 2261
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 9674 2048 9680 2100
rect 9732 2088 9738 2100
rect 25038 2088 25044 2100
rect 9732 2060 25044 2088
rect 9732 2048 9738 2060
rect 25038 2048 25044 2060
rect 25096 2048 25102 2100
rect 44174 484 44180 536
rect 44232 524 44238 536
rect 46842 524 46848 536
rect 44232 496 46848 524
rect 44232 484 44238 496
rect 46842 484 46848 496
rect 46900 484 46906 536
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 29368 47200 29420 47252
rect 17776 47132 17828 47184
rect 20260 47132 20312 47184
rect 11612 47064 11664 47116
rect 20076 47107 20128 47116
rect 20076 47073 20085 47107
rect 20085 47073 20119 47107
rect 20119 47073 20128 47107
rect 20076 47064 20128 47073
rect 30748 47107 30800 47116
rect 1952 47039 2004 47048
rect 1952 47005 1961 47039
rect 1961 47005 1995 47039
rect 1995 47005 2004 47039
rect 1952 46996 2004 47005
rect 2596 46996 2648 47048
rect 3240 46996 3292 47048
rect 4804 47039 4856 47048
rect 4804 47005 4813 47039
rect 4813 47005 4847 47039
rect 4847 47005 4856 47039
rect 4804 46996 4856 47005
rect 5816 46996 5868 47048
rect 7104 46996 7156 47048
rect 9036 46996 9088 47048
rect 11980 47039 12032 47048
rect 11980 47005 11989 47039
rect 11989 47005 12023 47039
rect 12023 47005 12032 47039
rect 11980 46996 12032 47005
rect 12900 46996 12952 47048
rect 13820 46996 13872 47048
rect 16488 46996 16540 47048
rect 4068 46971 4120 46980
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 7840 46928 7892 46980
rect 9496 46928 9548 46980
rect 14648 46928 14700 46980
rect 18696 46996 18748 47048
rect 19984 46996 20036 47048
rect 30748 47073 30757 47107
rect 30757 47073 30791 47107
rect 30791 47073 30800 47107
rect 30748 47064 30800 47073
rect 45100 47064 45152 47116
rect 48320 47064 48372 47116
rect 20444 46996 20496 47048
rect 25688 47039 25740 47048
rect 25688 47005 25697 47039
rect 25697 47005 25731 47039
rect 25731 47005 25740 47039
rect 25688 46996 25740 47005
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 31116 46996 31168 47048
rect 38108 46996 38160 47048
rect 42524 46996 42576 47048
rect 45192 47039 45244 47048
rect 45192 47005 45201 47039
rect 45201 47005 45235 47039
rect 45235 47005 45244 47039
rect 45192 46996 45244 47005
rect 47676 46996 47728 47048
rect 22928 46928 22980 46980
rect 2136 46903 2188 46912
rect 2136 46869 2145 46903
rect 2145 46869 2179 46903
rect 2179 46869 2188 46903
rect 2136 46860 2188 46869
rect 2872 46903 2924 46912
rect 2872 46869 2881 46903
rect 2881 46869 2915 46903
rect 2915 46869 2924 46903
rect 2872 46860 2924 46869
rect 4896 46903 4948 46912
rect 4896 46869 4905 46903
rect 4905 46869 4939 46903
rect 4939 46869 4948 46903
rect 4896 46860 4948 46869
rect 6920 46903 6972 46912
rect 6920 46869 6929 46903
rect 6929 46869 6963 46903
rect 6963 46869 6972 46903
rect 6920 46860 6972 46869
rect 27068 46860 27120 46912
rect 27620 46860 27672 46912
rect 28264 46860 28316 46912
rect 39304 46860 39356 46912
rect 40408 46928 40460 46980
rect 42800 46971 42852 46980
rect 42800 46937 42809 46971
rect 42809 46937 42843 46971
rect 42843 46937 42852 46971
rect 42800 46928 42852 46937
rect 45376 46971 45428 46980
rect 45376 46937 45385 46971
rect 45385 46937 45419 46971
rect 45419 46937 45428 46971
rect 45376 46928 45428 46937
rect 41236 46860 41288 46912
rect 41788 46860 41840 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 2872 46588 2924 46640
rect 1400 46563 1452 46572
rect 1400 46529 1409 46563
rect 1409 46529 1443 46563
rect 1443 46529 1452 46563
rect 1400 46520 1452 46529
rect 12256 46520 12308 46572
rect 28264 46563 28316 46572
rect 28264 46529 28273 46563
rect 28273 46529 28307 46563
rect 28307 46529 28316 46563
rect 28264 46520 28316 46529
rect 38108 46563 38160 46572
rect 38108 46529 38117 46563
rect 38117 46529 38151 46563
rect 38151 46529 38160 46563
rect 38108 46520 38160 46529
rect 47860 46563 47912 46572
rect 47860 46529 47869 46563
rect 47869 46529 47903 46563
rect 47903 46529 47912 46563
rect 47860 46520 47912 46529
rect 13544 46452 13596 46504
rect 14188 46452 14240 46504
rect 14280 46495 14332 46504
rect 14280 46461 14289 46495
rect 14289 46461 14323 46495
rect 14323 46461 14332 46495
rect 14280 46452 14332 46461
rect 19616 46495 19668 46504
rect 19616 46461 19625 46495
rect 19625 46461 19659 46495
rect 19659 46461 19668 46495
rect 19616 46452 19668 46461
rect 20628 46495 20680 46504
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 24952 46452 25004 46504
rect 25780 46495 25832 46504
rect 25780 46461 25789 46495
rect 25789 46461 25823 46495
rect 25823 46461 25832 46495
rect 25780 46452 25832 46461
rect 38292 46495 38344 46504
rect 38292 46461 38301 46495
rect 38301 46461 38335 46495
rect 38335 46461 38344 46495
rect 38292 46452 38344 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 42616 46495 42668 46504
rect 42616 46461 42625 46495
rect 42625 46461 42659 46495
rect 42659 46461 42668 46495
rect 42616 46452 42668 46461
rect 42708 46452 42760 46504
rect 44272 46384 44324 46436
rect 46020 46452 46072 46504
rect 46848 46495 46900 46504
rect 46848 46461 46857 46495
rect 46857 46461 46891 46495
rect 46891 46461 46900 46495
rect 46848 46452 46900 46461
rect 46940 46384 46992 46436
rect 1676 46316 1728 46368
rect 2320 46359 2372 46368
rect 2320 46325 2329 46359
rect 2329 46325 2363 46359
rect 2363 46325 2372 46359
rect 2320 46316 2372 46325
rect 4620 46316 4672 46368
rect 10416 46316 10468 46368
rect 12532 46359 12584 46368
rect 12532 46325 12541 46359
rect 12541 46325 12575 46359
rect 12575 46325 12584 46359
rect 12532 46316 12584 46325
rect 20076 46316 20128 46368
rect 31668 46316 31720 46368
rect 41236 46359 41288 46368
rect 41236 46325 41245 46359
rect 41245 46325 41279 46359
rect 41279 46325 41288 46359
rect 41236 46316 41288 46325
rect 48044 46359 48096 46368
rect 48044 46325 48053 46359
rect 48053 46325 48087 46359
rect 48087 46325 48096 46359
rect 48044 46316 48096 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 13544 46155 13596 46164
rect 13544 46121 13553 46155
rect 13553 46121 13587 46155
rect 13587 46121 13596 46155
rect 13544 46112 13596 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 19616 46112 19668 46164
rect 24952 46112 25004 46164
rect 25412 46112 25464 46164
rect 38292 46155 38344 46164
rect 38292 46121 38301 46155
rect 38301 46121 38335 46155
rect 38335 46121 38344 46155
rect 38292 46112 38344 46121
rect 3884 46044 3936 46096
rect 2320 45976 2372 46028
rect 2780 46019 2832 46028
rect 2780 45985 2789 46019
rect 2789 45985 2823 46019
rect 2823 45985 2832 46019
rect 2780 45976 2832 45985
rect 4620 45976 4672 46028
rect 25136 46044 25188 46096
rect 10416 46019 10468 46028
rect 10416 45985 10425 46019
rect 10425 45985 10459 46019
rect 10459 45985 10468 46019
rect 10416 45976 10468 45985
rect 10968 45976 11020 46028
rect 20076 46019 20128 46028
rect 20076 45985 20085 46019
rect 20085 45985 20119 46019
rect 20119 45985 20128 46019
rect 20076 45976 20128 45985
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 25688 45976 25740 46028
rect 31668 46019 31720 46028
rect 31668 45985 31677 46019
rect 31677 45985 31711 46019
rect 31711 45985 31720 46019
rect 31668 45976 31720 45985
rect 32220 46019 32272 46028
rect 32220 45985 32229 46019
rect 32229 45985 32263 46019
rect 32263 45985 32272 46019
rect 32220 45976 32272 45985
rect 45928 46044 45980 46096
rect 41236 46019 41288 46028
rect 41236 45985 41245 46019
rect 41245 45985 41279 46019
rect 41279 45985 41288 46019
rect 41236 45976 41288 45985
rect 41880 46019 41932 46028
rect 41880 45985 41889 46019
rect 41889 45985 41923 46019
rect 41923 45985 41932 46019
rect 41880 45976 41932 45985
rect 47032 46019 47084 46028
rect 47032 45985 47041 46019
rect 47041 45985 47075 46019
rect 47075 45985 47084 46019
rect 47032 45976 47084 45985
rect 14096 45951 14148 45960
rect 14096 45917 14105 45951
rect 14105 45917 14139 45951
rect 14139 45917 14148 45951
rect 14096 45908 14148 45917
rect 18788 45908 18840 45960
rect 38200 45951 38252 45960
rect 2320 45840 2372 45892
rect 5080 45840 5132 45892
rect 10600 45883 10652 45892
rect 10600 45849 10609 45883
rect 10609 45849 10643 45883
rect 10643 45849 10652 45883
rect 10600 45840 10652 45849
rect 16672 45840 16724 45892
rect 38200 45917 38209 45951
rect 38209 45917 38243 45951
rect 38243 45917 38252 45951
rect 38200 45908 38252 45917
rect 43812 45908 43864 45960
rect 45744 45908 45796 45960
rect 46296 45951 46348 45960
rect 46296 45917 46305 45951
rect 46305 45917 46339 45951
rect 46339 45917 46348 45951
rect 46296 45908 46348 45917
rect 27068 45840 27120 45892
rect 32220 45840 32272 45892
rect 41420 45883 41472 45892
rect 41420 45849 41429 45883
rect 41429 45849 41463 45883
rect 41463 45849 41472 45883
rect 41420 45840 41472 45849
rect 46480 45883 46532 45892
rect 46480 45849 46489 45883
rect 46489 45849 46523 45883
rect 46523 45849 46532 45883
rect 46480 45840 46532 45849
rect 43996 45772 44048 45824
rect 46572 45772 46624 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 2320 45611 2372 45620
rect 2320 45577 2329 45611
rect 2329 45577 2363 45611
rect 2363 45577 2372 45611
rect 2320 45568 2372 45577
rect 5080 45611 5132 45620
rect 5080 45577 5089 45611
rect 5089 45577 5123 45611
rect 5123 45577 5132 45611
rect 5080 45568 5132 45577
rect 10600 45611 10652 45620
rect 10600 45577 10609 45611
rect 10609 45577 10643 45611
rect 10643 45577 10652 45611
rect 10600 45568 10652 45577
rect 32220 45611 32272 45620
rect 32220 45577 32229 45611
rect 32229 45577 32263 45611
rect 32263 45577 32272 45611
rect 32220 45568 32272 45577
rect 41420 45611 41472 45620
rect 41420 45577 41429 45611
rect 41429 45577 41463 45611
rect 41463 45577 41472 45611
rect 41420 45568 41472 45577
rect 2320 45432 2372 45484
rect 18328 45500 18380 45552
rect 25412 45543 25464 45552
rect 25412 45509 25421 45543
rect 25421 45509 25455 45543
rect 25455 45509 25464 45543
rect 25412 45500 25464 45509
rect 27068 45543 27120 45552
rect 27068 45509 27077 45543
rect 27077 45509 27111 45543
rect 27111 45509 27120 45543
rect 27068 45500 27120 45509
rect 45100 45543 45152 45552
rect 45100 45509 45109 45543
rect 45109 45509 45143 45543
rect 45143 45509 45152 45543
rect 45100 45500 45152 45509
rect 45376 45500 45428 45552
rect 16672 45432 16724 45484
rect 25320 45475 25372 45484
rect 25320 45441 25329 45475
rect 25329 45441 25363 45475
rect 25363 45441 25372 45475
rect 25320 45432 25372 45441
rect 26516 45432 26568 45484
rect 31944 45432 31996 45484
rect 41328 45475 41380 45484
rect 41328 45441 41337 45475
rect 41337 45441 41371 45475
rect 41371 45441 41380 45475
rect 41328 45432 41380 45441
rect 46204 45475 46256 45484
rect 46204 45441 46213 45475
rect 46213 45441 46247 45475
rect 46247 45441 46256 45475
rect 46204 45432 46256 45441
rect 47492 45432 47544 45484
rect 42708 45407 42760 45416
rect 42708 45373 42717 45407
rect 42717 45373 42751 45407
rect 42751 45373 42760 45407
rect 42708 45364 42760 45373
rect 43812 45364 43864 45416
rect 44088 45407 44140 45416
rect 44088 45373 44097 45407
rect 44097 45373 44131 45407
rect 44131 45373 44140 45407
rect 44088 45364 44140 45373
rect 45836 45364 45888 45416
rect 25320 45296 25372 45348
rect 45652 45296 45704 45348
rect 45100 45228 45152 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 42616 45024 42668 45076
rect 42800 45024 42852 45076
rect 43812 45067 43864 45076
rect 43812 45033 43821 45067
rect 43821 45033 43855 45067
rect 43855 45033 43864 45067
rect 43812 45024 43864 45033
rect 46480 45024 46532 45076
rect 46296 44956 46348 45008
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 29552 44820 29604 44872
rect 42064 44820 42116 44872
rect 43076 44863 43128 44872
rect 43076 44829 43085 44863
rect 43085 44829 43119 44863
rect 43119 44829 43128 44863
rect 43076 44820 43128 44829
rect 45652 44863 45704 44872
rect 28080 44684 28132 44736
rect 45652 44829 45661 44863
rect 45661 44829 45695 44863
rect 45695 44829 45704 44863
rect 45652 44820 45704 44829
rect 45744 44820 45796 44872
rect 46664 44752 46716 44804
rect 47584 44684 47636 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 46020 44523 46072 44532
rect 46020 44489 46029 44523
rect 46029 44489 46063 44523
rect 46063 44489 46072 44523
rect 46020 44480 46072 44489
rect 46664 44523 46716 44532
rect 46664 44489 46673 44523
rect 46673 44489 46707 44523
rect 46707 44489 46716 44523
rect 46664 44480 46716 44489
rect 28080 44455 28132 44464
rect 28080 44421 28089 44455
rect 28089 44421 28123 44455
rect 28123 44421 28132 44455
rect 28080 44412 28132 44421
rect 41328 44412 41380 44464
rect 42708 44344 42760 44396
rect 45744 44344 45796 44396
rect 45928 44387 45980 44396
rect 45928 44353 45937 44387
rect 45937 44353 45971 44387
rect 45971 44353 45980 44387
rect 45928 44344 45980 44353
rect 47492 44344 47544 44396
rect 3516 44276 3568 44328
rect 27712 44276 27764 44328
rect 38660 44319 38712 44328
rect 38660 44285 38669 44319
rect 38669 44285 38703 44319
rect 38703 44285 38712 44319
rect 38660 44276 38712 44285
rect 38844 44319 38896 44328
rect 38844 44285 38853 44319
rect 38853 44285 38887 44319
rect 38887 44285 38896 44319
rect 38844 44276 38896 44285
rect 40040 44319 40092 44328
rect 40040 44285 40049 44319
rect 40049 44285 40083 44319
rect 40083 44285 40092 44319
rect 40040 44276 40092 44285
rect 42524 44276 42576 44328
rect 29552 44140 29604 44192
rect 31944 44140 31996 44192
rect 47676 44183 47728 44192
rect 47676 44149 47685 44183
rect 47685 44149 47719 44183
rect 47719 44149 47728 44183
rect 47676 44140 47728 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 38844 43979 38896 43988
rect 38844 43945 38853 43979
rect 38853 43945 38887 43979
rect 38887 43945 38896 43979
rect 38844 43936 38896 43945
rect 47676 43800 47728 43852
rect 48136 43843 48188 43852
rect 48136 43809 48145 43843
rect 48145 43809 48179 43843
rect 48179 43809 48188 43843
rect 48136 43800 48188 43809
rect 26976 43732 27028 43784
rect 29552 43775 29604 43784
rect 29552 43741 29561 43775
rect 29561 43741 29595 43775
rect 29595 43741 29604 43775
rect 29552 43732 29604 43741
rect 38752 43775 38804 43784
rect 38752 43741 38761 43775
rect 38761 43741 38795 43775
rect 38795 43741 38804 43775
rect 38752 43732 38804 43741
rect 27620 43664 27672 43716
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 2136 43188 2188 43240
rect 25596 43256 25648 43308
rect 45192 43256 45244 43308
rect 46940 43299 46992 43308
rect 46940 43265 46949 43299
rect 46949 43265 46983 43299
rect 46983 43265 46992 43299
rect 46940 43256 46992 43265
rect 26976 43231 27028 43240
rect 26976 43197 26985 43231
rect 26985 43197 27019 43231
rect 27019 43197 27028 43231
rect 26976 43188 27028 43197
rect 28816 43231 28868 43240
rect 28816 43197 28825 43231
rect 28825 43197 28859 43231
rect 28859 43197 28868 43231
rect 28816 43188 28868 43197
rect 1584 43095 1636 43104
rect 1584 43061 1593 43095
rect 1593 43061 1627 43095
rect 1627 43061 1636 43095
rect 1584 43052 1636 43061
rect 38660 43052 38712 43104
rect 47768 43095 47820 43104
rect 47768 43061 47777 43095
rect 47777 43061 47811 43095
rect 47811 43061 47820 43095
rect 47768 43052 47820 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 47768 42712 47820 42764
rect 47676 42576 47728 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 47676 42347 47728 42356
rect 47676 42313 47685 42347
rect 47685 42313 47719 42347
rect 47719 42313 47728 42347
rect 47676 42304 47728 42313
rect 1584 42100 1636 42152
rect 45652 42168 45704 42220
rect 47308 42168 47360 42220
rect 47584 42211 47636 42220
rect 47584 42177 47593 42211
rect 47593 42177 47627 42211
rect 47627 42177 47636 42211
rect 47584 42168 47636 42177
rect 26700 42100 26752 42152
rect 28816 42143 28868 42152
rect 28816 42109 28825 42143
rect 28825 42109 28859 42143
rect 28859 42109 28868 42143
rect 28816 42100 28868 42109
rect 1400 41964 1452 42016
rect 46480 41964 46532 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 46480 41667 46532 41676
rect 46480 41633 46489 41667
rect 46489 41633 46523 41667
rect 46523 41633 46532 41667
rect 46480 41624 46532 41633
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 47768 41488 47820 41540
rect 48136 41531 48188 41540
rect 48136 41497 48145 41531
rect 48145 41497 48179 41531
rect 48179 41497 48188 41531
rect 48136 41488 48188 41497
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 14096 41080 14148 41132
rect 46204 41123 46256 41132
rect 46204 41089 46213 41123
rect 46213 41089 46247 41123
rect 46247 41089 46256 41123
rect 46204 41080 46256 41089
rect 47768 41123 47820 41132
rect 47768 41089 47777 41123
rect 47777 41089 47811 41123
rect 47811 41089 47820 41123
rect 47768 41080 47820 41089
rect 43812 41012 43864 41064
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47768 40536 47820 40588
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 2044 40443 2096 40452
rect 2044 40409 2053 40443
rect 2053 40409 2087 40443
rect 2087 40409 2096 40443
rect 2044 40400 2096 40409
rect 45560 40400 45612 40452
rect 48136 40443 48188 40452
rect 48136 40409 48145 40443
rect 48145 40409 48179 40443
rect 48179 40409 48188 40443
rect 48136 40400 48188 40409
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 18972 40103 19024 40112
rect 18972 40069 18981 40103
rect 18981 40069 19015 40103
rect 19015 40069 19024 40103
rect 18972 40060 19024 40069
rect 38200 40060 38252 40112
rect 18420 40035 18472 40044
rect 18420 40001 18429 40035
rect 18429 40001 18463 40035
rect 18463 40001 18472 40035
rect 18420 39992 18472 40001
rect 19156 39992 19208 40044
rect 25320 39992 25372 40044
rect 43812 40060 43864 40112
rect 46020 40060 46072 40112
rect 47768 40035 47820 40044
rect 47768 40001 47777 40035
rect 47777 40001 47811 40035
rect 47811 40001 47820 40035
rect 47768 39992 47820 40001
rect 43720 39967 43772 39976
rect 43720 39933 43729 39967
rect 43729 39933 43763 39967
rect 43763 39933 43772 39967
rect 43720 39924 43772 39933
rect 26976 39856 27028 39908
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 18328 39448 18380 39500
rect 22744 39491 22796 39500
rect 18420 39380 18472 39432
rect 22744 39457 22753 39491
rect 22753 39457 22787 39491
rect 22787 39457 22796 39491
rect 22744 39448 22796 39457
rect 47860 39448 47912 39500
rect 38752 39380 38804 39432
rect 39948 39380 40000 39432
rect 16672 39312 16724 39364
rect 17592 39312 17644 39364
rect 20628 39312 20680 39364
rect 42064 39312 42116 39364
rect 47676 39312 47728 39364
rect 48136 39355 48188 39364
rect 48136 39321 48145 39355
rect 48145 39321 48179 39355
rect 48179 39321 48188 39355
rect 48136 39312 48188 39321
rect 22192 39287 22244 39296
rect 22192 39253 22201 39287
rect 22201 39253 22235 39287
rect 22235 39253 22244 39287
rect 22192 39244 22244 39253
rect 22468 39244 22520 39296
rect 22652 39287 22704 39296
rect 22652 39253 22661 39287
rect 22661 39253 22695 39287
rect 22695 39253 22704 39287
rect 22652 39244 22704 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 22468 39040 22520 39092
rect 47676 39083 47728 39092
rect 47676 39049 47685 39083
rect 47685 39049 47719 39083
rect 47719 39049 47728 39083
rect 47676 39040 47728 39049
rect 22560 38972 22612 39024
rect 18420 38947 18472 38956
rect 18420 38913 18429 38947
rect 18429 38913 18463 38947
rect 18463 38913 18472 38947
rect 18420 38904 18472 38913
rect 26976 38904 27028 38956
rect 30196 38904 30248 38956
rect 45652 38947 45704 38956
rect 45652 38913 45661 38947
rect 45661 38913 45695 38947
rect 45695 38913 45704 38947
rect 45652 38904 45704 38913
rect 45836 38947 45888 38956
rect 45836 38913 45845 38947
rect 45845 38913 45879 38947
rect 45879 38913 45888 38947
rect 45836 38904 45888 38913
rect 46388 38947 46440 38956
rect 46388 38913 46397 38947
rect 46397 38913 46431 38947
rect 46431 38913 46440 38947
rect 46388 38904 46440 38913
rect 47676 38904 47728 38956
rect 19156 38879 19208 38888
rect 19156 38845 19165 38879
rect 19165 38845 19199 38879
rect 19199 38845 19208 38879
rect 19156 38836 19208 38845
rect 21824 38879 21876 38888
rect 21824 38845 21833 38879
rect 21833 38845 21867 38879
rect 21867 38845 21876 38879
rect 21824 38836 21876 38845
rect 22100 38879 22152 38888
rect 22100 38845 22109 38879
rect 22109 38845 22143 38879
rect 22143 38845 22152 38879
rect 46848 38879 46900 38888
rect 22100 38836 22152 38845
rect 46848 38845 46857 38879
rect 46857 38845 46891 38879
rect 46891 38845 46900 38879
rect 46848 38836 46900 38845
rect 24860 38700 24912 38752
rect 45560 38700 45612 38752
rect 46112 38700 46164 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 18420 38496 18472 38548
rect 22652 38496 22704 38548
rect 24492 38496 24544 38548
rect 26976 38539 27028 38548
rect 20904 38360 20956 38412
rect 21088 38428 21140 38480
rect 21824 38428 21876 38480
rect 23480 38403 23532 38412
rect 19984 38292 20036 38344
rect 21180 38292 21232 38344
rect 22192 38292 22244 38344
rect 23480 38369 23489 38403
rect 23489 38369 23523 38403
rect 23523 38369 23532 38403
rect 23480 38360 23532 38369
rect 25412 38360 25464 38412
rect 26976 38505 26985 38539
rect 26985 38505 27019 38539
rect 27019 38505 27028 38539
rect 26976 38496 27028 38505
rect 11980 38224 12032 38276
rect 17132 38156 17184 38208
rect 18696 38156 18748 38208
rect 20536 38156 20588 38208
rect 22100 38156 22152 38208
rect 23296 38199 23348 38208
rect 23296 38165 23305 38199
rect 23305 38165 23339 38199
rect 23339 38165 23348 38199
rect 46572 38496 46624 38548
rect 45836 38428 45888 38480
rect 24860 38267 24912 38276
rect 24860 38233 24869 38267
rect 24869 38233 24903 38267
rect 24903 38233 24912 38267
rect 24860 38224 24912 38233
rect 25320 38224 25372 38276
rect 23296 38156 23348 38165
rect 26148 38156 26200 38208
rect 26332 38199 26384 38208
rect 26332 38165 26341 38199
rect 26341 38165 26375 38199
rect 26375 38165 26384 38199
rect 26332 38156 26384 38165
rect 26424 38156 26476 38208
rect 45652 38292 45704 38344
rect 45928 38292 45980 38344
rect 47860 38267 47912 38276
rect 47860 38233 47869 38267
rect 47869 38233 47903 38267
rect 47903 38233 47912 38267
rect 47860 38224 47912 38233
rect 46112 38156 46164 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 22560 37952 22612 38004
rect 23296 37952 23348 38004
rect 24492 37995 24544 38004
rect 24492 37961 24501 37995
rect 24501 37961 24535 37995
rect 24535 37961 24544 37995
rect 24492 37952 24544 37961
rect 25320 37952 25372 38004
rect 26148 37952 26200 38004
rect 46020 37995 46072 38004
rect 17132 37927 17184 37936
rect 17132 37893 17141 37927
rect 17141 37893 17175 37927
rect 17175 37893 17184 37927
rect 17132 37884 17184 37893
rect 18144 37884 18196 37936
rect 20536 37884 20588 37936
rect 21180 37816 21232 37868
rect 22468 37816 22520 37868
rect 22652 37816 22704 37868
rect 23480 37816 23532 37868
rect 24584 37816 24636 37868
rect 24676 37816 24728 37868
rect 26332 37816 26384 37868
rect 16304 37748 16356 37800
rect 18604 37655 18656 37664
rect 18604 37621 18613 37655
rect 18613 37621 18647 37655
rect 18647 37621 18656 37655
rect 20536 37748 20588 37800
rect 22100 37748 22152 37800
rect 20904 37680 20956 37732
rect 24308 37680 24360 37732
rect 24492 37680 24544 37732
rect 18604 37612 18656 37621
rect 20812 37612 20864 37664
rect 21088 37612 21140 37664
rect 21272 37655 21324 37664
rect 21272 37621 21281 37655
rect 21281 37621 21315 37655
rect 21315 37621 21324 37655
rect 21272 37612 21324 37621
rect 26424 37791 26476 37800
rect 26424 37757 26433 37791
rect 26433 37757 26467 37791
rect 26467 37757 26476 37791
rect 26424 37748 26476 37757
rect 26884 37816 26936 37868
rect 29552 37816 29604 37868
rect 27528 37748 27580 37800
rect 28172 37791 28224 37800
rect 28172 37757 28181 37791
rect 28181 37757 28215 37791
rect 28215 37757 28224 37791
rect 28172 37748 28224 37757
rect 28908 37748 28960 37800
rect 26332 37680 26384 37732
rect 46020 37961 46029 37995
rect 46029 37961 46063 37995
rect 46063 37961 46072 37995
rect 46020 37952 46072 37961
rect 39948 37884 40000 37936
rect 45560 37884 45612 37936
rect 45744 37859 45796 37868
rect 45744 37825 45753 37859
rect 45753 37825 45787 37859
rect 45787 37825 45796 37859
rect 45744 37816 45796 37825
rect 46112 37859 46164 37868
rect 46112 37825 46121 37859
rect 46121 37825 46155 37859
rect 46155 37825 46164 37859
rect 46112 37816 46164 37825
rect 45928 37748 45980 37800
rect 46020 37680 46072 37732
rect 26148 37612 26200 37664
rect 27160 37655 27212 37664
rect 27160 37621 27169 37655
rect 27169 37621 27203 37655
rect 27203 37621 27212 37655
rect 27160 37612 27212 37621
rect 28264 37612 28316 37664
rect 29920 37655 29972 37664
rect 29920 37621 29929 37655
rect 29929 37621 29963 37655
rect 29963 37621 29972 37655
rect 29920 37612 29972 37621
rect 46480 37612 46532 37664
rect 47768 37655 47820 37664
rect 47768 37621 47777 37655
rect 47777 37621 47811 37655
rect 47811 37621 47820 37655
rect 47768 37612 47820 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 9496 37408 9548 37460
rect 28908 37451 28960 37460
rect 2044 37340 2096 37392
rect 18696 37383 18748 37392
rect 18236 37315 18288 37324
rect 18236 37281 18245 37315
rect 18245 37281 18279 37315
rect 18279 37281 18288 37315
rect 18236 37272 18288 37281
rect 18696 37349 18705 37383
rect 18705 37349 18739 37383
rect 18739 37349 18748 37383
rect 18696 37340 18748 37349
rect 19984 37340 20036 37392
rect 20536 37383 20588 37392
rect 20536 37349 20545 37383
rect 20545 37349 20579 37383
rect 20579 37349 20588 37383
rect 20536 37340 20588 37349
rect 22100 37383 22152 37392
rect 22100 37349 22109 37383
rect 22109 37349 22143 37383
rect 22143 37349 22152 37383
rect 22100 37340 22152 37349
rect 21272 37272 21324 37324
rect 22652 37340 22704 37392
rect 1768 37204 1820 37256
rect 18512 37204 18564 37256
rect 19800 37247 19852 37256
rect 19800 37213 19809 37247
rect 19809 37213 19843 37247
rect 19843 37213 19852 37247
rect 19800 37204 19852 37213
rect 19340 37136 19392 37188
rect 20168 37247 20220 37256
rect 20168 37213 20177 37247
rect 20177 37213 20211 37247
rect 20211 37213 20220 37247
rect 20168 37204 20220 37213
rect 20352 37247 20404 37256
rect 20352 37213 20361 37247
rect 20361 37213 20395 37247
rect 20395 37213 20404 37247
rect 22284 37272 22336 37324
rect 27160 37272 27212 37324
rect 28908 37417 28917 37451
rect 28917 37417 28951 37451
rect 28951 37417 28960 37451
rect 28908 37408 28960 37417
rect 29552 37408 29604 37460
rect 45744 37451 45796 37460
rect 45744 37417 45753 37451
rect 45753 37417 45787 37451
rect 45787 37417 45796 37451
rect 45744 37408 45796 37417
rect 46020 37340 46072 37392
rect 46848 37340 46900 37392
rect 20352 37204 20404 37213
rect 28356 37247 28408 37256
rect 22284 37136 22336 37188
rect 22652 37179 22704 37188
rect 22652 37145 22661 37179
rect 22661 37145 22695 37179
rect 22695 37145 22704 37179
rect 22652 37136 22704 37145
rect 22744 37136 22796 37188
rect 26516 37136 26568 37188
rect 26884 37136 26936 37188
rect 28356 37213 28365 37247
rect 28365 37213 28399 37247
rect 28399 37213 28408 37247
rect 28356 37204 28408 37213
rect 29736 37272 29788 37324
rect 29920 37272 29972 37324
rect 45560 37272 45612 37324
rect 45744 37272 45796 37324
rect 46480 37315 46532 37324
rect 46480 37281 46489 37315
rect 46489 37281 46523 37315
rect 46523 37281 46532 37315
rect 46480 37272 46532 37281
rect 48136 37315 48188 37324
rect 48136 37281 48145 37315
rect 48145 37281 48179 37315
rect 48179 37281 48188 37315
rect 48136 37272 48188 37281
rect 28724 37247 28776 37256
rect 28724 37213 28733 37247
rect 28733 37213 28767 37247
rect 28767 37213 28776 37247
rect 28724 37204 28776 37213
rect 29184 37136 29236 37188
rect 21732 37111 21784 37120
rect 21732 37077 21741 37111
rect 21741 37077 21775 37111
rect 21775 37077 21784 37111
rect 21732 37068 21784 37077
rect 23204 37068 23256 37120
rect 26976 37068 27028 37120
rect 30748 37204 30800 37256
rect 45652 37247 45704 37256
rect 45652 37213 45661 37247
rect 45661 37213 45695 37247
rect 45695 37213 45704 37247
rect 45652 37204 45704 37213
rect 45836 37247 45888 37256
rect 45836 37213 45845 37247
rect 45845 37213 45879 37247
rect 45879 37213 45888 37247
rect 45836 37204 45888 37213
rect 47768 37136 47820 37188
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 18144 36864 18196 36916
rect 19984 36864 20036 36916
rect 23848 36864 23900 36916
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 17684 36771 17736 36780
rect 17684 36737 17693 36771
rect 17693 36737 17727 36771
rect 17727 36737 17736 36771
rect 17684 36728 17736 36737
rect 17776 36728 17828 36780
rect 18696 36728 18748 36780
rect 21732 36728 21784 36780
rect 24676 36728 24728 36780
rect 28172 36728 28224 36780
rect 28540 36771 28592 36780
rect 28540 36737 28549 36771
rect 28549 36737 28583 36771
rect 28583 36737 28592 36771
rect 28540 36728 28592 36737
rect 30748 36771 30800 36780
rect 30748 36737 30757 36771
rect 30757 36737 30791 36771
rect 30791 36737 30800 36771
rect 30748 36728 30800 36737
rect 2228 36660 2280 36712
rect 2780 36703 2832 36712
rect 2780 36669 2789 36703
rect 2789 36669 2823 36703
rect 2823 36669 2832 36703
rect 2780 36660 2832 36669
rect 29460 36660 29512 36712
rect 23388 36592 23440 36644
rect 26976 36592 27028 36644
rect 23480 36524 23532 36576
rect 24400 36567 24452 36576
rect 24400 36533 24409 36567
rect 24409 36533 24443 36567
rect 24443 36533 24452 36567
rect 24400 36524 24452 36533
rect 30288 36567 30340 36576
rect 30288 36533 30297 36567
rect 30297 36533 30331 36567
rect 30331 36533 30340 36567
rect 30288 36524 30340 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2228 36363 2280 36372
rect 2228 36329 2237 36363
rect 2237 36329 2271 36363
rect 2271 36329 2280 36363
rect 2228 36320 2280 36329
rect 20352 36252 20404 36304
rect 19248 36184 19300 36236
rect 22928 36184 22980 36236
rect 23572 36184 23624 36236
rect 2136 36159 2188 36168
rect 2136 36125 2145 36159
rect 2145 36125 2179 36159
rect 2179 36125 2188 36159
rect 2136 36116 2188 36125
rect 15660 36116 15712 36168
rect 16304 36159 16356 36168
rect 16304 36125 16313 36159
rect 16313 36125 16347 36159
rect 16347 36125 16356 36159
rect 16304 36116 16356 36125
rect 22468 36116 22520 36168
rect 22744 36116 22796 36168
rect 23296 36159 23348 36168
rect 17316 36048 17368 36100
rect 23296 36125 23305 36159
rect 23305 36125 23339 36159
rect 23339 36125 23348 36159
rect 23296 36116 23348 36125
rect 25412 36227 25464 36236
rect 25412 36193 25421 36227
rect 25421 36193 25455 36227
rect 25455 36193 25464 36227
rect 25412 36184 25464 36193
rect 26424 36184 26476 36236
rect 23572 36048 23624 36100
rect 27068 36048 27120 36100
rect 27896 36048 27948 36100
rect 29736 36159 29788 36168
rect 29736 36125 29745 36159
rect 29745 36125 29779 36159
rect 29779 36125 29788 36159
rect 29736 36116 29788 36125
rect 29920 36159 29972 36168
rect 29920 36125 29929 36159
rect 29929 36125 29963 36159
rect 29963 36125 29972 36159
rect 29920 36116 29972 36125
rect 30012 36159 30064 36168
rect 30012 36125 30021 36159
rect 30021 36125 30055 36159
rect 30055 36125 30064 36159
rect 30012 36116 30064 36125
rect 28724 36048 28776 36100
rect 29644 36048 29696 36100
rect 18052 36023 18104 36032
rect 18052 35989 18061 36023
rect 18061 35989 18095 36023
rect 18095 35989 18104 36023
rect 18052 35980 18104 35989
rect 19064 35980 19116 36032
rect 22928 35980 22980 36032
rect 23296 35980 23348 36032
rect 23664 35980 23716 36032
rect 27160 36023 27212 36032
rect 27160 35989 27169 36023
rect 27169 35989 27203 36023
rect 27203 35989 27212 36023
rect 27160 35980 27212 35989
rect 28080 35980 28132 36032
rect 29000 35980 29052 36032
rect 29828 35980 29880 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 17316 35819 17368 35828
rect 17316 35785 17325 35819
rect 17325 35785 17359 35819
rect 17359 35785 17368 35819
rect 17316 35776 17368 35785
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 16672 35640 16724 35692
rect 17684 35640 17736 35692
rect 17868 35683 17920 35692
rect 17868 35649 17877 35683
rect 17877 35649 17911 35683
rect 17911 35649 17920 35683
rect 17868 35640 17920 35649
rect 18052 35683 18104 35692
rect 18052 35649 18061 35683
rect 18061 35649 18095 35683
rect 18095 35649 18104 35683
rect 18052 35640 18104 35649
rect 19064 35708 19116 35760
rect 19248 35776 19300 35828
rect 23756 35776 23808 35828
rect 24676 35776 24728 35828
rect 27068 35819 27120 35828
rect 27068 35785 27077 35819
rect 27077 35785 27111 35819
rect 27111 35785 27120 35819
rect 27068 35776 27120 35785
rect 29460 35819 29512 35828
rect 19340 35708 19392 35760
rect 23664 35751 23716 35760
rect 23664 35717 23673 35751
rect 23673 35717 23707 35751
rect 23707 35717 23716 35751
rect 23664 35708 23716 35717
rect 24400 35708 24452 35760
rect 28264 35708 28316 35760
rect 20352 35640 20404 35692
rect 22468 35683 22520 35692
rect 22468 35649 22477 35683
rect 22477 35649 22511 35683
rect 22511 35649 22520 35683
rect 22468 35640 22520 35649
rect 22560 35683 22612 35692
rect 22560 35649 22569 35683
rect 22569 35649 22603 35683
rect 22603 35649 22612 35683
rect 22836 35683 22888 35692
rect 22560 35640 22612 35649
rect 22836 35649 22845 35683
rect 22845 35649 22879 35683
rect 22879 35649 22888 35683
rect 22836 35640 22888 35649
rect 26976 35683 27028 35692
rect 26976 35649 26985 35683
rect 26985 35649 27019 35683
rect 27019 35649 27028 35683
rect 26976 35640 27028 35649
rect 27804 35640 27856 35692
rect 27988 35683 28040 35692
rect 27988 35649 27997 35683
rect 27997 35649 28031 35683
rect 28031 35649 28040 35683
rect 27988 35640 28040 35649
rect 29460 35785 29469 35819
rect 29469 35785 29503 35819
rect 29503 35785 29512 35819
rect 29460 35776 29512 35785
rect 29552 35776 29604 35828
rect 43996 35776 44048 35828
rect 29092 35708 29144 35760
rect 19064 35615 19116 35624
rect 19064 35581 19073 35615
rect 19073 35581 19107 35615
rect 19107 35581 19116 35615
rect 19064 35572 19116 35581
rect 20720 35572 20772 35624
rect 22376 35572 22428 35624
rect 27620 35572 27672 35624
rect 29000 35683 29052 35692
rect 29000 35649 29009 35683
rect 29009 35649 29043 35683
rect 29043 35649 29052 35683
rect 29644 35708 29696 35760
rect 29000 35640 29052 35649
rect 29920 35683 29972 35692
rect 29920 35649 29929 35683
rect 29929 35649 29963 35683
rect 29963 35649 29972 35683
rect 30932 35683 30984 35692
rect 29920 35640 29972 35649
rect 29460 35572 29512 35624
rect 29736 35572 29788 35624
rect 30932 35649 30941 35683
rect 30941 35649 30975 35683
rect 30975 35649 30984 35683
rect 30932 35640 30984 35649
rect 31852 35640 31904 35692
rect 31760 35572 31812 35624
rect 19800 35504 19852 35556
rect 27804 35504 27856 35556
rect 31300 35547 31352 35556
rect 31300 35513 31309 35547
rect 31309 35513 31343 35547
rect 31343 35513 31352 35547
rect 31300 35504 31352 35513
rect 1492 35436 1544 35488
rect 18328 35436 18380 35488
rect 22284 35479 22336 35488
rect 22284 35445 22293 35479
rect 22293 35445 22327 35479
rect 22327 35445 22336 35479
rect 22284 35436 22336 35445
rect 29092 35436 29144 35488
rect 29736 35436 29788 35488
rect 30012 35436 30064 35488
rect 30932 35436 30984 35488
rect 32128 35436 32180 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 18236 35275 18288 35284
rect 18236 35241 18245 35275
rect 18245 35241 18279 35275
rect 18279 35241 18288 35275
rect 18236 35232 18288 35241
rect 19800 35275 19852 35284
rect 19800 35241 19809 35275
rect 19809 35241 19843 35275
rect 19843 35241 19852 35275
rect 19800 35232 19852 35241
rect 22192 35232 22244 35284
rect 22560 35232 22612 35284
rect 24952 35232 25004 35284
rect 18052 35096 18104 35148
rect 18420 35096 18472 35148
rect 19064 35096 19116 35148
rect 23572 35164 23624 35216
rect 26424 35232 26476 35284
rect 27160 35232 27212 35284
rect 28264 35232 28316 35284
rect 29184 35232 29236 35284
rect 29644 35275 29696 35284
rect 29644 35241 29653 35275
rect 29653 35241 29687 35275
rect 29687 35241 29696 35275
rect 29644 35232 29696 35241
rect 27068 35164 27120 35216
rect 27804 35164 27856 35216
rect 20720 35139 20772 35148
rect 20720 35105 20729 35139
rect 20729 35105 20763 35139
rect 20763 35105 20772 35139
rect 20720 35096 20772 35105
rect 21088 35096 21140 35148
rect 25964 35096 26016 35148
rect 27160 35096 27212 35148
rect 27344 35139 27396 35148
rect 27344 35105 27353 35139
rect 27353 35105 27387 35139
rect 27387 35105 27396 35139
rect 27344 35096 27396 35105
rect 17868 35028 17920 35080
rect 18512 35071 18564 35080
rect 18052 34960 18104 35012
rect 18512 35037 18521 35071
rect 18521 35037 18555 35071
rect 18555 35037 18564 35071
rect 18512 35028 18564 35037
rect 18604 35028 18656 35080
rect 23112 35071 23164 35080
rect 23112 35037 23121 35071
rect 23121 35037 23155 35071
rect 23155 35037 23164 35071
rect 23112 35028 23164 35037
rect 23388 35071 23440 35080
rect 23388 35037 23397 35071
rect 23397 35037 23431 35071
rect 23431 35037 23440 35071
rect 23388 35028 23440 35037
rect 24676 35028 24728 35080
rect 27436 35028 27488 35080
rect 27528 35071 27580 35080
rect 27528 35037 27537 35071
rect 27537 35037 27571 35071
rect 27571 35037 27580 35071
rect 27528 35028 27580 35037
rect 20352 34960 20404 35012
rect 20996 35003 21048 35012
rect 20996 34969 21005 35003
rect 21005 34969 21039 35003
rect 21039 34969 21048 35003
rect 20996 34960 21048 34969
rect 21456 34960 21508 35012
rect 19064 34892 19116 34944
rect 19984 34892 20036 34944
rect 23204 34960 23256 35012
rect 25320 34960 25372 35012
rect 27252 35003 27304 35012
rect 22468 34892 22520 34944
rect 25780 34892 25832 34944
rect 27252 34969 27261 35003
rect 27261 34969 27295 35003
rect 27295 34969 27304 35003
rect 27252 34960 27304 34969
rect 28540 35096 28592 35148
rect 29736 35139 29788 35148
rect 29736 35105 29745 35139
rect 29745 35105 29779 35139
rect 29779 35105 29788 35139
rect 29736 35096 29788 35105
rect 29644 35028 29696 35080
rect 30288 35028 30340 35080
rect 48136 35071 48188 35080
rect 48136 35037 48145 35071
rect 48145 35037 48179 35071
rect 48179 35037 48188 35071
rect 48136 35028 48188 35037
rect 30104 34960 30156 35012
rect 31024 34960 31076 35012
rect 32128 34960 32180 35012
rect 28632 34892 28684 34944
rect 32864 34935 32916 34944
rect 32864 34901 32873 34935
rect 32873 34901 32907 34935
rect 32907 34901 32916 34935
rect 32864 34892 32916 34901
rect 47124 34892 47176 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 18604 34731 18656 34740
rect 18604 34697 18613 34731
rect 18613 34697 18647 34731
rect 18647 34697 18656 34731
rect 18604 34688 18656 34697
rect 21088 34688 21140 34740
rect 21456 34688 21508 34740
rect 24952 34731 25004 34740
rect 24952 34697 24961 34731
rect 24961 34697 24995 34731
rect 24995 34697 25004 34731
rect 24952 34688 25004 34697
rect 27436 34688 27488 34740
rect 17500 34620 17552 34672
rect 18696 34620 18748 34672
rect 19064 34663 19116 34672
rect 19064 34629 19073 34663
rect 19073 34629 19107 34663
rect 19107 34629 19116 34663
rect 19064 34620 19116 34629
rect 17132 34595 17184 34604
rect 17132 34561 17141 34595
rect 17141 34561 17175 34595
rect 17175 34561 17184 34595
rect 17132 34552 17184 34561
rect 17960 34552 18012 34604
rect 18328 34595 18380 34604
rect 18328 34561 18337 34595
rect 18337 34561 18371 34595
rect 18371 34561 18380 34595
rect 18328 34552 18380 34561
rect 18880 34552 18932 34604
rect 19984 34620 20036 34672
rect 20352 34552 20404 34604
rect 22560 34620 22612 34672
rect 25964 34663 26016 34672
rect 25964 34629 25973 34663
rect 25973 34629 26007 34663
rect 26007 34629 26016 34663
rect 25964 34620 26016 34629
rect 21088 34595 21140 34604
rect 21088 34561 21097 34595
rect 21097 34561 21131 34595
rect 21131 34561 21140 34595
rect 21088 34552 21140 34561
rect 22100 34552 22152 34604
rect 23112 34552 23164 34604
rect 24676 34552 24728 34604
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 26148 34595 26200 34604
rect 26148 34561 26157 34595
rect 26157 34561 26191 34595
rect 26191 34561 26200 34595
rect 26148 34552 26200 34561
rect 27344 34620 27396 34672
rect 27620 34620 27672 34672
rect 31760 34688 31812 34740
rect 32128 34688 32180 34740
rect 18052 34416 18104 34468
rect 19248 34416 19300 34468
rect 22468 34484 22520 34536
rect 27160 34552 27212 34604
rect 27896 34595 27948 34604
rect 27896 34561 27905 34595
rect 27905 34561 27939 34595
rect 27939 34561 27948 34595
rect 27896 34552 27948 34561
rect 30932 34620 30984 34672
rect 28356 34552 28408 34604
rect 28632 34595 28684 34604
rect 28632 34561 28641 34595
rect 28641 34561 28675 34595
rect 28675 34561 28684 34595
rect 28632 34552 28684 34561
rect 29920 34552 29972 34604
rect 30104 34552 30156 34604
rect 32864 34620 32916 34672
rect 28356 34416 28408 34468
rect 30288 34484 30340 34536
rect 48136 34595 48188 34604
rect 48136 34561 48145 34595
rect 48145 34561 48179 34595
rect 48179 34561 48188 34595
rect 48136 34552 48188 34561
rect 46572 34484 46624 34536
rect 16948 34391 17000 34400
rect 16948 34357 16957 34391
rect 16957 34357 16991 34391
rect 16991 34357 17000 34391
rect 16948 34348 17000 34357
rect 18420 34391 18472 34400
rect 18420 34357 18429 34391
rect 18429 34357 18463 34391
rect 18463 34357 18472 34391
rect 18420 34348 18472 34357
rect 21732 34348 21784 34400
rect 26148 34348 26200 34400
rect 27160 34391 27212 34400
rect 27160 34357 27169 34391
rect 27169 34357 27203 34391
rect 27203 34357 27212 34391
rect 27160 34348 27212 34357
rect 27436 34391 27488 34400
rect 27436 34357 27445 34391
rect 27445 34357 27479 34391
rect 27479 34357 27488 34391
rect 27436 34348 27488 34357
rect 27896 34348 27948 34400
rect 29000 34348 29052 34400
rect 31208 34348 31260 34400
rect 47216 34348 47268 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 17960 34187 18012 34196
rect 17960 34153 17969 34187
rect 17969 34153 18003 34187
rect 18003 34153 18012 34187
rect 17960 34144 18012 34153
rect 18144 34076 18196 34128
rect 16948 34008 17000 34060
rect 1308 33940 1360 33992
rect 15660 33983 15712 33992
rect 15660 33949 15669 33983
rect 15669 33949 15703 33983
rect 15703 33949 15712 33983
rect 15660 33940 15712 33949
rect 18144 33983 18196 33992
rect 18144 33949 18153 33983
rect 18153 33949 18187 33983
rect 18187 33949 18196 33983
rect 18144 33940 18196 33949
rect 18236 33940 18288 33992
rect 18604 33940 18656 33992
rect 16028 33872 16080 33924
rect 19340 33872 19392 33924
rect 1584 33804 1636 33856
rect 18604 33804 18656 33856
rect 20996 34144 21048 34196
rect 21732 34187 21784 34196
rect 21732 34153 21741 34187
rect 21741 34153 21775 34187
rect 21775 34153 21784 34187
rect 21732 34144 21784 34153
rect 22376 34144 22428 34196
rect 22836 34144 22888 34196
rect 27804 34144 27856 34196
rect 30288 34144 30340 34196
rect 31024 34187 31076 34196
rect 31024 34153 31033 34187
rect 31033 34153 31067 34187
rect 31067 34153 31076 34187
rect 31024 34144 31076 34153
rect 31300 34144 31352 34196
rect 28080 34076 28132 34128
rect 28356 34076 28408 34128
rect 46112 34076 46164 34128
rect 22284 34008 22336 34060
rect 21088 33872 21140 33924
rect 23480 33940 23532 33992
rect 27436 34008 27488 34060
rect 27896 34008 27948 34060
rect 47124 34051 47176 34060
rect 47124 34017 47133 34051
rect 47133 34017 47167 34051
rect 47167 34017 47176 34051
rect 47124 34008 47176 34017
rect 26792 33940 26844 33992
rect 27252 33940 27304 33992
rect 27620 33940 27672 33992
rect 29920 33983 29972 33992
rect 23296 33872 23348 33924
rect 24584 33872 24636 33924
rect 26516 33872 26568 33924
rect 27528 33872 27580 33924
rect 29920 33949 29929 33983
rect 29929 33949 29963 33983
rect 29963 33949 29972 33983
rect 29920 33940 29972 33949
rect 30104 33983 30156 33992
rect 30104 33949 30113 33983
rect 30113 33949 30147 33983
rect 30147 33949 30156 33983
rect 30104 33940 30156 33949
rect 31208 33983 31260 33992
rect 31208 33949 31217 33983
rect 31217 33949 31251 33983
rect 31251 33949 31260 33983
rect 31208 33940 31260 33949
rect 32128 33983 32180 33992
rect 32128 33949 32137 33983
rect 32137 33949 32171 33983
rect 32171 33949 32180 33983
rect 32128 33940 32180 33949
rect 47216 33915 47268 33924
rect 47216 33881 47225 33915
rect 47225 33881 47259 33915
rect 47259 33881 47268 33915
rect 47216 33872 47268 33881
rect 22468 33804 22520 33856
rect 23756 33847 23808 33856
rect 23756 33813 23765 33847
rect 23765 33813 23799 33847
rect 23799 33813 23808 33847
rect 23756 33804 23808 33813
rect 26148 33847 26200 33856
rect 26148 33813 26157 33847
rect 26157 33813 26191 33847
rect 26191 33813 26200 33847
rect 26148 33804 26200 33813
rect 27988 33804 28040 33856
rect 30840 33804 30892 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 16028 33643 16080 33652
rect 16028 33609 16037 33643
rect 16037 33609 16071 33643
rect 16071 33609 16080 33643
rect 16028 33600 16080 33609
rect 17132 33600 17184 33652
rect 18604 33643 18656 33652
rect 18604 33609 18613 33643
rect 18613 33609 18647 33643
rect 18647 33609 18656 33643
rect 18604 33600 18656 33609
rect 19248 33643 19300 33652
rect 19248 33609 19257 33643
rect 19257 33609 19291 33643
rect 19291 33609 19300 33643
rect 19248 33600 19300 33609
rect 22836 33600 22888 33652
rect 26148 33643 26200 33652
rect 26148 33609 26173 33643
rect 26173 33609 26200 33643
rect 26332 33643 26384 33652
rect 26148 33600 26200 33609
rect 26332 33609 26341 33643
rect 26341 33609 26375 33643
rect 26375 33609 26384 33643
rect 26332 33600 26384 33609
rect 28540 33643 28592 33652
rect 28540 33609 28549 33643
rect 28549 33609 28583 33643
rect 28583 33609 28592 33643
rect 28540 33600 28592 33609
rect 18144 33532 18196 33584
rect 18236 33532 18288 33584
rect 16672 33464 16724 33516
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 1676 33439 1728 33448
rect 1676 33405 1685 33439
rect 1685 33405 1719 33439
rect 1719 33405 1728 33439
rect 1676 33396 1728 33405
rect 17316 33507 17368 33516
rect 17316 33473 17325 33507
rect 17325 33473 17359 33507
rect 17359 33473 17368 33507
rect 17316 33464 17368 33473
rect 18512 33507 18564 33516
rect 17040 33396 17092 33448
rect 18512 33473 18521 33507
rect 18521 33473 18555 33507
rect 18555 33473 18564 33507
rect 18512 33464 18564 33473
rect 23756 33532 23808 33584
rect 18972 33464 19024 33516
rect 19340 33507 19392 33516
rect 19340 33473 19349 33507
rect 19349 33473 19383 33507
rect 19383 33473 19392 33507
rect 19340 33464 19392 33473
rect 22376 33464 22428 33516
rect 24952 33464 25004 33516
rect 26976 33575 27028 33584
rect 26976 33541 26985 33575
rect 26985 33541 27019 33575
rect 27019 33541 27028 33575
rect 26976 33532 27028 33541
rect 27436 33532 27488 33584
rect 32128 33600 32180 33652
rect 25596 33464 25648 33516
rect 25872 33464 25924 33516
rect 27160 33507 27212 33516
rect 27160 33473 27169 33507
rect 27169 33473 27203 33507
rect 27203 33473 27212 33507
rect 27160 33464 27212 33473
rect 28448 33507 28500 33516
rect 28448 33473 28457 33507
rect 28457 33473 28491 33507
rect 28491 33473 28500 33507
rect 28448 33464 28500 33473
rect 30656 33507 30708 33516
rect 23112 33439 23164 33448
rect 23112 33405 23121 33439
rect 23121 33405 23155 33439
rect 23155 33405 23164 33439
rect 23112 33396 23164 33405
rect 25044 33439 25096 33448
rect 25044 33405 25053 33439
rect 25053 33405 25087 33439
rect 25087 33405 25096 33439
rect 25044 33396 25096 33405
rect 26884 33396 26936 33448
rect 30656 33473 30665 33507
rect 30665 33473 30699 33507
rect 30699 33473 30708 33507
rect 30656 33464 30708 33473
rect 30840 33507 30892 33516
rect 30840 33473 30847 33507
rect 30847 33473 30892 33507
rect 30840 33464 30892 33473
rect 30104 33396 30156 33448
rect 32772 33532 32824 33584
rect 31208 33464 31260 33516
rect 31852 33464 31904 33516
rect 47768 33507 47820 33516
rect 47768 33473 47777 33507
rect 47777 33473 47811 33507
rect 47811 33473 47820 33507
rect 47768 33464 47820 33473
rect 18236 33328 18288 33380
rect 19432 33328 19484 33380
rect 18512 33260 18564 33312
rect 18696 33260 18748 33312
rect 22284 33303 22336 33312
rect 22284 33269 22293 33303
rect 22293 33269 22327 33303
rect 22327 33269 22336 33303
rect 22284 33260 22336 33269
rect 23756 33260 23808 33312
rect 25228 33303 25280 33312
rect 25228 33269 25237 33303
rect 25237 33269 25271 33303
rect 25271 33269 25280 33303
rect 25228 33260 25280 33269
rect 26148 33303 26200 33312
rect 26148 33269 26157 33303
rect 26157 33269 26191 33303
rect 26191 33269 26200 33303
rect 26148 33260 26200 33269
rect 26516 33260 26568 33312
rect 27528 33260 27580 33312
rect 29184 33303 29236 33312
rect 29184 33269 29193 33303
rect 29193 33269 29227 33303
rect 29227 33269 29236 33303
rect 29184 33260 29236 33269
rect 31300 33303 31352 33312
rect 31300 33269 31309 33303
rect 31309 33269 31343 33303
rect 31343 33269 31352 33303
rect 31300 33260 31352 33269
rect 32312 33260 32364 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 17500 33056 17552 33108
rect 22284 33056 22336 33108
rect 23020 33056 23072 33108
rect 25228 33056 25280 33108
rect 26332 33056 26384 33108
rect 26792 33099 26844 33108
rect 26792 33065 26801 33099
rect 26801 33065 26835 33099
rect 26835 33065 26844 33099
rect 26792 33056 26844 33065
rect 28172 33056 28224 33108
rect 30104 33056 30156 33108
rect 31852 33056 31904 33108
rect 32772 33099 32824 33108
rect 32772 33065 32781 33099
rect 32781 33065 32815 33099
rect 32815 33065 32824 33099
rect 32772 33056 32824 33065
rect 1492 32988 1544 33040
rect 16672 32988 16724 33040
rect 1584 32963 1636 32972
rect 1584 32929 1593 32963
rect 1593 32929 1627 32963
rect 1627 32929 1636 32963
rect 1584 32920 1636 32929
rect 12532 32920 12584 32972
rect 18420 32920 18472 32972
rect 20812 32920 20864 32972
rect 18236 32852 18288 32904
rect 18512 32895 18564 32904
rect 18512 32861 18521 32895
rect 18521 32861 18555 32895
rect 18555 32861 18564 32895
rect 18512 32852 18564 32861
rect 18604 32852 18656 32904
rect 18880 32852 18932 32904
rect 21548 32920 21600 32972
rect 23204 32988 23256 33040
rect 23480 32988 23532 33040
rect 24676 32988 24728 33040
rect 26424 32988 26476 33040
rect 22284 32920 22336 32972
rect 25044 32920 25096 32972
rect 3240 32827 3292 32836
rect 3240 32793 3249 32827
rect 3249 32793 3283 32827
rect 3283 32793 3292 32827
rect 3240 32784 3292 32793
rect 17960 32784 18012 32836
rect 19340 32827 19392 32836
rect 19340 32793 19349 32827
rect 19349 32793 19383 32827
rect 19383 32793 19392 32827
rect 19340 32784 19392 32793
rect 23940 32852 23992 32904
rect 25504 32895 25556 32904
rect 25504 32861 25513 32895
rect 25513 32861 25547 32895
rect 25547 32861 25556 32895
rect 25504 32852 25556 32861
rect 26516 32852 26568 32904
rect 28540 32920 28592 32972
rect 31300 32963 31352 32972
rect 31300 32929 31309 32963
rect 31309 32929 31343 32963
rect 31343 32929 31352 32963
rect 31300 32920 31352 32929
rect 28908 32852 28960 32904
rect 46296 32895 46348 32904
rect 46296 32861 46305 32895
rect 46305 32861 46339 32895
rect 46339 32861 46348 32895
rect 46296 32852 46348 32861
rect 16856 32759 16908 32768
rect 16856 32725 16865 32759
rect 16865 32725 16899 32759
rect 16899 32725 16908 32759
rect 16856 32716 16908 32725
rect 18052 32716 18104 32768
rect 18972 32716 19024 32768
rect 20996 32716 21048 32768
rect 22376 32716 22428 32768
rect 27160 32784 27212 32836
rect 27620 32784 27672 32836
rect 29184 32784 29236 32836
rect 32312 32784 32364 32836
rect 47676 32784 47728 32836
rect 48136 32827 48188 32836
rect 48136 32793 48145 32827
rect 48145 32793 48179 32827
rect 48179 32793 48188 32827
rect 48136 32784 48188 32793
rect 30104 32759 30156 32768
rect 30104 32725 30113 32759
rect 30113 32725 30147 32759
rect 30147 32725 30156 32759
rect 30104 32716 30156 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 18880 32512 18932 32564
rect 19064 32555 19116 32564
rect 19064 32521 19073 32555
rect 19073 32521 19107 32555
rect 19107 32521 19116 32555
rect 19064 32512 19116 32521
rect 1676 32444 1728 32496
rect 16856 32444 16908 32496
rect 18236 32444 18288 32496
rect 20996 32512 21048 32564
rect 19432 32444 19484 32496
rect 22284 32512 22336 32564
rect 25228 32512 25280 32564
rect 27620 32555 27672 32564
rect 27620 32521 27629 32555
rect 27629 32521 27663 32555
rect 27663 32521 27672 32555
rect 27620 32512 27672 32521
rect 30656 32512 30708 32564
rect 47676 32555 47728 32564
rect 47676 32521 47685 32555
rect 47685 32521 47719 32555
rect 47719 32521 47728 32555
rect 47676 32512 47728 32521
rect 15660 32376 15712 32428
rect 23112 32444 23164 32496
rect 25596 32444 25648 32496
rect 26148 32444 26200 32496
rect 27528 32444 27580 32496
rect 27896 32444 27948 32496
rect 2412 32308 2464 32360
rect 3240 32351 3292 32360
rect 3240 32317 3249 32351
rect 3249 32317 3283 32351
rect 3283 32317 3292 32351
rect 3240 32308 3292 32317
rect 16948 32351 17000 32360
rect 16948 32317 16957 32351
rect 16957 32317 16991 32351
rect 16991 32317 17000 32351
rect 16948 32308 17000 32317
rect 22836 32376 22888 32428
rect 23204 32419 23256 32428
rect 23204 32385 23213 32419
rect 23213 32385 23247 32419
rect 23247 32385 23256 32419
rect 23204 32376 23256 32385
rect 23848 32419 23900 32428
rect 23848 32385 23857 32419
rect 23857 32385 23891 32419
rect 23891 32385 23900 32419
rect 23848 32376 23900 32385
rect 24676 32419 24728 32428
rect 24676 32385 24685 32419
rect 24685 32385 24719 32419
rect 24719 32385 24728 32419
rect 24676 32376 24728 32385
rect 24860 32419 24912 32428
rect 24860 32385 24869 32419
rect 24869 32385 24903 32419
rect 24903 32385 24912 32419
rect 24860 32376 24912 32385
rect 24952 32376 25004 32428
rect 25504 32376 25556 32428
rect 26976 32419 27028 32428
rect 19524 32351 19576 32360
rect 19524 32317 19533 32351
rect 19533 32317 19567 32351
rect 19567 32317 19576 32351
rect 19524 32308 19576 32317
rect 22192 32351 22244 32360
rect 22192 32317 22201 32351
rect 22201 32317 22235 32351
rect 22235 32317 22244 32351
rect 22192 32308 22244 32317
rect 22560 32308 22612 32360
rect 23296 32308 23348 32360
rect 1400 32172 1452 32224
rect 18880 32215 18932 32224
rect 18880 32181 18889 32215
rect 18889 32181 18923 32215
rect 18923 32181 18932 32215
rect 18880 32172 18932 32181
rect 19248 32172 19300 32224
rect 22100 32283 22152 32292
rect 22100 32249 22109 32283
rect 22109 32249 22143 32283
rect 22143 32249 22152 32283
rect 22100 32240 22152 32249
rect 22376 32240 22428 32292
rect 25780 32283 25832 32292
rect 19708 32172 19760 32224
rect 20168 32215 20220 32224
rect 20168 32181 20177 32215
rect 20177 32181 20211 32215
rect 20211 32181 20220 32215
rect 20168 32172 20220 32181
rect 22744 32172 22796 32224
rect 23020 32172 23072 32224
rect 25780 32249 25789 32283
rect 25789 32249 25823 32283
rect 25823 32249 25832 32283
rect 25780 32240 25832 32249
rect 26976 32385 26985 32419
rect 26985 32385 27019 32419
rect 27019 32385 27028 32419
rect 26976 32376 27028 32385
rect 27160 32419 27212 32428
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27160 32376 27212 32385
rect 27804 32419 27856 32428
rect 27804 32385 27813 32419
rect 27813 32385 27847 32419
rect 27847 32385 27856 32419
rect 27988 32419 28040 32428
rect 27804 32376 27856 32385
rect 27988 32385 27997 32419
rect 27997 32385 28031 32419
rect 28031 32385 28040 32419
rect 27988 32376 28040 32385
rect 31576 32376 31628 32428
rect 46296 32376 46348 32428
rect 47492 32376 47544 32428
rect 26424 32351 26476 32360
rect 26424 32317 26433 32351
rect 26433 32317 26467 32351
rect 26467 32317 26476 32351
rect 26424 32308 26476 32317
rect 28264 32308 28316 32360
rect 30472 32351 30524 32360
rect 30472 32317 30481 32351
rect 30481 32317 30515 32351
rect 30515 32317 30524 32351
rect 30472 32308 30524 32317
rect 26792 32240 26844 32292
rect 27160 32240 27212 32292
rect 28172 32240 28224 32292
rect 29092 32240 29144 32292
rect 29460 32240 29512 32292
rect 28908 32172 28960 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 16948 31968 17000 32020
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 1860 31875 1912 31884
rect 1860 31841 1869 31875
rect 1869 31841 1903 31875
rect 1903 31841 1912 31875
rect 1860 31832 1912 31841
rect 17316 31875 17368 31884
rect 17316 31841 17325 31875
rect 17325 31841 17359 31875
rect 17359 31841 17368 31875
rect 17316 31832 17368 31841
rect 1584 31739 1636 31748
rect 1584 31705 1593 31739
rect 1593 31705 1627 31739
rect 1627 31705 1636 31739
rect 1584 31696 1636 31705
rect 17500 31764 17552 31816
rect 17960 31764 18012 31816
rect 18880 31832 18932 31884
rect 18972 31832 19024 31884
rect 20996 31968 21048 32020
rect 21180 31968 21232 32020
rect 20168 31832 20220 31884
rect 18696 31764 18748 31816
rect 19708 31807 19760 31816
rect 19708 31773 19717 31807
rect 19717 31773 19751 31807
rect 19751 31773 19760 31807
rect 19708 31764 19760 31773
rect 23204 31968 23256 32020
rect 26516 32011 26568 32020
rect 26516 31977 26525 32011
rect 26525 31977 26559 32011
rect 26559 31977 26568 32011
rect 26516 31968 26568 31977
rect 26792 31968 26844 32020
rect 30472 31968 30524 32020
rect 27896 31900 27948 31952
rect 28448 31943 28500 31952
rect 28448 31909 28457 31943
rect 28457 31909 28491 31943
rect 28491 31909 28500 31943
rect 28448 31900 28500 31909
rect 32312 31900 32364 31952
rect 22284 31875 22336 31884
rect 22284 31841 22293 31875
rect 22293 31841 22327 31875
rect 22327 31841 22336 31875
rect 22744 31875 22796 31884
rect 22284 31832 22336 31841
rect 22744 31841 22753 31875
rect 22753 31841 22787 31875
rect 22787 31841 22796 31875
rect 22744 31832 22796 31841
rect 30104 31832 30156 31884
rect 47308 31875 47360 31884
rect 23020 31764 23072 31816
rect 23204 31807 23256 31816
rect 23204 31773 23213 31807
rect 23213 31773 23247 31807
rect 23247 31773 23256 31807
rect 25228 31807 25280 31816
rect 23204 31764 23256 31773
rect 25228 31773 25237 31807
rect 25237 31773 25271 31807
rect 25271 31773 25280 31807
rect 25228 31764 25280 31773
rect 26516 31764 26568 31816
rect 30656 31807 30708 31816
rect 30656 31773 30665 31807
rect 30665 31773 30699 31807
rect 30699 31773 30708 31807
rect 30656 31764 30708 31773
rect 47308 31841 47317 31875
rect 47317 31841 47351 31875
rect 47351 31841 47360 31875
rect 47308 31832 47360 31841
rect 31116 31764 31168 31816
rect 46572 31764 46624 31816
rect 16856 31671 16908 31680
rect 16856 31637 16865 31671
rect 16865 31637 16899 31671
rect 16899 31637 16908 31671
rect 16856 31628 16908 31637
rect 17960 31628 18012 31680
rect 20720 31696 20772 31748
rect 23112 31739 23164 31748
rect 23112 31705 23121 31739
rect 23121 31705 23155 31739
rect 23155 31705 23164 31739
rect 23112 31696 23164 31705
rect 25596 31696 25648 31748
rect 26148 31696 26200 31748
rect 27528 31739 27580 31748
rect 27528 31705 27537 31739
rect 27537 31705 27571 31739
rect 27571 31705 27580 31739
rect 27528 31696 27580 31705
rect 20536 31628 20588 31680
rect 29552 31696 29604 31748
rect 30564 31696 30616 31748
rect 31208 31696 31260 31748
rect 29000 31628 29052 31680
rect 29460 31628 29512 31680
rect 30104 31628 30156 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1584 31424 1636 31476
rect 18604 31424 18656 31476
rect 18696 31424 18748 31476
rect 23204 31467 23256 31476
rect 16856 31356 16908 31408
rect 2320 31288 2372 31340
rect 18052 31288 18104 31340
rect 20444 31356 20496 31408
rect 23204 31433 23213 31467
rect 23213 31433 23247 31467
rect 23247 31433 23256 31467
rect 23204 31424 23256 31433
rect 23664 31424 23716 31476
rect 24308 31424 24360 31476
rect 24768 31424 24820 31476
rect 20996 31331 21048 31340
rect 20996 31297 21005 31331
rect 21005 31297 21039 31331
rect 21039 31297 21048 31331
rect 20996 31288 21048 31297
rect 22008 31288 22060 31340
rect 24860 31356 24912 31408
rect 24952 31356 25004 31408
rect 27804 31424 27856 31476
rect 29460 31424 29512 31476
rect 19340 31263 19392 31272
rect 19340 31229 19349 31263
rect 19349 31229 19383 31263
rect 19383 31229 19392 31263
rect 19340 31220 19392 31229
rect 23112 31288 23164 31340
rect 20812 31152 20864 31204
rect 21088 31195 21140 31204
rect 21088 31161 21097 31195
rect 21097 31161 21131 31195
rect 21131 31161 21140 31195
rect 21088 31152 21140 31161
rect 22468 31220 22520 31272
rect 23572 31288 23624 31340
rect 25412 31288 25464 31340
rect 24768 31220 24820 31272
rect 24952 31220 25004 31272
rect 25504 31152 25556 31204
rect 26148 31331 26200 31340
rect 26148 31297 26157 31331
rect 26157 31297 26191 31331
rect 26191 31297 26200 31331
rect 26148 31288 26200 31297
rect 27988 31288 28040 31340
rect 28172 31331 28224 31340
rect 28172 31297 28181 31331
rect 28181 31297 28215 31331
rect 28215 31297 28224 31331
rect 28172 31288 28224 31297
rect 28356 31288 28408 31340
rect 29552 31288 29604 31340
rect 45100 31424 45152 31476
rect 32128 31356 32180 31408
rect 30564 31331 30616 31340
rect 30104 31220 30156 31272
rect 30564 31297 30573 31331
rect 30573 31297 30607 31331
rect 30607 31297 30616 31331
rect 30564 31288 30616 31297
rect 32312 31331 32364 31340
rect 29920 31152 29972 31204
rect 32312 31297 32321 31331
rect 32321 31297 32355 31331
rect 32355 31297 32364 31331
rect 32312 31288 32364 31297
rect 32588 31331 32640 31340
rect 32588 31297 32597 31331
rect 32597 31297 32631 31331
rect 32631 31297 32640 31331
rect 32588 31288 32640 31297
rect 45560 31152 45612 31204
rect 46020 31152 46072 31204
rect 17960 31084 18012 31136
rect 22008 31084 22060 31136
rect 22652 31084 22704 31136
rect 28632 31084 28684 31136
rect 30012 31084 30064 31136
rect 32036 31084 32088 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 22376 30880 22428 30932
rect 24860 30880 24912 30932
rect 26976 30880 27028 30932
rect 29276 30880 29328 30932
rect 32588 30880 32640 30932
rect 28264 30812 28316 30864
rect 29828 30812 29880 30864
rect 8300 30744 8352 30796
rect 14648 30744 14700 30796
rect 14004 30676 14056 30728
rect 23388 30744 23440 30796
rect 14280 30651 14332 30660
rect 14280 30617 14289 30651
rect 14289 30617 14323 30651
rect 14323 30617 14332 30651
rect 14280 30608 14332 30617
rect 20720 30676 20772 30728
rect 21916 30676 21968 30728
rect 23848 30676 23900 30728
rect 24584 30676 24636 30728
rect 25412 30719 25464 30728
rect 25412 30685 25421 30719
rect 25421 30685 25455 30719
rect 25455 30685 25464 30719
rect 25412 30676 25464 30685
rect 26240 30719 26292 30728
rect 26240 30685 26249 30719
rect 26249 30685 26283 30719
rect 26283 30685 26292 30719
rect 26240 30676 26292 30685
rect 26792 30676 26844 30728
rect 29276 30744 29328 30796
rect 32036 30787 32088 30796
rect 17868 30651 17920 30660
rect 17868 30617 17877 30651
rect 17877 30617 17911 30651
rect 17911 30617 17920 30651
rect 17868 30608 17920 30617
rect 18144 30608 18196 30660
rect 20536 30608 20588 30660
rect 21272 30651 21324 30660
rect 21272 30617 21281 30651
rect 21281 30617 21315 30651
rect 21315 30617 21324 30651
rect 21272 30608 21324 30617
rect 22284 30608 22336 30660
rect 22652 30608 22704 30660
rect 27160 30608 27212 30660
rect 27528 30608 27580 30660
rect 29828 30676 29880 30728
rect 30012 30719 30064 30728
rect 30012 30685 30021 30719
rect 30021 30685 30055 30719
rect 30055 30685 30064 30719
rect 30012 30676 30064 30685
rect 30288 30719 30340 30728
rect 30288 30685 30297 30719
rect 30297 30685 30331 30719
rect 30331 30685 30340 30719
rect 30288 30676 30340 30685
rect 30656 30676 30708 30728
rect 30932 30719 30984 30728
rect 30932 30685 30941 30719
rect 30941 30685 30975 30719
rect 30975 30685 30984 30719
rect 30932 30676 30984 30685
rect 29184 30608 29236 30660
rect 30472 30608 30524 30660
rect 32036 30753 32045 30787
rect 32045 30753 32079 30787
rect 32079 30753 32088 30787
rect 32036 30744 32088 30753
rect 32496 30608 32548 30660
rect 18052 30540 18104 30592
rect 18236 30583 18288 30592
rect 18236 30549 18245 30583
rect 18245 30549 18279 30583
rect 18279 30549 18288 30583
rect 18236 30540 18288 30549
rect 21180 30540 21232 30592
rect 23020 30540 23072 30592
rect 23112 30540 23164 30592
rect 29000 30583 29052 30592
rect 29000 30549 29009 30583
rect 29009 30549 29043 30583
rect 29043 30549 29052 30583
rect 29000 30540 29052 30549
rect 30748 30540 30800 30592
rect 30932 30540 30984 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 17408 30336 17460 30388
rect 17868 30336 17920 30388
rect 30564 30336 30616 30388
rect 14280 30268 14332 30320
rect 16120 30311 16172 30320
rect 16120 30277 16129 30311
rect 16129 30277 16163 30311
rect 16163 30277 16172 30311
rect 16120 30268 16172 30277
rect 23296 30268 23348 30320
rect 26240 30268 26292 30320
rect 13636 30243 13688 30252
rect 13636 30209 13645 30243
rect 13645 30209 13679 30243
rect 13679 30209 13688 30243
rect 13636 30200 13688 30209
rect 18236 30243 18288 30252
rect 18236 30209 18245 30243
rect 18245 30209 18279 30243
rect 18279 30209 18288 30243
rect 18236 30200 18288 30209
rect 13912 30132 13964 30184
rect 14648 30132 14700 30184
rect 18512 30243 18564 30252
rect 18512 30209 18521 30243
rect 18521 30209 18555 30243
rect 18555 30209 18564 30243
rect 18512 30200 18564 30209
rect 21916 30200 21968 30252
rect 22468 30200 22520 30252
rect 22836 30243 22888 30252
rect 22836 30209 22845 30243
rect 22845 30209 22879 30243
rect 22879 30209 22888 30243
rect 22836 30200 22888 30209
rect 23020 30243 23072 30252
rect 23020 30209 23029 30243
rect 23029 30209 23063 30243
rect 23063 30209 23072 30243
rect 23020 30200 23072 30209
rect 23572 30200 23624 30252
rect 24584 30243 24636 30252
rect 24584 30209 24593 30243
rect 24593 30209 24627 30243
rect 24627 30209 24636 30243
rect 24584 30200 24636 30209
rect 25504 30243 25556 30252
rect 25504 30209 25513 30243
rect 25513 30209 25547 30243
rect 25547 30209 25556 30243
rect 25504 30200 25556 30209
rect 25780 30200 25832 30252
rect 27436 30200 27488 30252
rect 22376 30132 22428 30184
rect 23112 30175 23164 30184
rect 23112 30141 23121 30175
rect 23121 30141 23155 30175
rect 23155 30141 23164 30175
rect 23112 30132 23164 30141
rect 28448 30200 28500 30252
rect 29184 30243 29236 30252
rect 29184 30209 29193 30243
rect 29193 30209 29227 30243
rect 29227 30209 29236 30243
rect 29184 30200 29236 30209
rect 29736 30200 29788 30252
rect 29828 30200 29880 30252
rect 30288 30200 30340 30252
rect 30564 30200 30616 30252
rect 25688 30064 25740 30116
rect 18052 30039 18104 30048
rect 18052 30005 18061 30039
rect 18061 30005 18095 30039
rect 18095 30005 18104 30039
rect 18052 29996 18104 30005
rect 21272 29996 21324 30048
rect 22100 29996 22152 30048
rect 22652 29996 22704 30048
rect 25136 29996 25188 30048
rect 26976 30039 27028 30048
rect 26976 30005 26985 30039
rect 26985 30005 27019 30039
rect 27019 30005 27028 30039
rect 26976 29996 27028 30005
rect 27068 29996 27120 30048
rect 29644 30132 29696 30184
rect 32128 30268 32180 30320
rect 32496 30311 32548 30320
rect 32496 30277 32505 30311
rect 32505 30277 32539 30311
rect 32539 30277 32548 30311
rect 32496 30268 32548 30277
rect 32220 30200 32272 30252
rect 29276 29996 29328 30048
rect 30656 30064 30708 30116
rect 30380 30039 30432 30048
rect 30380 30005 30389 30039
rect 30389 30005 30423 30039
rect 30423 30005 30432 30039
rect 30380 29996 30432 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 14648 29835 14700 29844
rect 14648 29801 14657 29835
rect 14657 29801 14691 29835
rect 14691 29801 14700 29835
rect 14648 29792 14700 29801
rect 18512 29792 18564 29844
rect 22468 29835 22520 29844
rect 22468 29801 22477 29835
rect 22477 29801 22511 29835
rect 22511 29801 22520 29835
rect 22468 29792 22520 29801
rect 22192 29656 22244 29708
rect 13636 29588 13688 29640
rect 18144 29631 18196 29640
rect 18144 29597 18153 29631
rect 18153 29597 18187 29631
rect 18187 29597 18196 29631
rect 18144 29588 18196 29597
rect 20720 29588 20772 29640
rect 20904 29631 20956 29640
rect 20904 29597 20913 29631
rect 20913 29597 20947 29631
rect 20947 29597 20956 29631
rect 20904 29588 20956 29597
rect 22100 29631 22152 29640
rect 22100 29597 22109 29631
rect 22109 29597 22143 29631
rect 22143 29597 22152 29631
rect 22468 29631 22520 29640
rect 22100 29588 22152 29597
rect 22468 29597 22477 29631
rect 22477 29597 22511 29631
rect 22511 29597 22520 29631
rect 22468 29588 22520 29597
rect 22836 29656 22888 29708
rect 27252 29792 27304 29844
rect 28448 29792 28500 29844
rect 29920 29792 29972 29844
rect 30564 29792 30616 29844
rect 25688 29724 25740 29776
rect 28080 29724 28132 29776
rect 29644 29724 29696 29776
rect 30472 29699 30524 29708
rect 30472 29665 30481 29699
rect 30481 29665 30515 29699
rect 30515 29665 30524 29699
rect 30472 29656 30524 29665
rect 30748 29699 30800 29708
rect 30748 29665 30757 29699
rect 30757 29665 30791 29699
rect 30791 29665 30800 29699
rect 30748 29656 30800 29665
rect 23296 29631 23348 29640
rect 23296 29597 23305 29631
rect 23305 29597 23339 29631
rect 23339 29597 23348 29631
rect 23296 29588 23348 29597
rect 23572 29588 23624 29640
rect 18328 29520 18380 29572
rect 19984 29520 20036 29572
rect 21548 29452 21600 29504
rect 22192 29520 22244 29572
rect 23940 29588 23992 29640
rect 27068 29588 27120 29640
rect 25136 29520 25188 29572
rect 28172 29588 28224 29640
rect 28356 29588 28408 29640
rect 22928 29452 22980 29504
rect 23296 29452 23348 29504
rect 27712 29495 27764 29504
rect 27712 29461 27721 29495
rect 27721 29461 27755 29495
rect 27755 29461 27764 29495
rect 27712 29452 27764 29461
rect 27804 29452 27856 29504
rect 29000 29588 29052 29640
rect 47308 29631 47360 29640
rect 47308 29597 47317 29631
rect 47317 29597 47351 29631
rect 47351 29597 47360 29631
rect 47308 29588 47360 29597
rect 47400 29588 47452 29640
rect 29552 29563 29604 29572
rect 29552 29529 29561 29563
rect 29561 29529 29595 29563
rect 29595 29529 29604 29563
rect 29552 29520 29604 29529
rect 30380 29520 30432 29572
rect 32128 29520 32180 29572
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 7840 29180 7892 29232
rect 20536 29248 20588 29300
rect 20720 29248 20772 29300
rect 22100 29248 22152 29300
rect 24492 29248 24544 29300
rect 10876 29112 10928 29164
rect 13544 29112 13596 29164
rect 13912 29155 13964 29164
rect 13912 29121 13921 29155
rect 13921 29121 13955 29155
rect 13955 29121 13964 29155
rect 13912 29112 13964 29121
rect 20168 29153 20220 29164
rect 20168 29119 20177 29153
rect 20177 29119 20211 29153
rect 20211 29119 20220 29153
rect 20168 29112 20220 29119
rect 22192 29180 22244 29232
rect 22284 29155 22336 29164
rect 15844 29044 15896 29096
rect 16856 29087 16908 29096
rect 16856 29053 16865 29087
rect 16865 29053 16899 29087
rect 16899 29053 16908 29087
rect 16856 29044 16908 29053
rect 14096 28976 14148 29028
rect 16580 28976 16632 29028
rect 19984 29044 20036 29096
rect 22284 29121 22293 29155
rect 22293 29121 22327 29155
rect 22327 29121 22336 29155
rect 22284 29112 22336 29121
rect 22836 29180 22888 29232
rect 20536 29087 20588 29096
rect 20536 29053 20545 29087
rect 20545 29053 20579 29087
rect 20579 29053 20588 29087
rect 20536 29044 20588 29053
rect 20168 28976 20220 29028
rect 22008 28976 22060 29028
rect 22100 28976 22152 29028
rect 22468 28976 22520 29028
rect 13820 28951 13872 28960
rect 13820 28917 13829 28951
rect 13829 28917 13863 28951
rect 13863 28917 13872 28951
rect 13820 28908 13872 28917
rect 20904 28951 20956 28960
rect 20904 28917 20913 28951
rect 20913 28917 20947 28951
rect 20947 28917 20956 28951
rect 20904 28908 20956 28917
rect 22284 28951 22336 28960
rect 22284 28917 22293 28951
rect 22293 28917 22327 28951
rect 22327 28917 22336 28951
rect 22284 28908 22336 28917
rect 22376 28908 22428 28960
rect 23296 29155 23348 29164
rect 23296 29121 23305 29155
rect 23305 29121 23339 29155
rect 23339 29121 23348 29155
rect 23296 29112 23348 29121
rect 24952 29112 25004 29164
rect 27804 29112 27856 29164
rect 32128 29248 32180 29300
rect 28724 29180 28776 29232
rect 28080 29112 28132 29164
rect 28448 29112 28500 29164
rect 38292 29180 38344 29232
rect 27160 29087 27212 29096
rect 27160 29053 27169 29087
rect 27169 29053 27203 29087
rect 27203 29053 27212 29087
rect 27160 29044 27212 29053
rect 27712 29044 27764 29096
rect 25964 29019 26016 29028
rect 25964 28985 25973 29019
rect 25973 28985 26007 29019
rect 26007 28985 26016 29019
rect 25964 28976 26016 28985
rect 27896 28976 27948 29028
rect 29644 29044 29696 29096
rect 28264 28976 28316 29028
rect 29828 29112 29880 29164
rect 30380 29155 30432 29164
rect 30380 29121 30389 29155
rect 30389 29121 30423 29155
rect 30423 29121 30432 29155
rect 30380 29112 30432 29121
rect 32128 29155 32180 29164
rect 32128 29121 32137 29155
rect 32137 29121 32171 29155
rect 32171 29121 32180 29155
rect 32128 29112 32180 29121
rect 30840 28976 30892 29028
rect 27712 28908 27764 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 15844 28747 15896 28756
rect 15844 28713 15853 28747
rect 15853 28713 15887 28747
rect 15887 28713 15896 28747
rect 15844 28704 15896 28713
rect 18236 28704 18288 28756
rect 20720 28704 20772 28756
rect 21548 28747 21600 28756
rect 21548 28713 21557 28747
rect 21557 28713 21591 28747
rect 21591 28713 21600 28747
rect 21548 28704 21600 28713
rect 22008 28747 22060 28756
rect 22008 28713 22017 28747
rect 22017 28713 22051 28747
rect 22051 28713 22060 28747
rect 22008 28704 22060 28713
rect 22376 28704 22428 28756
rect 26792 28704 26844 28756
rect 20812 28636 20864 28688
rect 3700 28568 3752 28620
rect 13820 28568 13872 28620
rect 14096 28611 14148 28620
rect 14096 28577 14105 28611
rect 14105 28577 14139 28611
rect 14139 28577 14148 28611
rect 14096 28568 14148 28577
rect 17960 28568 18012 28620
rect 20904 28568 20956 28620
rect 22100 28568 22152 28620
rect 25964 28568 26016 28620
rect 28724 28704 28776 28756
rect 30380 28704 30432 28756
rect 28080 28636 28132 28688
rect 12072 28543 12124 28552
rect 12072 28509 12081 28543
rect 12081 28509 12115 28543
rect 12115 28509 12124 28543
rect 12072 28500 12124 28509
rect 13084 28500 13136 28552
rect 13176 28543 13228 28552
rect 13176 28509 13185 28543
rect 13185 28509 13219 28543
rect 13219 28509 13228 28543
rect 19248 28543 19300 28552
rect 13176 28500 13228 28509
rect 19248 28509 19257 28543
rect 19257 28509 19291 28543
rect 19291 28509 19300 28543
rect 19248 28500 19300 28509
rect 10048 28432 10100 28484
rect 9956 28364 10008 28416
rect 11796 28364 11848 28416
rect 14832 28432 14884 28484
rect 18880 28432 18932 28484
rect 19984 28432 20036 28484
rect 22192 28500 22244 28552
rect 22652 28543 22704 28552
rect 22652 28509 22661 28543
rect 22661 28509 22695 28543
rect 22695 28509 22704 28543
rect 22652 28500 22704 28509
rect 23296 28500 23348 28552
rect 27896 28543 27948 28552
rect 27896 28509 27905 28543
rect 27905 28509 27939 28543
rect 27939 28509 27948 28543
rect 27896 28500 27948 28509
rect 30840 28611 30892 28620
rect 30840 28577 30849 28611
rect 30849 28577 30883 28611
rect 30883 28577 30892 28611
rect 30840 28568 30892 28577
rect 47400 28568 47452 28620
rect 47676 28611 47728 28620
rect 47676 28577 47685 28611
rect 47685 28577 47719 28611
rect 47719 28577 47728 28611
rect 47676 28568 47728 28577
rect 28172 28543 28224 28552
rect 28172 28509 28181 28543
rect 28181 28509 28215 28543
rect 28215 28509 28224 28543
rect 28172 28500 28224 28509
rect 28356 28500 28408 28552
rect 28540 28500 28592 28552
rect 18052 28364 18104 28416
rect 27436 28432 27488 28484
rect 29736 28432 29788 28484
rect 30472 28432 30524 28484
rect 32220 28432 32272 28484
rect 46572 28432 46624 28484
rect 22468 28364 22520 28416
rect 28448 28364 28500 28416
rect 28724 28364 28776 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 10048 28203 10100 28212
rect 10048 28169 10057 28203
rect 10057 28169 10091 28203
rect 10091 28169 10100 28203
rect 10048 28160 10100 28169
rect 14832 28160 14884 28212
rect 16856 28160 16908 28212
rect 18880 28160 18932 28212
rect 19984 28203 20036 28212
rect 19984 28169 19993 28203
rect 19993 28169 20027 28203
rect 20027 28169 20036 28203
rect 19984 28160 20036 28169
rect 22100 28160 22152 28212
rect 23204 28160 23256 28212
rect 28172 28160 28224 28212
rect 32220 28203 32272 28212
rect 32220 28169 32229 28203
rect 32229 28169 32263 28203
rect 32263 28169 32272 28203
rect 32220 28160 32272 28169
rect 11796 28135 11848 28144
rect 11796 28101 11805 28135
rect 11805 28101 11839 28135
rect 11839 28101 11848 28135
rect 11796 28092 11848 28101
rect 20720 28092 20772 28144
rect 23756 28092 23808 28144
rect 25596 28092 25648 28144
rect 25872 28135 25924 28144
rect 25872 28101 25881 28135
rect 25881 28101 25915 28135
rect 25915 28101 25924 28135
rect 25872 28092 25924 28101
rect 25964 28092 26016 28144
rect 28724 28135 28776 28144
rect 10876 28067 10928 28076
rect 10876 28033 10885 28067
rect 10885 28033 10919 28067
rect 10919 28033 10928 28067
rect 10876 28024 10928 28033
rect 14096 28024 14148 28076
rect 18604 28024 18656 28076
rect 20812 28067 20864 28076
rect 20812 28033 20821 28067
rect 20821 28033 20855 28067
rect 20855 28033 20864 28067
rect 20812 28024 20864 28033
rect 22652 28067 22704 28076
rect 22652 28033 22661 28067
rect 22661 28033 22695 28067
rect 22695 28033 22704 28067
rect 22652 28024 22704 28033
rect 16028 27956 16080 28008
rect 16672 27999 16724 28008
rect 16672 27965 16681 27999
rect 16681 27965 16715 27999
rect 16715 27965 16724 27999
rect 16672 27956 16724 27965
rect 16856 27999 16908 28008
rect 16856 27965 16865 27999
rect 16865 27965 16899 27999
rect 16899 27965 16908 27999
rect 16856 27956 16908 27965
rect 21088 27956 21140 28008
rect 26792 28024 26844 28076
rect 28724 28101 28733 28135
rect 28733 28101 28767 28135
rect 28767 28101 28776 28135
rect 28724 28092 28776 28101
rect 30840 28092 30892 28144
rect 27344 28024 27396 28076
rect 28448 28067 28500 28076
rect 28448 28033 28457 28067
rect 28457 28033 28491 28067
rect 28491 28033 28500 28067
rect 28448 28024 28500 28033
rect 30656 28024 30708 28076
rect 32128 28067 32180 28076
rect 32128 28033 32137 28067
rect 32137 28033 32171 28067
rect 32171 28033 32180 28067
rect 32128 28024 32180 28033
rect 27896 27956 27948 28008
rect 28816 27956 28868 28008
rect 47676 28160 47728 28212
rect 47124 28024 47176 28076
rect 47584 28067 47636 28076
rect 47584 28033 47593 28067
rect 47593 28033 47627 28067
rect 47627 28033 47636 28067
rect 47584 28024 47636 28033
rect 3976 27820 4028 27872
rect 13268 27863 13320 27872
rect 13268 27829 13277 27863
rect 13277 27829 13311 27863
rect 13311 27829 13320 27863
rect 13268 27820 13320 27829
rect 22192 27820 22244 27872
rect 24492 27888 24544 27940
rect 24216 27863 24268 27872
rect 24216 27829 24225 27863
rect 24225 27829 24259 27863
rect 24259 27829 24268 27863
rect 24216 27820 24268 27829
rect 27068 27863 27120 27872
rect 27068 27829 27077 27863
rect 27077 27829 27111 27863
rect 27111 27829 27120 27863
rect 27068 27820 27120 27829
rect 29460 27820 29512 27872
rect 47032 27863 47084 27872
rect 47032 27829 47041 27863
rect 47041 27829 47075 27863
rect 47075 27829 47084 27863
rect 47032 27820 47084 27829
rect 47676 27863 47728 27872
rect 47676 27829 47685 27863
rect 47685 27829 47719 27863
rect 47719 27829 47728 27863
rect 47676 27820 47728 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 12072 27616 12124 27668
rect 9772 27480 9824 27532
rect 10876 27480 10928 27532
rect 10600 27412 10652 27464
rect 13176 27616 13228 27668
rect 13084 27548 13136 27600
rect 14004 27548 14056 27600
rect 11980 27344 12032 27396
rect 13268 27412 13320 27464
rect 15844 27616 15896 27668
rect 16856 27616 16908 27668
rect 22376 27616 22428 27668
rect 27068 27616 27120 27668
rect 28356 27616 28408 27668
rect 30012 27616 30064 27668
rect 43536 27616 43588 27668
rect 46204 27616 46256 27668
rect 25596 27548 25648 27600
rect 22192 27523 22244 27532
rect 22192 27489 22201 27523
rect 22201 27489 22235 27523
rect 22235 27489 22244 27523
rect 22192 27480 22244 27489
rect 27252 27480 27304 27532
rect 30656 27548 30708 27600
rect 30840 27591 30892 27600
rect 30840 27557 30849 27591
rect 30849 27557 30883 27591
rect 30883 27557 30892 27591
rect 30840 27548 30892 27557
rect 15752 27455 15804 27464
rect 15752 27421 15761 27455
rect 15761 27421 15795 27455
rect 15795 27421 15804 27455
rect 15752 27412 15804 27421
rect 17776 27412 17828 27464
rect 13544 27344 13596 27396
rect 13912 27344 13964 27396
rect 9128 27276 9180 27328
rect 10876 27276 10928 27328
rect 14648 27319 14700 27328
rect 14648 27285 14657 27319
rect 14657 27285 14691 27319
rect 14691 27285 14700 27319
rect 14648 27276 14700 27285
rect 15936 27319 15988 27328
rect 15936 27285 15945 27319
rect 15945 27285 15979 27319
rect 15979 27285 15988 27319
rect 15936 27276 15988 27285
rect 22744 27344 22796 27396
rect 22284 27276 22336 27328
rect 22652 27276 22704 27328
rect 23756 27412 23808 27464
rect 24216 27412 24268 27464
rect 26792 27412 26844 27464
rect 26976 27455 27028 27464
rect 26976 27421 26985 27455
rect 26985 27421 27019 27455
rect 27019 27421 27028 27455
rect 26976 27412 27028 27421
rect 28908 27412 28960 27464
rect 29460 27412 29512 27464
rect 27988 27344 28040 27396
rect 28172 27344 28224 27396
rect 23388 27276 23440 27328
rect 25688 27276 25740 27328
rect 25872 27276 25924 27328
rect 30012 27412 30064 27464
rect 47032 27480 47084 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 40408 27344 40460 27396
rect 47676 27344 47728 27396
rect 29828 27276 29880 27328
rect 30104 27276 30156 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 1768 27072 1820 27124
rect 10416 27004 10468 27056
rect 9128 26979 9180 26988
rect 9128 26945 9137 26979
rect 9137 26945 9171 26979
rect 9171 26945 9180 26979
rect 9128 26936 9180 26945
rect 12808 26979 12860 26988
rect 12808 26945 12817 26979
rect 12817 26945 12851 26979
rect 12851 26945 12860 26979
rect 12808 26936 12860 26945
rect 12992 26979 13044 26988
rect 12992 26945 13001 26979
rect 13001 26945 13035 26979
rect 13035 26945 13044 26979
rect 12992 26936 13044 26945
rect 13544 26979 13596 26988
rect 13544 26945 13553 26979
rect 13553 26945 13587 26979
rect 13587 26945 13596 26979
rect 13544 26936 13596 26945
rect 14648 27004 14700 27056
rect 15200 27004 15252 27056
rect 16120 27004 16172 27056
rect 13820 26936 13872 26988
rect 15936 26936 15988 26988
rect 16580 26936 16632 26988
rect 9404 26911 9456 26920
rect 9404 26877 9413 26911
rect 9413 26877 9447 26911
rect 9447 26877 9456 26911
rect 9404 26868 9456 26877
rect 14004 26868 14056 26920
rect 10600 26800 10652 26852
rect 15660 26800 15712 26852
rect 16764 26800 16816 26852
rect 10876 26775 10928 26784
rect 10876 26741 10885 26775
rect 10885 26741 10919 26775
rect 10919 26741 10928 26775
rect 10876 26732 10928 26741
rect 12072 26732 12124 26784
rect 16396 26732 16448 26784
rect 22376 27004 22428 27056
rect 20720 26936 20772 26988
rect 22284 26979 22336 26988
rect 22284 26945 22293 26979
rect 22293 26945 22327 26979
rect 22327 26945 22336 26979
rect 22284 26936 22336 26945
rect 22744 26936 22796 26988
rect 24216 27072 24268 27124
rect 24676 27072 24728 27124
rect 24860 27004 24912 27056
rect 26792 27004 26844 27056
rect 25780 26936 25832 26988
rect 26884 26936 26936 26988
rect 26976 26979 27028 26988
rect 26976 26945 26985 26979
rect 26985 26945 27019 26979
rect 27019 26945 27028 26979
rect 28356 27004 28408 27056
rect 29828 27072 29880 27124
rect 30104 27047 30156 27056
rect 26976 26936 27028 26945
rect 30104 27013 30113 27047
rect 30113 27013 30147 27047
rect 30147 27013 30156 27047
rect 30104 27004 30156 27013
rect 29736 26936 29788 26988
rect 32128 26979 32180 26988
rect 32128 26945 32137 26979
rect 32137 26945 32171 26979
rect 32171 26945 32180 26979
rect 32128 26936 32180 26945
rect 22100 26800 22152 26852
rect 22192 26800 22244 26852
rect 25320 26868 25372 26920
rect 28264 26868 28316 26920
rect 27252 26800 27304 26852
rect 27436 26843 27488 26852
rect 27436 26809 27445 26843
rect 27445 26809 27479 26843
rect 27479 26809 27488 26843
rect 27436 26800 27488 26809
rect 20812 26732 20864 26784
rect 23756 26732 23808 26784
rect 25688 26732 25740 26784
rect 26884 26732 26936 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 9404 26528 9456 26580
rect 14004 26528 14056 26580
rect 16580 26528 16632 26580
rect 22284 26528 22336 26580
rect 24952 26571 25004 26580
rect 24952 26537 24961 26571
rect 24961 26537 24995 26571
rect 24995 26537 25004 26571
rect 24952 26528 25004 26537
rect 26608 26528 26660 26580
rect 10600 26392 10652 26444
rect 12072 26435 12124 26444
rect 12072 26401 12081 26435
rect 12081 26401 12115 26435
rect 12115 26401 12124 26435
rect 12072 26392 12124 26401
rect 10876 26324 10928 26376
rect 14096 26367 14148 26376
rect 14096 26333 14105 26367
rect 14105 26333 14139 26367
rect 14139 26333 14148 26367
rect 14096 26324 14148 26333
rect 16028 26392 16080 26444
rect 16396 26435 16448 26444
rect 16396 26401 16405 26435
rect 16405 26401 16439 26435
rect 16439 26401 16448 26435
rect 16396 26392 16448 26401
rect 15660 26367 15712 26376
rect 15660 26333 15669 26367
rect 15669 26333 15703 26367
rect 15703 26333 15712 26367
rect 15660 26324 15712 26333
rect 17500 26324 17552 26376
rect 18328 26367 18380 26376
rect 18328 26333 18337 26367
rect 18337 26333 18371 26367
rect 18371 26333 18380 26367
rect 18328 26324 18380 26333
rect 23664 26460 23716 26512
rect 24676 26460 24728 26512
rect 23388 26392 23440 26444
rect 21640 26324 21692 26376
rect 22100 26324 22152 26376
rect 27160 26460 27212 26512
rect 27436 26460 27488 26512
rect 25320 26392 25372 26444
rect 26976 26392 27028 26444
rect 47124 26460 47176 26512
rect 25688 26367 25740 26376
rect 25688 26333 25697 26367
rect 25697 26333 25731 26367
rect 25731 26333 25740 26367
rect 25688 26324 25740 26333
rect 25780 26324 25832 26376
rect 27252 26367 27304 26376
rect 27252 26333 27261 26367
rect 27261 26333 27295 26367
rect 27295 26333 27304 26367
rect 27252 26324 27304 26333
rect 27436 26324 27488 26376
rect 28264 26367 28316 26376
rect 28264 26333 28273 26367
rect 28273 26333 28307 26367
rect 28307 26333 28316 26367
rect 28264 26324 28316 26333
rect 46940 26392 46992 26444
rect 47768 26435 47820 26444
rect 47768 26401 47777 26435
rect 47777 26401 47811 26435
rect 47811 26401 47820 26435
rect 47768 26392 47820 26401
rect 32128 26324 32180 26376
rect 12716 26188 12768 26240
rect 16672 26256 16724 26308
rect 21272 26256 21324 26308
rect 21824 26256 21876 26308
rect 25872 26299 25924 26308
rect 25872 26265 25881 26299
rect 25881 26265 25915 26299
rect 25915 26265 25924 26299
rect 25872 26256 25924 26265
rect 26884 26256 26936 26308
rect 32312 26256 32364 26308
rect 43444 26256 43496 26308
rect 46296 26256 46348 26308
rect 48044 26256 48096 26308
rect 16764 26188 16816 26240
rect 17868 26231 17920 26240
rect 17868 26197 17877 26231
rect 17877 26197 17911 26231
rect 17911 26197 17920 26231
rect 17868 26188 17920 26197
rect 18512 26188 18564 26240
rect 19432 26188 19484 26240
rect 20996 26231 21048 26240
rect 20996 26197 21005 26231
rect 21005 26197 21039 26231
rect 21039 26197 21048 26231
rect 26240 26231 26292 26240
rect 20996 26188 21048 26197
rect 26240 26197 26249 26231
rect 26249 26197 26283 26231
rect 26283 26197 26292 26231
rect 26240 26188 26292 26197
rect 27988 26188 28040 26240
rect 32036 26188 32088 26240
rect 45652 26188 45704 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 10416 25984 10468 26036
rect 12716 26027 12768 26036
rect 12716 25993 12725 26027
rect 12725 25993 12759 26027
rect 12759 25993 12768 26027
rect 12716 25984 12768 25993
rect 15752 26027 15804 26036
rect 15752 25993 15761 26027
rect 15761 25993 15795 26027
rect 15795 25993 15804 26027
rect 15752 25984 15804 25993
rect 16764 25984 16816 26036
rect 20720 25984 20772 26036
rect 16028 25916 16080 25968
rect 16580 25916 16632 25968
rect 17868 25916 17920 25968
rect 18512 25959 18564 25968
rect 18512 25925 18521 25959
rect 18521 25925 18555 25959
rect 18555 25925 18564 25959
rect 18512 25916 18564 25925
rect 46204 25984 46256 26036
rect 26976 25959 27028 25968
rect 26976 25925 26985 25959
rect 26985 25925 27019 25959
rect 27019 25925 27028 25959
rect 26976 25916 27028 25925
rect 27252 25916 27304 25968
rect 28356 25916 28408 25968
rect 10232 25891 10284 25900
rect 10232 25857 10241 25891
rect 10241 25857 10275 25891
rect 10275 25857 10284 25891
rect 10232 25848 10284 25857
rect 13452 25848 13504 25900
rect 15568 25891 15620 25900
rect 15568 25857 15577 25891
rect 15577 25857 15611 25891
rect 15611 25857 15620 25891
rect 15568 25848 15620 25857
rect 15108 25780 15160 25832
rect 15568 25712 15620 25764
rect 21732 25848 21784 25900
rect 21824 25891 21876 25900
rect 21824 25857 21833 25891
rect 21833 25857 21867 25891
rect 21867 25857 21876 25891
rect 21824 25848 21876 25857
rect 18328 25823 18380 25832
rect 18328 25789 18337 25823
rect 18337 25789 18371 25823
rect 18371 25789 18380 25823
rect 18328 25780 18380 25789
rect 21272 25823 21324 25832
rect 21272 25789 21281 25823
rect 21281 25789 21315 25823
rect 21315 25789 21324 25823
rect 27988 25891 28040 25900
rect 21272 25780 21324 25789
rect 22100 25712 22152 25764
rect 22468 25780 22520 25832
rect 27988 25857 27997 25891
rect 27997 25857 28031 25891
rect 28031 25857 28040 25891
rect 27988 25848 28040 25857
rect 28172 25891 28224 25900
rect 28172 25857 28181 25891
rect 28181 25857 28215 25891
rect 28215 25857 28224 25891
rect 28172 25848 28224 25857
rect 32128 25916 32180 25968
rect 32312 25959 32364 25968
rect 32312 25925 32321 25959
rect 32321 25925 32355 25959
rect 32355 25925 32364 25959
rect 32312 25916 32364 25925
rect 43444 25916 43496 25968
rect 45652 25848 45704 25900
rect 28264 25823 28316 25832
rect 28264 25789 28273 25823
rect 28273 25789 28307 25823
rect 28307 25789 28316 25823
rect 28264 25780 28316 25789
rect 28356 25823 28408 25832
rect 28356 25789 28365 25823
rect 28365 25789 28399 25823
rect 28399 25789 28408 25823
rect 31300 25823 31352 25832
rect 28356 25780 28408 25789
rect 31300 25789 31309 25823
rect 31309 25789 31343 25823
rect 31343 25789 31352 25823
rect 31300 25780 31352 25789
rect 23388 25712 23440 25764
rect 24032 25712 24084 25764
rect 21180 25687 21232 25696
rect 21180 25653 21189 25687
rect 21189 25653 21223 25687
rect 21223 25653 21232 25687
rect 21180 25644 21232 25653
rect 22284 25687 22336 25696
rect 22284 25653 22293 25687
rect 22293 25653 22327 25687
rect 22327 25653 22336 25687
rect 22284 25644 22336 25653
rect 22744 25644 22796 25696
rect 27528 25644 27580 25696
rect 31300 25644 31352 25696
rect 47400 25780 47452 25832
rect 46296 25712 46348 25764
rect 46480 25644 46532 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 16672 25483 16724 25492
rect 16672 25449 16681 25483
rect 16681 25449 16715 25483
rect 16715 25449 16724 25483
rect 16672 25440 16724 25449
rect 17500 25440 17552 25492
rect 20996 25440 21048 25492
rect 22284 25440 22336 25492
rect 28264 25440 28316 25492
rect 21732 25415 21784 25424
rect 21732 25381 21741 25415
rect 21741 25381 21775 25415
rect 21775 25381 21784 25415
rect 21732 25372 21784 25381
rect 22100 25372 22152 25424
rect 22560 25372 22612 25424
rect 12808 25304 12860 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 9864 25279 9916 25288
rect 9864 25245 9873 25279
rect 9873 25245 9907 25279
rect 9907 25245 9916 25279
rect 9864 25236 9916 25245
rect 12348 25236 12400 25288
rect 15476 25236 15528 25288
rect 18328 25304 18380 25356
rect 15844 25236 15896 25288
rect 16580 25279 16632 25288
rect 16580 25245 16589 25279
rect 16589 25245 16623 25279
rect 16623 25245 16632 25279
rect 16580 25236 16632 25245
rect 17500 25279 17552 25288
rect 17500 25245 17509 25279
rect 17509 25245 17543 25279
rect 17543 25245 17552 25279
rect 17500 25236 17552 25245
rect 18604 25236 18656 25288
rect 19248 25279 19300 25288
rect 19248 25245 19257 25279
rect 19257 25245 19291 25279
rect 19291 25245 19300 25279
rect 19248 25236 19300 25245
rect 21272 25236 21324 25288
rect 21732 25236 21784 25288
rect 22744 25279 22796 25288
rect 1676 25211 1728 25220
rect 1676 25177 1685 25211
rect 1685 25177 1719 25211
rect 1719 25177 1728 25211
rect 1676 25168 1728 25177
rect 10140 25211 10192 25220
rect 10140 25177 10149 25211
rect 10149 25177 10183 25211
rect 10183 25177 10192 25211
rect 10140 25168 10192 25177
rect 11428 25168 11480 25220
rect 19432 25168 19484 25220
rect 22744 25245 22753 25279
rect 22753 25245 22787 25279
rect 22787 25245 22796 25279
rect 22744 25236 22796 25245
rect 26240 25304 26292 25356
rect 46480 25347 46532 25356
rect 46480 25313 46489 25347
rect 46489 25313 46523 25347
rect 46523 25313 46532 25347
rect 46480 25304 46532 25313
rect 48136 25347 48188 25356
rect 48136 25313 48145 25347
rect 48145 25313 48179 25347
rect 48179 25313 48188 25347
rect 48136 25304 48188 25313
rect 25596 25279 25648 25288
rect 25596 25245 25605 25279
rect 25605 25245 25639 25279
rect 25639 25245 25648 25279
rect 25596 25236 25648 25245
rect 27252 25279 27304 25288
rect 27252 25245 27261 25279
rect 27261 25245 27295 25279
rect 27295 25245 27304 25279
rect 27252 25236 27304 25245
rect 32128 25279 32180 25288
rect 32128 25245 32137 25279
rect 32137 25245 32171 25279
rect 32171 25245 32180 25279
rect 32128 25236 32180 25245
rect 45652 25279 45704 25288
rect 45652 25245 45661 25279
rect 45661 25245 45695 25279
rect 45695 25245 45704 25279
rect 45652 25236 45704 25245
rect 11060 25100 11112 25152
rect 12992 25143 13044 25152
rect 12992 25109 13001 25143
rect 13001 25109 13035 25143
rect 13035 25109 13044 25143
rect 12992 25100 13044 25109
rect 15568 25143 15620 25152
rect 15568 25109 15577 25143
rect 15577 25109 15611 25143
rect 15611 25109 15620 25143
rect 15568 25100 15620 25109
rect 15660 25100 15712 25152
rect 22836 25168 22888 25220
rect 24860 25168 24912 25220
rect 27528 25211 27580 25220
rect 27528 25177 27537 25211
rect 27537 25177 27571 25211
rect 27571 25177 27580 25211
rect 27528 25168 27580 25177
rect 28080 25168 28132 25220
rect 31208 25168 31260 25220
rect 32772 25211 32824 25220
rect 21180 25100 21232 25152
rect 25412 25100 25464 25152
rect 32772 25177 32781 25211
rect 32781 25177 32815 25211
rect 32815 25177 32824 25211
rect 32772 25168 32824 25177
rect 43076 25168 43128 25220
rect 46572 25168 46624 25220
rect 41236 25100 41288 25152
rect 45560 25100 45612 25152
rect 46020 25100 46072 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9864 24939 9916 24948
rect 9864 24905 9873 24939
rect 9873 24905 9907 24939
rect 9907 24905 9916 24939
rect 9864 24896 9916 24905
rect 10140 24896 10192 24948
rect 11704 24896 11756 24948
rect 12348 24896 12400 24948
rect 15292 24896 15344 24948
rect 16764 24896 16816 24948
rect 18328 24896 18380 24948
rect 21272 24939 21324 24948
rect 21272 24905 21281 24939
rect 21281 24905 21315 24939
rect 21315 24905 21324 24939
rect 21272 24896 21324 24905
rect 22836 24896 22888 24948
rect 25320 24896 25372 24948
rect 12992 24828 13044 24880
rect 13544 24828 13596 24880
rect 15476 24871 15528 24880
rect 15476 24837 15485 24871
rect 15485 24837 15519 24871
rect 15519 24837 15528 24871
rect 15476 24828 15528 24837
rect 15660 24871 15712 24880
rect 15660 24837 15669 24871
rect 15669 24837 15703 24871
rect 15703 24837 15712 24871
rect 15660 24828 15712 24837
rect 9772 24803 9824 24812
rect 9772 24769 9781 24803
rect 9781 24769 9815 24803
rect 9815 24769 9824 24803
rect 9772 24760 9824 24769
rect 10416 24803 10468 24812
rect 10416 24769 10425 24803
rect 10425 24769 10459 24803
rect 10459 24769 10468 24803
rect 10416 24760 10468 24769
rect 10600 24803 10652 24812
rect 10600 24769 10609 24803
rect 10609 24769 10643 24803
rect 10643 24769 10652 24803
rect 10600 24760 10652 24769
rect 10232 24692 10284 24744
rect 15200 24760 15252 24812
rect 17684 24828 17736 24880
rect 20444 24828 20496 24880
rect 24492 24828 24544 24880
rect 22560 24803 22612 24812
rect 22560 24769 22569 24803
rect 22569 24769 22603 24803
rect 22603 24769 22612 24803
rect 22560 24760 22612 24769
rect 23112 24760 23164 24812
rect 25044 24760 25096 24812
rect 28080 24803 28132 24812
rect 28080 24769 28089 24803
rect 28089 24769 28123 24803
rect 28123 24769 28132 24803
rect 32128 24803 32180 24812
rect 28080 24760 28132 24769
rect 32128 24769 32137 24803
rect 32137 24769 32171 24803
rect 32171 24769 32180 24803
rect 32128 24760 32180 24769
rect 11428 24692 11480 24744
rect 14096 24692 14148 24744
rect 16672 24735 16724 24744
rect 16672 24701 16681 24735
rect 16681 24701 16715 24735
rect 16715 24701 16724 24735
rect 16672 24692 16724 24701
rect 16948 24735 17000 24744
rect 16948 24701 16957 24735
rect 16957 24701 16991 24735
rect 16991 24701 17000 24735
rect 16948 24692 17000 24701
rect 19248 24692 19300 24744
rect 23756 24735 23808 24744
rect 3516 24624 3568 24676
rect 12532 24624 12584 24676
rect 12440 24556 12492 24608
rect 18420 24556 18472 24608
rect 23756 24701 23765 24735
rect 23765 24701 23799 24735
rect 23799 24701 23808 24735
rect 23756 24692 23808 24701
rect 25228 24692 25280 24744
rect 29276 24692 29328 24744
rect 29644 24692 29696 24744
rect 29828 24735 29880 24744
rect 29828 24701 29837 24735
rect 29837 24701 29871 24735
rect 29871 24701 29880 24735
rect 29828 24692 29880 24701
rect 32036 24692 32088 24744
rect 45376 24735 45428 24744
rect 45008 24624 45060 24676
rect 26424 24556 26476 24608
rect 45376 24701 45385 24735
rect 45385 24701 45419 24735
rect 45419 24701 45428 24735
rect 45376 24692 45428 24701
rect 46848 24735 46900 24744
rect 46848 24701 46857 24735
rect 46857 24701 46891 24735
rect 46891 24701 46900 24735
rect 46848 24692 46900 24701
rect 45284 24624 45336 24676
rect 46204 24624 46256 24676
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 10416 24352 10468 24404
rect 3884 24284 3936 24336
rect 13544 24284 13596 24336
rect 14096 24327 14148 24336
rect 14096 24293 14105 24327
rect 14105 24293 14139 24327
rect 14139 24293 14148 24327
rect 14096 24284 14148 24293
rect 15292 24327 15344 24336
rect 15292 24293 15301 24327
rect 15301 24293 15335 24327
rect 15335 24293 15344 24327
rect 15292 24284 15344 24293
rect 1952 24216 2004 24268
rect 12440 24216 12492 24268
rect 12532 24259 12584 24268
rect 12532 24225 12541 24259
rect 12541 24225 12575 24259
rect 12575 24225 12584 24259
rect 12532 24216 12584 24225
rect 9588 24148 9640 24200
rect 10140 24148 10192 24200
rect 11060 24191 11112 24200
rect 11060 24157 11069 24191
rect 11069 24157 11103 24191
rect 11103 24157 11112 24191
rect 11060 24148 11112 24157
rect 12716 24148 12768 24200
rect 14004 24148 14056 24200
rect 15568 24216 15620 24268
rect 16948 24284 17000 24336
rect 17684 24284 17736 24336
rect 20444 24327 20496 24336
rect 20444 24293 20453 24327
rect 20453 24293 20487 24327
rect 20487 24293 20496 24327
rect 20444 24284 20496 24293
rect 24492 24352 24544 24404
rect 26884 24327 26936 24336
rect 26884 24293 26893 24327
rect 26893 24293 26927 24327
rect 26927 24293 26936 24327
rect 26884 24284 26936 24293
rect 29644 24327 29696 24336
rect 29644 24293 29653 24327
rect 29653 24293 29687 24327
rect 29687 24293 29696 24327
rect 29644 24284 29696 24293
rect 33140 24284 33192 24336
rect 16580 24216 16632 24268
rect 18604 24216 18656 24268
rect 10232 24080 10284 24132
rect 11244 24123 11296 24132
rect 11244 24089 11253 24123
rect 11253 24089 11287 24123
rect 11287 24089 11296 24123
rect 11244 24080 11296 24089
rect 13452 24080 13504 24132
rect 15752 24148 15804 24200
rect 16856 24148 16908 24200
rect 17500 24148 17552 24200
rect 19432 24191 19484 24200
rect 15200 24080 15252 24132
rect 15936 24080 15988 24132
rect 19432 24157 19441 24191
rect 19441 24157 19475 24191
rect 19475 24157 19484 24191
rect 19432 24148 19484 24157
rect 27252 24216 27304 24268
rect 46020 24259 46072 24268
rect 46020 24225 46029 24259
rect 46029 24225 46063 24259
rect 46063 24225 46072 24259
rect 46020 24216 46072 24225
rect 47308 24259 47360 24268
rect 47308 24225 47317 24259
rect 47317 24225 47351 24259
rect 47351 24225 47360 24259
rect 47308 24216 47360 24225
rect 25044 24148 25096 24200
rect 29184 24148 29236 24200
rect 30196 24148 30248 24200
rect 8208 24012 8260 24064
rect 9772 24055 9824 24064
rect 9772 24021 9781 24055
rect 9781 24021 9815 24055
rect 9815 24021 9824 24055
rect 9772 24012 9824 24021
rect 10508 24055 10560 24064
rect 10508 24021 10517 24055
rect 10517 24021 10551 24055
rect 10551 24021 10560 24055
rect 10508 24012 10560 24021
rect 15476 24055 15528 24064
rect 15476 24021 15485 24055
rect 15485 24021 15519 24055
rect 15519 24021 15528 24055
rect 15476 24012 15528 24021
rect 15844 24055 15896 24064
rect 15844 24021 15853 24055
rect 15853 24021 15887 24055
rect 15887 24021 15896 24055
rect 15844 24012 15896 24021
rect 16764 24012 16816 24064
rect 20076 24080 20128 24132
rect 25412 24123 25464 24132
rect 25412 24089 25421 24123
rect 25421 24089 25455 24123
rect 25455 24089 25464 24123
rect 25412 24080 25464 24089
rect 26424 24080 26476 24132
rect 47032 24080 47084 24132
rect 21916 24012 21968 24064
rect 45560 24012 45612 24064
rect 45836 24012 45888 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1952 23851 2004 23860
rect 1952 23817 1961 23851
rect 1961 23817 1995 23851
rect 1995 23817 2004 23851
rect 1952 23808 2004 23817
rect 3424 23808 3476 23860
rect 9772 23740 9824 23792
rect 29828 23808 29880 23860
rect 45376 23808 45428 23860
rect 11060 23740 11112 23792
rect 14556 23740 14608 23792
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 8208 23715 8260 23724
rect 8208 23681 8217 23715
rect 8217 23681 8251 23715
rect 8251 23681 8260 23715
rect 8208 23672 8260 23681
rect 12992 23672 13044 23724
rect 15292 23715 15344 23724
rect 15292 23681 15301 23715
rect 15301 23681 15335 23715
rect 15335 23681 15344 23715
rect 15292 23672 15344 23681
rect 16120 23672 16172 23724
rect 16580 23672 16632 23724
rect 17592 23672 17644 23724
rect 21916 23740 21968 23792
rect 8484 23647 8536 23656
rect 8484 23613 8493 23647
rect 8493 23613 8527 23647
rect 8527 23613 8536 23647
rect 8484 23604 8536 23613
rect 9956 23647 10008 23656
rect 9956 23613 9965 23647
rect 9965 23613 9999 23647
rect 9999 23613 10008 23647
rect 9956 23604 10008 23613
rect 15476 23604 15528 23656
rect 17684 23604 17736 23656
rect 17868 23604 17920 23656
rect 9680 23536 9732 23588
rect 10600 23536 10652 23588
rect 15108 23536 15160 23588
rect 16672 23579 16724 23588
rect 16672 23545 16681 23579
rect 16681 23545 16715 23579
rect 16715 23545 16724 23579
rect 16672 23536 16724 23545
rect 18604 23536 18656 23588
rect 23480 23672 23532 23724
rect 37280 23740 37332 23792
rect 23388 23604 23440 23656
rect 28724 23672 28776 23724
rect 45836 23715 45888 23724
rect 23848 23604 23900 23656
rect 26424 23604 26476 23656
rect 31116 23647 31168 23656
rect 31116 23613 31125 23647
rect 31125 23613 31159 23647
rect 31159 23613 31168 23647
rect 31116 23604 31168 23613
rect 45836 23681 45845 23715
rect 45845 23681 45879 23715
rect 45879 23681 45888 23715
rect 45836 23672 45888 23681
rect 46664 23672 46716 23724
rect 47492 23672 47544 23724
rect 20076 23536 20128 23588
rect 23204 23536 23256 23588
rect 28908 23536 28960 23588
rect 31760 23536 31812 23588
rect 33048 23604 33100 23656
rect 33140 23647 33192 23656
rect 33140 23613 33149 23647
rect 33149 23613 33183 23647
rect 33183 23613 33192 23647
rect 33140 23604 33192 23613
rect 44732 23647 44784 23656
rect 32496 23536 32548 23588
rect 44732 23613 44741 23647
rect 44741 23613 44775 23647
rect 44775 23613 44784 23647
rect 44732 23604 44784 23613
rect 46388 23604 46440 23656
rect 46848 23536 46900 23588
rect 10508 23468 10560 23520
rect 13452 23511 13504 23520
rect 13452 23477 13461 23511
rect 13461 23477 13495 23511
rect 13495 23477 13504 23511
rect 13452 23468 13504 23477
rect 19340 23468 19392 23520
rect 20168 23511 20220 23520
rect 20168 23477 20177 23511
rect 20177 23477 20211 23511
rect 20211 23477 20220 23511
rect 20168 23468 20220 23477
rect 23020 23511 23072 23520
rect 23020 23477 23029 23511
rect 23029 23477 23063 23511
rect 23063 23477 23072 23511
rect 23020 23468 23072 23477
rect 23572 23511 23624 23520
rect 23572 23477 23581 23511
rect 23581 23477 23615 23511
rect 23615 23477 23624 23511
rect 23572 23468 23624 23477
rect 32036 23468 32088 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 8484 23264 8536 23316
rect 9956 23264 10008 23316
rect 10232 23264 10284 23316
rect 10508 23307 10560 23316
rect 10508 23273 10517 23307
rect 10517 23273 10551 23307
rect 10551 23273 10560 23307
rect 10508 23264 10560 23273
rect 11244 23264 11296 23316
rect 14556 23307 14608 23316
rect 14556 23273 14565 23307
rect 14565 23273 14599 23307
rect 14599 23273 14608 23307
rect 14556 23264 14608 23273
rect 18236 23307 18288 23316
rect 18236 23273 18245 23307
rect 18245 23273 18279 23307
rect 18279 23273 18288 23307
rect 18236 23264 18288 23273
rect 20260 23264 20312 23316
rect 47584 23264 47636 23316
rect 10692 23196 10744 23248
rect 10600 23128 10652 23180
rect 15844 23196 15896 23248
rect 15752 23171 15804 23180
rect 15752 23137 15761 23171
rect 15761 23137 15795 23171
rect 15795 23137 15804 23171
rect 15752 23128 15804 23137
rect 19432 23128 19484 23180
rect 23572 23128 23624 23180
rect 24124 23128 24176 23180
rect 30288 23128 30340 23180
rect 31760 23171 31812 23180
rect 31760 23137 31769 23171
rect 31769 23137 31803 23171
rect 31803 23137 31812 23171
rect 31760 23128 31812 23137
rect 32036 23171 32088 23180
rect 32036 23137 32045 23171
rect 32045 23137 32079 23171
rect 32079 23137 32088 23171
rect 32036 23128 32088 23137
rect 32496 23128 32548 23180
rect 9772 23060 9824 23112
rect 11060 23060 11112 23112
rect 15660 23060 15712 23112
rect 16120 23060 16172 23112
rect 9956 22992 10008 23044
rect 12992 22992 13044 23044
rect 15292 22992 15344 23044
rect 10048 22924 10100 22976
rect 10324 22967 10376 22976
rect 10324 22933 10349 22967
rect 10349 22933 10376 22967
rect 10324 22924 10376 22933
rect 15200 22924 15252 22976
rect 15384 22924 15436 22976
rect 19432 23035 19484 23044
rect 19432 23001 19441 23035
rect 19441 23001 19475 23035
rect 19475 23001 19484 23035
rect 19432 22992 19484 23001
rect 21180 22992 21232 23044
rect 28540 23060 28592 23112
rect 31484 23060 31536 23112
rect 22284 22992 22336 23044
rect 23020 22992 23072 23044
rect 29828 23035 29880 23044
rect 19984 22924 20036 22976
rect 29828 23001 29837 23035
rect 29837 23001 29871 23035
rect 29871 23001 29880 23035
rect 29828 22992 29880 23001
rect 32496 22992 32548 23044
rect 41512 23128 41564 23180
rect 41788 23171 41840 23180
rect 41788 23137 41797 23171
rect 41797 23137 41831 23171
rect 41831 23137 41840 23171
rect 41788 23128 41840 23137
rect 46296 23171 46348 23180
rect 46296 23137 46305 23171
rect 46305 23137 46339 23171
rect 46339 23137 46348 23171
rect 46296 23128 46348 23137
rect 46756 23171 46808 23180
rect 46756 23137 46765 23171
rect 46765 23137 46799 23171
rect 46799 23137 46808 23171
rect 46756 23128 46808 23137
rect 33416 23060 33468 23112
rect 39764 23060 39816 23112
rect 39948 23103 40000 23112
rect 39948 23069 39957 23103
rect 39957 23069 39991 23103
rect 39991 23069 40000 23103
rect 39948 23060 40000 23069
rect 46020 23060 46072 23112
rect 40132 23035 40184 23044
rect 40132 23001 40141 23035
rect 40141 23001 40175 23035
rect 40175 23001 40184 23035
rect 40132 22992 40184 23001
rect 47676 22992 47728 23044
rect 33876 22924 33928 22976
rect 42800 22924 42852 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9772 22720 9824 22772
rect 12716 22763 12768 22772
rect 12716 22729 12725 22763
rect 12725 22729 12759 22763
rect 12759 22729 12768 22763
rect 12716 22720 12768 22729
rect 13360 22720 13412 22772
rect 9680 22652 9732 22704
rect 10232 22695 10284 22704
rect 10232 22661 10241 22695
rect 10241 22661 10275 22695
rect 10275 22661 10284 22695
rect 10232 22652 10284 22661
rect 10692 22652 10744 22704
rect 15752 22720 15804 22772
rect 22928 22720 22980 22772
rect 24124 22763 24176 22772
rect 15384 22652 15436 22704
rect 24124 22729 24133 22763
rect 24133 22729 24167 22763
rect 24167 22729 24176 22763
rect 28540 22763 28592 22772
rect 24124 22720 24176 22729
rect 9496 22448 9548 22500
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 9864 22380 9916 22432
rect 10324 22380 10376 22432
rect 11888 22380 11940 22432
rect 13452 22516 13504 22568
rect 16672 22584 16724 22636
rect 18236 22584 18288 22636
rect 18788 22627 18840 22636
rect 14096 22559 14148 22568
rect 14096 22525 14105 22559
rect 14105 22525 14139 22559
rect 14139 22525 14148 22559
rect 14096 22516 14148 22525
rect 17684 22516 17736 22568
rect 18788 22593 18797 22627
rect 18797 22593 18831 22627
rect 18831 22593 18840 22627
rect 18788 22584 18840 22593
rect 19984 22584 20036 22636
rect 20260 22584 20312 22636
rect 20904 22627 20956 22636
rect 20904 22593 20913 22627
rect 20913 22593 20947 22627
rect 20947 22593 20956 22627
rect 20904 22584 20956 22593
rect 28540 22729 28549 22763
rect 28549 22729 28583 22763
rect 28583 22729 28592 22763
rect 28540 22720 28592 22729
rect 30748 22763 30800 22772
rect 30748 22729 30757 22763
rect 30757 22729 30791 22763
rect 30791 22729 30800 22763
rect 30748 22720 30800 22729
rect 31116 22720 31168 22772
rect 31484 22763 31536 22772
rect 31484 22729 31493 22763
rect 31493 22729 31527 22763
rect 31527 22729 31536 22763
rect 31484 22720 31536 22729
rect 32496 22720 32548 22772
rect 33048 22763 33100 22772
rect 33048 22729 33057 22763
rect 33057 22729 33091 22763
rect 33091 22729 33100 22763
rect 33048 22720 33100 22729
rect 40132 22763 40184 22772
rect 40132 22729 40141 22763
rect 40141 22729 40175 22763
rect 40175 22729 40184 22763
rect 40132 22720 40184 22729
rect 45836 22720 45888 22772
rect 47676 22763 47728 22772
rect 47676 22729 47685 22763
rect 47685 22729 47719 22763
rect 47719 22729 47728 22763
rect 47676 22720 47728 22729
rect 22376 22584 22428 22636
rect 23848 22627 23900 22636
rect 20812 22559 20864 22568
rect 20812 22525 20821 22559
rect 20821 22525 20855 22559
rect 20855 22525 20864 22559
rect 23848 22593 23857 22627
rect 23857 22593 23891 22627
rect 23891 22593 23900 22627
rect 23848 22584 23900 22593
rect 23940 22584 23992 22636
rect 39948 22652 40000 22704
rect 41512 22695 41564 22704
rect 41512 22661 41521 22695
rect 41521 22661 41555 22695
rect 41555 22661 41564 22695
rect 41512 22652 41564 22661
rect 20812 22516 20864 22525
rect 15936 22448 15988 22500
rect 17868 22491 17920 22500
rect 17868 22457 17877 22491
rect 17877 22457 17911 22491
rect 17911 22457 17920 22491
rect 17868 22448 17920 22457
rect 16120 22380 16172 22432
rect 16856 22423 16908 22432
rect 16856 22389 16865 22423
rect 16865 22389 16899 22423
rect 16899 22389 16908 22423
rect 16856 22380 16908 22389
rect 20812 22380 20864 22432
rect 21088 22380 21140 22432
rect 21272 22423 21324 22432
rect 21272 22389 21281 22423
rect 21281 22389 21315 22423
rect 21315 22389 21324 22423
rect 21272 22380 21324 22389
rect 21824 22380 21876 22432
rect 22836 22448 22888 22500
rect 23480 22516 23532 22568
rect 23388 22491 23440 22500
rect 23388 22457 23397 22491
rect 23397 22457 23431 22491
rect 23431 22457 23440 22491
rect 23388 22448 23440 22457
rect 23020 22380 23072 22432
rect 25964 22584 26016 22636
rect 28540 22627 28592 22636
rect 28540 22593 28549 22627
rect 28549 22593 28583 22627
rect 28583 22593 28592 22627
rect 28540 22584 28592 22593
rect 28724 22584 28776 22636
rect 29276 22627 29328 22636
rect 29276 22593 29285 22627
rect 29285 22593 29319 22627
rect 29319 22593 29328 22627
rect 29276 22584 29328 22593
rect 30288 22584 30340 22636
rect 30564 22627 30616 22636
rect 30564 22593 30573 22627
rect 30573 22593 30607 22627
rect 30607 22593 30616 22627
rect 30564 22584 30616 22593
rect 31392 22627 31444 22636
rect 29828 22516 29880 22568
rect 31392 22593 31401 22627
rect 31401 22593 31435 22627
rect 31435 22593 31444 22627
rect 31392 22584 31444 22593
rect 33416 22584 33468 22636
rect 39764 22584 39816 22636
rect 31116 22516 31168 22568
rect 33876 22559 33928 22568
rect 33876 22525 33885 22559
rect 33885 22525 33919 22559
rect 33919 22525 33928 22559
rect 33876 22516 33928 22525
rect 30288 22448 30340 22500
rect 41604 22516 41656 22568
rect 45836 22584 45888 22636
rect 47584 22627 47636 22636
rect 47584 22593 47593 22627
rect 47593 22593 47627 22627
rect 47627 22593 47636 22627
rect 47584 22584 47636 22593
rect 43536 22448 43588 22500
rect 25228 22423 25280 22432
rect 25228 22389 25237 22423
rect 25237 22389 25271 22423
rect 25271 22389 25280 22423
rect 25228 22380 25280 22389
rect 25688 22423 25740 22432
rect 25688 22389 25697 22423
rect 25697 22389 25731 22423
rect 25731 22389 25740 22423
rect 25688 22380 25740 22389
rect 26240 22380 26292 22432
rect 31208 22380 31260 22432
rect 41604 22423 41656 22432
rect 41604 22389 41613 22423
rect 41613 22389 41647 22423
rect 41647 22389 41656 22423
rect 41604 22380 41656 22389
rect 46204 22516 46256 22568
rect 46756 22559 46808 22568
rect 46756 22525 46765 22559
rect 46765 22525 46799 22559
rect 46799 22525 46808 22559
rect 46756 22516 46808 22525
rect 45928 22491 45980 22500
rect 45928 22457 45937 22491
rect 45937 22457 45971 22491
rect 45971 22457 45980 22491
rect 45928 22448 45980 22457
rect 47492 22380 47544 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 9496 22219 9548 22228
rect 9496 22185 9505 22219
rect 9505 22185 9539 22219
rect 9539 22185 9548 22219
rect 9496 22176 9548 22185
rect 14096 22219 14148 22228
rect 14096 22185 14105 22219
rect 14105 22185 14139 22219
rect 14139 22185 14148 22219
rect 14096 22176 14148 22185
rect 21272 22176 21324 22228
rect 22284 22219 22336 22228
rect 22284 22185 22293 22219
rect 22293 22185 22327 22219
rect 22327 22185 22336 22219
rect 22284 22176 22336 22185
rect 22376 22176 22428 22228
rect 26240 22176 26292 22228
rect 26424 22219 26476 22228
rect 26424 22185 26433 22219
rect 26433 22185 26467 22219
rect 26467 22185 26476 22219
rect 26424 22176 26476 22185
rect 9772 22040 9824 22092
rect 10048 22040 10100 22092
rect 11888 22083 11940 22092
rect 11888 22049 11897 22083
rect 11897 22049 11931 22083
rect 11931 22049 11940 22083
rect 11888 22040 11940 22049
rect 13360 22040 13412 22092
rect 10692 21972 10744 22024
rect 11704 22015 11756 22024
rect 11704 21981 11713 22015
rect 11713 21981 11747 22015
rect 11747 21981 11756 22015
rect 11704 21972 11756 21981
rect 13544 21972 13596 22024
rect 15384 22040 15436 22092
rect 17960 22083 18012 22092
rect 9772 21904 9824 21956
rect 10140 21904 10192 21956
rect 11428 21904 11480 21956
rect 13452 21904 13504 21956
rect 17960 22049 17969 22083
rect 17969 22049 18003 22083
rect 18003 22049 18012 22083
rect 17960 22040 18012 22049
rect 23848 22108 23900 22160
rect 19248 22015 19300 22024
rect 8208 21879 8260 21888
rect 8208 21845 8217 21879
rect 8217 21845 8251 21879
rect 8251 21845 8260 21879
rect 8208 21836 8260 21845
rect 9956 21836 10008 21888
rect 10600 21836 10652 21888
rect 19248 21981 19257 22015
rect 19257 21981 19291 22015
rect 19291 21981 19300 22015
rect 19248 21972 19300 21981
rect 16948 21947 17000 21956
rect 16948 21913 16957 21947
rect 16957 21913 16991 21947
rect 16991 21913 17000 21947
rect 16948 21904 17000 21913
rect 20904 22040 20956 22092
rect 21732 22083 21784 22092
rect 21732 22049 21741 22083
rect 21741 22049 21775 22083
rect 21775 22049 21784 22083
rect 21732 22040 21784 22049
rect 19984 22015 20036 22024
rect 19984 21981 19993 22015
rect 19993 21981 20027 22015
rect 20027 21981 20036 22015
rect 19984 21972 20036 21981
rect 22560 21972 22612 22024
rect 25688 22040 25740 22092
rect 27712 22040 27764 22092
rect 30288 22176 30340 22228
rect 41512 22176 41564 22228
rect 45836 22219 45888 22228
rect 45836 22185 45845 22219
rect 45845 22185 45879 22219
rect 45879 22185 45888 22219
rect 45836 22176 45888 22185
rect 31116 22108 31168 22160
rect 23664 21972 23716 22024
rect 26884 22015 26936 22024
rect 26884 21981 26893 22015
rect 26893 21981 26927 22015
rect 26927 21981 26936 22015
rect 26884 21972 26936 21981
rect 28264 21972 28316 22024
rect 20996 21904 21048 21956
rect 20076 21836 20128 21888
rect 21824 21836 21876 21888
rect 23296 21836 23348 21888
rect 24676 21904 24728 21956
rect 24860 21904 24912 21956
rect 26240 21904 26292 21956
rect 23940 21836 23992 21888
rect 27344 21836 27396 21888
rect 44732 22040 44784 22092
rect 47768 22083 47820 22092
rect 47768 22049 47777 22083
rect 47777 22049 47811 22083
rect 47811 22049 47820 22083
rect 47768 22040 47820 22049
rect 30748 21972 30800 22024
rect 41236 22015 41288 22024
rect 41236 21981 41245 22015
rect 41245 21981 41279 22015
rect 41279 21981 41288 22015
rect 41236 21972 41288 21981
rect 45560 21972 45612 22024
rect 45836 21972 45888 22024
rect 46296 22015 46348 22024
rect 46296 21981 46305 22015
rect 46305 21981 46339 22015
rect 46339 21981 46348 22015
rect 46296 21972 46348 21981
rect 30564 21904 30616 21956
rect 31944 21904 31996 21956
rect 29920 21836 29972 21888
rect 30380 21836 30432 21888
rect 31116 21836 31168 21888
rect 43996 21879 44048 21888
rect 43996 21845 44005 21879
rect 44005 21845 44039 21879
rect 44039 21845 44048 21879
rect 43996 21836 44048 21845
rect 45928 21836 45980 21888
rect 46296 21836 46348 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4620 21632 4672 21684
rect 10048 21632 10100 21684
rect 16948 21632 17000 21684
rect 20444 21632 20496 21684
rect 22560 21632 22612 21684
rect 23296 21632 23348 21684
rect 24860 21675 24912 21684
rect 8208 21564 8260 21616
rect 10140 21564 10192 21616
rect 13452 21496 13504 21548
rect 16672 21564 16724 21616
rect 16856 21607 16908 21616
rect 16856 21573 16865 21607
rect 16865 21573 16899 21607
rect 16899 21573 16908 21607
rect 16856 21564 16908 21573
rect 19248 21564 19300 21616
rect 22284 21564 22336 21616
rect 22468 21564 22520 21616
rect 15936 21539 15988 21548
rect 15936 21505 15945 21539
rect 15945 21505 15979 21539
rect 15979 21505 15988 21539
rect 15936 21496 15988 21505
rect 19892 21496 19944 21548
rect 22192 21539 22244 21548
rect 22192 21505 22201 21539
rect 22201 21505 22235 21539
rect 22235 21505 22244 21539
rect 22192 21496 22244 21505
rect 22560 21496 22612 21548
rect 9128 21471 9180 21480
rect 9128 21437 9137 21471
rect 9137 21437 9171 21471
rect 9171 21437 9180 21471
rect 9128 21428 9180 21437
rect 9772 21428 9824 21480
rect 18328 21471 18380 21480
rect 18328 21437 18337 21471
rect 18337 21437 18371 21471
rect 18371 21437 18380 21471
rect 18328 21428 18380 21437
rect 23388 21428 23440 21480
rect 22100 21360 22152 21412
rect 24860 21641 24869 21675
rect 24869 21641 24903 21675
rect 24903 21641 24912 21675
rect 24860 21632 24912 21641
rect 26240 21675 26292 21684
rect 26240 21641 26249 21675
rect 26249 21641 26283 21675
rect 26283 21641 26292 21675
rect 26240 21632 26292 21641
rect 28264 21675 28316 21684
rect 28264 21641 28273 21675
rect 28273 21641 28307 21675
rect 28307 21641 28316 21675
rect 28264 21632 28316 21641
rect 28356 21632 28408 21684
rect 24676 21496 24728 21548
rect 25228 21496 25280 21548
rect 25964 21360 26016 21412
rect 29920 21564 29972 21616
rect 27344 21539 27396 21548
rect 27344 21505 27353 21539
rect 27353 21505 27387 21539
rect 27387 21505 27396 21539
rect 27344 21496 27396 21505
rect 30380 21564 30432 21616
rect 30288 21539 30340 21548
rect 27712 21471 27764 21480
rect 27712 21437 27721 21471
rect 27721 21437 27755 21471
rect 27755 21437 27764 21471
rect 27712 21428 27764 21437
rect 30288 21505 30297 21539
rect 30297 21505 30331 21539
rect 30331 21505 30340 21539
rect 30288 21496 30340 21505
rect 31392 21496 31444 21548
rect 42064 21632 42116 21684
rect 46204 21675 46256 21684
rect 43996 21607 44048 21616
rect 43996 21573 44005 21607
rect 44005 21573 44039 21607
rect 44039 21573 44048 21607
rect 43996 21564 44048 21573
rect 46204 21641 46213 21675
rect 46213 21641 46247 21675
rect 46247 21641 46256 21675
rect 46204 21632 46256 21641
rect 47952 21607 48004 21616
rect 47952 21573 47961 21607
rect 47961 21573 47995 21607
rect 47995 21573 48004 21607
rect 47952 21564 48004 21573
rect 45836 21496 45888 21548
rect 45928 21496 45980 21548
rect 46296 21539 46348 21548
rect 46296 21505 46305 21539
rect 46305 21505 46339 21539
rect 46339 21505 46348 21539
rect 46296 21496 46348 21505
rect 46664 21496 46716 21548
rect 45376 21471 45428 21480
rect 45376 21437 45385 21471
rect 45385 21437 45419 21471
rect 45419 21437 45428 21471
rect 45376 21428 45428 21437
rect 10416 21292 10468 21344
rect 13360 21335 13412 21344
rect 13360 21301 13369 21335
rect 13369 21301 13403 21335
rect 13403 21301 13412 21335
rect 13360 21292 13412 21301
rect 15844 21292 15896 21344
rect 21088 21292 21140 21344
rect 22376 21292 22428 21344
rect 23664 21292 23716 21344
rect 30472 21292 30524 21344
rect 31208 21292 31260 21344
rect 46480 21292 46532 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 9128 21088 9180 21140
rect 10140 21088 10192 21140
rect 15936 21088 15988 21140
rect 19984 21088 20036 21140
rect 20996 21088 21048 21140
rect 20 20816 72 20868
rect 15844 20995 15896 21004
rect 15844 20961 15853 20995
rect 15853 20961 15887 20995
rect 15887 20961 15896 20995
rect 15844 20952 15896 20961
rect 26884 21020 26936 21072
rect 20076 20952 20128 21004
rect 9404 20927 9456 20936
rect 9404 20893 9413 20927
rect 9413 20893 9447 20927
rect 9447 20893 9456 20927
rect 9404 20884 9456 20893
rect 10416 20884 10468 20936
rect 11060 20884 11112 20936
rect 11520 20927 11572 20936
rect 11520 20893 11529 20927
rect 11529 20893 11563 20927
rect 11563 20893 11572 20927
rect 11520 20884 11572 20893
rect 13360 20884 13412 20936
rect 15660 20927 15712 20936
rect 15660 20893 15669 20927
rect 15669 20893 15703 20927
rect 15703 20893 15712 20927
rect 15660 20884 15712 20893
rect 17868 20884 17920 20936
rect 19432 20884 19484 20936
rect 20444 20927 20496 20936
rect 20444 20893 20453 20927
rect 20453 20893 20487 20927
rect 20487 20893 20496 20927
rect 20444 20884 20496 20893
rect 22100 20995 22152 21004
rect 22100 20961 22109 20995
rect 22109 20961 22143 20995
rect 22143 20961 22152 20995
rect 22376 20995 22428 21004
rect 22100 20952 22152 20961
rect 22376 20961 22385 20995
rect 22385 20961 22419 20995
rect 22419 20961 22428 20995
rect 22376 20952 22428 20961
rect 30472 20995 30524 21004
rect 30472 20961 30481 20995
rect 30481 20961 30515 20995
rect 30515 20961 30524 20995
rect 30472 20952 30524 20961
rect 46388 21020 46440 21072
rect 46480 20995 46532 21004
rect 46480 20961 46489 20995
rect 46489 20961 46523 20995
rect 46523 20961 46532 20995
rect 46480 20952 46532 20961
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 21824 20884 21876 20936
rect 25964 20927 26016 20936
rect 25964 20893 25973 20927
rect 25973 20893 26007 20927
rect 26007 20893 26016 20927
rect 25964 20884 26016 20893
rect 30196 20927 30248 20936
rect 30196 20893 30205 20927
rect 30205 20893 30239 20927
rect 30239 20893 30248 20927
rect 30196 20884 30248 20893
rect 33416 20884 33468 20936
rect 45560 20884 45612 20936
rect 23664 20816 23716 20868
rect 31208 20816 31260 20868
rect 47768 20816 47820 20868
rect 14648 20791 14700 20800
rect 14648 20757 14657 20791
rect 14657 20757 14691 20791
rect 14691 20757 14700 20791
rect 14648 20748 14700 20757
rect 19340 20791 19392 20800
rect 19340 20757 19349 20791
rect 19349 20757 19383 20791
rect 19383 20757 19392 20791
rect 19340 20748 19392 20757
rect 22192 20748 22244 20800
rect 23940 20748 23992 20800
rect 31944 20791 31996 20800
rect 31944 20757 31953 20791
rect 31953 20757 31987 20791
rect 31987 20757 31996 20791
rect 31944 20748 31996 20757
rect 33324 20748 33376 20800
rect 43812 20791 43864 20800
rect 43812 20757 43821 20791
rect 43821 20757 43855 20791
rect 43855 20757 43864 20791
rect 43812 20748 43864 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 3976 20544 4028 20596
rect 9404 20476 9456 20528
rect 10416 20408 10468 20460
rect 13084 20476 13136 20528
rect 12992 20408 13044 20460
rect 14188 20476 14240 20528
rect 14648 20476 14700 20528
rect 15660 20544 15712 20596
rect 17776 20544 17828 20596
rect 17960 20476 18012 20528
rect 20168 20476 20220 20528
rect 17224 20408 17276 20460
rect 17868 20408 17920 20460
rect 21088 20544 21140 20596
rect 21824 20544 21876 20596
rect 28540 20544 28592 20596
rect 30196 20587 30248 20596
rect 30196 20553 30205 20587
rect 30205 20553 30239 20587
rect 30239 20553 30248 20587
rect 30196 20544 30248 20553
rect 20444 20476 20496 20528
rect 27896 20476 27948 20528
rect 22376 20408 22428 20460
rect 23020 20408 23072 20460
rect 23204 20408 23256 20460
rect 26240 20451 26292 20460
rect 26240 20417 26249 20451
rect 26249 20417 26283 20451
rect 26283 20417 26292 20451
rect 26240 20408 26292 20417
rect 27436 20451 27488 20460
rect 27436 20417 27445 20451
rect 27445 20417 27479 20451
rect 27479 20417 27488 20451
rect 27436 20408 27488 20417
rect 27712 20408 27764 20460
rect 33324 20519 33376 20528
rect 33324 20485 33333 20519
rect 33333 20485 33367 20519
rect 33367 20485 33376 20519
rect 33324 20476 33376 20485
rect 43812 20519 43864 20528
rect 43812 20485 43821 20519
rect 43821 20485 43855 20519
rect 43855 20485 43864 20519
rect 43812 20476 43864 20485
rect 31944 20408 31996 20460
rect 46388 20451 46440 20460
rect 46388 20417 46397 20451
rect 46397 20417 46431 20451
rect 46431 20417 46440 20451
rect 46388 20408 46440 20417
rect 46940 20408 46992 20460
rect 47768 20451 47820 20460
rect 47768 20417 47777 20451
rect 47777 20417 47811 20451
rect 47811 20417 47820 20451
rect 47768 20408 47820 20417
rect 13912 20383 13964 20392
rect 13912 20349 13921 20383
rect 13921 20349 13955 20383
rect 13955 20349 13964 20383
rect 13912 20340 13964 20349
rect 17684 20383 17736 20392
rect 17684 20349 17693 20383
rect 17693 20349 17727 20383
rect 17727 20349 17736 20383
rect 17684 20340 17736 20349
rect 18052 20340 18104 20392
rect 19340 20340 19392 20392
rect 3240 20272 3292 20324
rect 8944 20204 8996 20256
rect 9956 20204 10008 20256
rect 13084 20247 13136 20256
rect 13084 20213 13093 20247
rect 13093 20213 13127 20247
rect 13127 20213 13136 20247
rect 13084 20204 13136 20213
rect 25964 20340 26016 20392
rect 35440 20340 35492 20392
rect 19984 20272 20036 20324
rect 24584 20272 24636 20324
rect 25044 20315 25096 20324
rect 25044 20281 25053 20315
rect 25053 20281 25087 20315
rect 25087 20281 25096 20315
rect 25044 20272 25096 20281
rect 26700 20272 26752 20324
rect 45468 20383 45520 20392
rect 45468 20349 45477 20383
rect 45477 20349 45511 20383
rect 45511 20349 45520 20383
rect 45468 20340 45520 20349
rect 45560 20340 45612 20392
rect 46756 20315 46808 20324
rect 46756 20281 46765 20315
rect 46765 20281 46799 20315
rect 46799 20281 46808 20315
rect 46756 20272 46808 20281
rect 20076 20247 20128 20256
rect 20076 20213 20085 20247
rect 20085 20213 20119 20247
rect 20119 20213 20128 20247
rect 20076 20204 20128 20213
rect 21916 20247 21968 20256
rect 21916 20213 21925 20247
rect 21925 20213 21959 20247
rect 21959 20213 21968 20247
rect 21916 20204 21968 20213
rect 23020 20204 23072 20256
rect 23388 20204 23440 20256
rect 27344 20204 27396 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 10600 20000 10652 20052
rect 13912 20000 13964 20052
rect 14556 20000 14608 20052
rect 20352 20000 20404 20052
rect 8944 19907 8996 19916
rect 8944 19873 8953 19907
rect 8953 19873 8987 19907
rect 8987 19873 8996 19907
rect 8944 19864 8996 19873
rect 11520 19864 11572 19916
rect 13176 19932 13228 19984
rect 14188 19932 14240 19984
rect 20076 19932 20128 19984
rect 21456 19932 21508 19984
rect 1768 19796 1820 19848
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 14464 19864 14516 19916
rect 17776 19864 17828 19916
rect 18052 19864 18104 19916
rect 20444 19864 20496 19916
rect 21916 19907 21968 19916
rect 21916 19873 21925 19907
rect 21925 19873 21959 19907
rect 21959 19873 21968 19907
rect 21916 19864 21968 19873
rect 9220 19771 9272 19780
rect 9220 19737 9229 19771
rect 9229 19737 9263 19771
rect 9263 19737 9272 19771
rect 9220 19728 9272 19737
rect 9956 19728 10008 19780
rect 13912 19796 13964 19848
rect 15660 19796 15712 19848
rect 17224 19839 17276 19848
rect 17224 19805 17233 19839
rect 17233 19805 17267 19839
rect 17267 19805 17276 19839
rect 17224 19796 17276 19805
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 13728 19728 13780 19780
rect 14188 19728 14240 19780
rect 17684 19728 17736 19780
rect 20352 19728 20404 19780
rect 11244 19703 11296 19712
rect 11244 19669 11253 19703
rect 11253 19669 11287 19703
rect 11287 19669 11296 19703
rect 11244 19660 11296 19669
rect 11336 19660 11388 19712
rect 13084 19660 13136 19712
rect 14096 19660 14148 19712
rect 15660 19660 15712 19712
rect 18420 19660 18472 19712
rect 20168 19660 20220 19712
rect 22192 19728 22244 19780
rect 23204 19660 23256 19712
rect 23388 20000 23440 20052
rect 24584 19864 24636 19916
rect 26056 19864 26108 19916
rect 27436 20000 27488 20052
rect 26516 19932 26568 19984
rect 41328 20000 41380 20052
rect 46940 20000 46992 20052
rect 27712 19975 27764 19984
rect 27712 19941 27721 19975
rect 27721 19941 27755 19975
rect 27755 19941 27764 19975
rect 27712 19932 27764 19941
rect 29184 19864 29236 19916
rect 45560 19864 45612 19916
rect 46572 19864 46624 19916
rect 25964 19839 26016 19848
rect 25964 19805 25973 19839
rect 25973 19805 26007 19839
rect 26007 19805 26016 19839
rect 25964 19796 26016 19805
rect 26424 19796 26476 19848
rect 26608 19839 26660 19848
rect 26608 19805 26617 19839
rect 26617 19805 26651 19839
rect 26651 19805 26660 19839
rect 26608 19796 26660 19805
rect 27160 19796 27212 19848
rect 27344 19796 27396 19848
rect 27528 19796 27580 19848
rect 28816 19839 28868 19848
rect 28816 19805 28825 19839
rect 28825 19805 28859 19839
rect 28859 19805 28868 19839
rect 28816 19796 28868 19805
rect 29000 19796 29052 19848
rect 44272 19839 44324 19848
rect 44272 19805 44281 19839
rect 44281 19805 44315 19839
rect 44315 19805 44324 19839
rect 44272 19796 44324 19805
rect 31392 19771 31444 19780
rect 31392 19737 31401 19771
rect 31401 19737 31435 19771
rect 31435 19737 31444 19771
rect 31392 19728 31444 19737
rect 46020 19796 46072 19848
rect 46388 19839 46440 19848
rect 46388 19805 46397 19839
rect 46397 19805 46431 19839
rect 46431 19805 46440 19839
rect 46388 19796 46440 19805
rect 46572 19728 46624 19780
rect 26240 19660 26292 19712
rect 27344 19660 27396 19712
rect 44272 19660 44324 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 2412 19456 2464 19508
rect 11244 19388 11296 19440
rect 12532 19388 12584 19440
rect 13176 19456 13228 19508
rect 19984 19456 20036 19508
rect 22192 19456 22244 19508
rect 13912 19431 13964 19440
rect 13912 19397 13921 19431
rect 13921 19397 13955 19431
rect 13955 19397 13964 19431
rect 13912 19388 13964 19397
rect 14280 19431 14332 19440
rect 14280 19397 14289 19431
rect 14289 19397 14323 19431
rect 14323 19397 14332 19431
rect 14280 19388 14332 19397
rect 16580 19388 16632 19440
rect 20076 19388 20128 19440
rect 20352 19388 20404 19440
rect 26516 19456 26568 19508
rect 26608 19456 26660 19508
rect 27344 19499 27396 19508
rect 27344 19465 27353 19499
rect 27353 19465 27387 19499
rect 27387 19465 27396 19499
rect 27344 19456 27396 19465
rect 29368 19456 29420 19508
rect 27528 19431 27580 19440
rect 27528 19397 27537 19431
rect 27537 19397 27571 19431
rect 27571 19397 27580 19431
rect 27528 19388 27580 19397
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 8852 19363 8904 19372
rect 8852 19329 8861 19363
rect 8861 19329 8895 19363
rect 8895 19329 8904 19363
rect 8852 19320 8904 19329
rect 10600 19320 10652 19372
rect 11336 19320 11388 19372
rect 14096 19363 14148 19372
rect 14096 19329 14105 19363
rect 14105 19329 14139 19363
rect 14139 19329 14148 19363
rect 14096 19320 14148 19329
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 17224 19320 17276 19372
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 20812 19320 20864 19372
rect 20996 19320 21048 19372
rect 21364 19320 21416 19372
rect 24584 19320 24636 19372
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 9220 19295 9272 19304
rect 9220 19261 9229 19295
rect 9229 19261 9263 19295
rect 9263 19261 9272 19295
rect 9220 19252 9272 19261
rect 13728 19252 13780 19304
rect 18696 19295 18748 19304
rect 18696 19261 18705 19295
rect 18705 19261 18739 19295
rect 18739 19261 18748 19295
rect 18696 19252 18748 19261
rect 18788 19252 18840 19304
rect 19064 19252 19116 19304
rect 19248 19252 19300 19304
rect 24032 19252 24084 19304
rect 25964 19320 26016 19372
rect 26424 19363 26476 19372
rect 26424 19329 26433 19363
rect 26433 19329 26467 19363
rect 26467 19329 26476 19363
rect 26424 19320 26476 19329
rect 26976 19320 27028 19372
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 39304 19431 39356 19440
rect 39304 19397 39313 19431
rect 39313 19397 39347 19431
rect 39347 19397 39356 19431
rect 39304 19388 39356 19397
rect 46848 19456 46900 19508
rect 42800 19320 42852 19372
rect 47216 19388 47268 19440
rect 11428 19184 11480 19236
rect 7564 19116 7616 19168
rect 18420 19184 18472 19236
rect 17316 19116 17368 19168
rect 21088 19184 21140 19236
rect 29368 19184 29420 19236
rect 20812 19159 20864 19168
rect 20812 19125 20821 19159
rect 20821 19125 20855 19159
rect 20855 19125 20864 19159
rect 20812 19116 20864 19125
rect 26884 19116 26936 19168
rect 30564 19184 30616 19236
rect 46940 19320 46992 19372
rect 47492 19320 47544 19372
rect 47768 19320 47820 19372
rect 46020 19252 46072 19304
rect 47032 19295 47084 19304
rect 47032 19261 47041 19295
rect 47041 19261 47075 19295
rect 47075 19261 47084 19295
rect 47032 19252 47084 19261
rect 47676 19159 47728 19168
rect 47676 19125 47685 19159
rect 47685 19125 47719 19159
rect 47719 19125 47728 19159
rect 47676 19116 47728 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 4896 18912 4948 18964
rect 12532 18912 12584 18964
rect 14188 18912 14240 18964
rect 14464 18955 14516 18964
rect 14464 18921 14473 18955
rect 14473 18921 14507 18955
rect 14507 18921 14516 18955
rect 14464 18912 14516 18921
rect 15200 18912 15252 18964
rect 18696 18912 18748 18964
rect 4896 18776 4948 18828
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 8208 18751 8260 18760
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 8852 18708 8904 18760
rect 13360 18776 13412 18828
rect 15200 18776 15252 18828
rect 19248 18819 19300 18828
rect 13084 18708 13136 18760
rect 15384 18751 15436 18760
rect 15384 18717 15393 18751
rect 15393 18717 15427 18751
rect 15427 18717 15436 18751
rect 15384 18708 15436 18717
rect 19248 18785 19257 18819
rect 19257 18785 19291 18819
rect 19291 18785 19300 18819
rect 19248 18776 19300 18785
rect 19432 18776 19484 18828
rect 19984 18776 20036 18828
rect 20720 18819 20772 18828
rect 20720 18785 20729 18819
rect 20729 18785 20763 18819
rect 20763 18785 20772 18819
rect 20720 18776 20772 18785
rect 21088 18776 21140 18828
rect 27160 18912 27212 18964
rect 14096 18683 14148 18692
rect 14096 18649 14105 18683
rect 14105 18649 14139 18683
rect 14139 18649 14148 18683
rect 14096 18640 14148 18649
rect 14648 18640 14700 18692
rect 17316 18683 17368 18692
rect 17316 18649 17325 18683
rect 17325 18649 17359 18683
rect 17359 18649 17368 18683
rect 17316 18640 17368 18649
rect 18236 18640 18288 18692
rect 19340 18708 19392 18760
rect 19432 18640 19484 18692
rect 12900 18572 12952 18624
rect 14280 18615 14332 18624
rect 14280 18581 14315 18615
rect 14315 18581 14332 18615
rect 14280 18572 14332 18581
rect 17684 18615 17736 18624
rect 17684 18581 17693 18615
rect 17693 18581 17727 18615
rect 17727 18581 17736 18615
rect 20536 18615 20588 18624
rect 17684 18572 17736 18581
rect 20536 18581 20545 18615
rect 20545 18581 20579 18615
rect 20579 18581 20588 18615
rect 20536 18572 20588 18581
rect 20904 18751 20956 18760
rect 20904 18717 20913 18751
rect 20913 18717 20947 18751
rect 20947 18717 20956 18751
rect 20904 18708 20956 18717
rect 22008 18708 22060 18760
rect 25044 18708 25096 18760
rect 26056 18751 26108 18760
rect 26056 18717 26065 18751
rect 26065 18717 26099 18751
rect 26099 18717 26108 18751
rect 26056 18708 26108 18717
rect 26884 18751 26936 18760
rect 26884 18717 26893 18751
rect 26893 18717 26927 18751
rect 26927 18717 26936 18751
rect 26884 18708 26936 18717
rect 47676 18776 47728 18828
rect 48136 18819 48188 18828
rect 48136 18785 48145 18819
rect 48145 18785 48179 18819
rect 48179 18785 48188 18819
rect 48136 18776 48188 18785
rect 27160 18708 27212 18760
rect 27620 18708 27672 18760
rect 27804 18640 27856 18692
rect 28080 18683 28132 18692
rect 28080 18649 28089 18683
rect 28089 18649 28123 18683
rect 28123 18649 28132 18683
rect 28080 18640 28132 18649
rect 29552 18640 29604 18692
rect 20996 18572 21048 18624
rect 22284 18615 22336 18624
rect 22284 18581 22293 18615
rect 22293 18581 22327 18615
rect 22327 18581 22336 18615
rect 22284 18572 22336 18581
rect 22468 18572 22520 18624
rect 23572 18572 23624 18624
rect 24492 18615 24544 18624
rect 24492 18581 24501 18615
rect 24501 18581 24535 18615
rect 24535 18581 24544 18615
rect 24492 18572 24544 18581
rect 26240 18572 26292 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 7564 18368 7616 18420
rect 2136 18300 2188 18352
rect 6644 18300 6696 18352
rect 13912 18300 13964 18352
rect 14464 18300 14516 18352
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 15108 18275 15160 18284
rect 15108 18241 15117 18275
rect 15117 18241 15151 18275
rect 15151 18241 15160 18275
rect 15108 18232 15160 18241
rect 17316 18300 17368 18352
rect 19340 18343 19392 18352
rect 19340 18309 19349 18343
rect 19349 18309 19383 18343
rect 19383 18309 19392 18343
rect 19340 18300 19392 18309
rect 20076 18343 20128 18352
rect 20076 18309 20085 18343
rect 20085 18309 20119 18343
rect 20119 18309 20128 18343
rect 20076 18300 20128 18309
rect 24492 18300 24544 18352
rect 15660 18232 15712 18284
rect 16120 18232 16172 18284
rect 19064 18232 19116 18284
rect 18788 18164 18840 18216
rect 19248 18275 19300 18284
rect 19248 18241 19257 18275
rect 19257 18241 19291 18275
rect 19291 18241 19300 18275
rect 19248 18232 19300 18241
rect 20168 18232 20220 18284
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 26608 18300 26660 18352
rect 26884 18300 26936 18352
rect 27160 18343 27212 18352
rect 27160 18309 27169 18343
rect 27169 18309 27203 18343
rect 27203 18309 27212 18343
rect 27160 18300 27212 18309
rect 28080 18368 28132 18420
rect 46940 18411 46992 18420
rect 46940 18377 46949 18411
rect 46949 18377 46983 18411
rect 46983 18377 46992 18411
rect 46940 18368 46992 18377
rect 26056 18275 26108 18284
rect 20812 18207 20864 18216
rect 20812 18173 20821 18207
rect 20821 18173 20855 18207
rect 20855 18173 20864 18207
rect 20812 18164 20864 18173
rect 14648 18071 14700 18080
rect 14648 18037 14657 18071
rect 14657 18037 14691 18071
rect 14691 18037 14700 18071
rect 14648 18028 14700 18037
rect 15384 18028 15436 18080
rect 18144 18028 18196 18080
rect 19340 18028 19392 18080
rect 19524 18071 19576 18080
rect 19524 18037 19533 18071
rect 19533 18037 19567 18071
rect 19567 18037 19576 18071
rect 19524 18028 19576 18037
rect 26056 18241 26065 18275
rect 26065 18241 26099 18275
rect 26099 18241 26108 18275
rect 26056 18232 26108 18241
rect 26240 18275 26292 18284
rect 26240 18241 26249 18275
rect 26249 18241 26283 18275
rect 26283 18241 26292 18275
rect 26240 18232 26292 18241
rect 32772 18232 32824 18284
rect 46848 18275 46900 18284
rect 46848 18241 46857 18275
rect 46857 18241 46891 18275
rect 46891 18241 46900 18275
rect 46848 18232 46900 18241
rect 47216 18232 47268 18284
rect 47492 18232 47544 18284
rect 47768 18275 47820 18284
rect 47768 18241 47777 18275
rect 47777 18241 47811 18275
rect 47811 18241 47820 18275
rect 47768 18232 47820 18241
rect 26424 18164 26476 18216
rect 27804 18207 27856 18216
rect 27804 18173 27813 18207
rect 27813 18173 27847 18207
rect 27847 18173 27856 18207
rect 27804 18164 27856 18173
rect 28080 18164 28132 18216
rect 27436 18096 27488 18148
rect 29000 18096 29052 18148
rect 28724 18071 28776 18080
rect 28724 18037 28733 18071
rect 28733 18037 28767 18071
rect 28767 18037 28776 18071
rect 28724 18028 28776 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 15108 17824 15160 17876
rect 19432 17824 19484 17876
rect 21364 17867 21416 17876
rect 21364 17833 21373 17867
rect 21373 17833 21407 17867
rect 21407 17833 21416 17867
rect 21364 17824 21416 17833
rect 24032 17824 24084 17876
rect 26424 17867 26476 17876
rect 26424 17833 26433 17867
rect 26433 17833 26467 17867
rect 26467 17833 26476 17867
rect 26424 17824 26476 17833
rect 47216 17824 47268 17876
rect 20536 17756 20588 17808
rect 3976 17688 4028 17740
rect 14648 17688 14700 17740
rect 17868 17688 17920 17740
rect 19340 17688 19392 17740
rect 19524 17688 19576 17740
rect 20812 17688 20864 17740
rect 22284 17688 22336 17740
rect 14372 17663 14424 17672
rect 14372 17629 14381 17663
rect 14381 17629 14415 17663
rect 14415 17629 14424 17663
rect 14372 17620 14424 17629
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 11704 17552 11756 17604
rect 15200 17552 15252 17604
rect 17224 17595 17276 17604
rect 17224 17561 17233 17595
rect 17233 17561 17267 17595
rect 17267 17561 17276 17595
rect 17224 17552 17276 17561
rect 17776 17552 17828 17604
rect 19248 17552 19300 17604
rect 27436 17620 27488 17672
rect 28080 17663 28132 17672
rect 28080 17629 28089 17663
rect 28089 17629 28123 17663
rect 28123 17629 28132 17663
rect 28080 17620 28132 17629
rect 47032 17620 47084 17672
rect 11980 17484 12032 17536
rect 14188 17484 14240 17536
rect 18144 17527 18196 17536
rect 18144 17493 18153 17527
rect 18153 17493 18187 17527
rect 18187 17493 18196 17527
rect 22192 17552 22244 17604
rect 23572 17552 23624 17604
rect 25688 17552 25740 17604
rect 26056 17595 26108 17604
rect 26056 17561 26065 17595
rect 26065 17561 26099 17595
rect 26099 17561 26108 17595
rect 26056 17552 26108 17561
rect 26240 17595 26292 17604
rect 26240 17561 26249 17595
rect 26249 17561 26283 17595
rect 26283 17561 26292 17595
rect 26240 17552 26292 17561
rect 27712 17552 27764 17604
rect 47768 17620 47820 17672
rect 47492 17552 47544 17604
rect 48044 17552 48096 17604
rect 18144 17484 18196 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 11704 17323 11756 17332
rect 11704 17289 11713 17323
rect 11713 17289 11747 17323
rect 11747 17289 11756 17323
rect 11704 17280 11756 17289
rect 13912 17280 13964 17332
rect 15200 17323 15252 17332
rect 15200 17289 15209 17323
rect 15209 17289 15243 17323
rect 15243 17289 15252 17323
rect 15200 17280 15252 17289
rect 19064 17280 19116 17332
rect 19984 17280 20036 17332
rect 22008 17323 22060 17332
rect 22008 17289 22017 17323
rect 22017 17289 22051 17323
rect 22051 17289 22060 17323
rect 22008 17280 22060 17289
rect 8208 17144 8260 17196
rect 17316 17212 17368 17264
rect 17776 17212 17828 17264
rect 18144 17212 18196 17264
rect 28724 17212 28776 17264
rect 11060 17144 11112 17196
rect 11612 17187 11664 17196
rect 11612 17153 11621 17187
rect 11621 17153 11655 17187
rect 11655 17153 11664 17187
rect 11612 17144 11664 17153
rect 10416 17119 10468 17128
rect 10416 17085 10425 17119
rect 10425 17085 10459 17119
rect 10459 17085 10468 17119
rect 10416 17076 10468 17085
rect 8208 17008 8260 17060
rect 13360 17144 13412 17196
rect 14832 17144 14884 17196
rect 15660 17144 15712 17196
rect 19984 17144 20036 17196
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 47584 17187 47636 17196
rect 47584 17153 47593 17187
rect 47593 17153 47627 17187
rect 47627 17153 47636 17187
rect 47584 17144 47636 17153
rect 16580 17076 16632 17128
rect 27712 17119 27764 17128
rect 27712 17085 27721 17119
rect 27721 17085 27755 17119
rect 27755 17085 27764 17119
rect 27712 17076 27764 17085
rect 28172 17119 28224 17128
rect 28172 17085 28181 17119
rect 28181 17085 28215 17119
rect 28215 17085 28224 17119
rect 28172 17076 28224 17085
rect 18236 17008 18288 17060
rect 1400 16940 1452 16992
rect 11612 16940 11664 16992
rect 15660 16940 15712 16992
rect 15752 16940 15804 16992
rect 18512 16940 18564 16992
rect 19432 16940 19484 16992
rect 46296 16940 46348 16992
rect 47676 16983 47728 16992
rect 47676 16949 47685 16983
rect 47685 16949 47719 16983
rect 47719 16949 47728 16983
rect 47676 16940 47728 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3332 16736 3384 16788
rect 28172 16736 28224 16788
rect 18052 16668 18104 16720
rect 18328 16668 18380 16720
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 19340 16643 19392 16652
rect 15108 16532 15160 16584
rect 17224 16532 17276 16584
rect 19340 16609 19349 16643
rect 19349 16609 19383 16643
rect 19383 16609 19392 16643
rect 19340 16600 19392 16609
rect 19984 16600 20036 16652
rect 46296 16643 46348 16652
rect 46296 16609 46305 16643
rect 46305 16609 46339 16643
rect 46339 16609 46348 16643
rect 46296 16600 46348 16609
rect 48136 16643 48188 16652
rect 48136 16609 48145 16643
rect 48145 16609 48179 16643
rect 48179 16609 48188 16643
rect 48136 16600 48188 16609
rect 2136 16464 2188 16516
rect 17500 16464 17552 16516
rect 18144 16507 18196 16516
rect 18144 16473 18153 16507
rect 18153 16473 18187 16507
rect 18187 16473 18196 16507
rect 18144 16464 18196 16473
rect 18512 16532 18564 16584
rect 19248 16532 19300 16584
rect 21824 16464 21876 16516
rect 17960 16396 18012 16448
rect 18512 16396 18564 16448
rect 20444 16439 20496 16448
rect 20444 16405 20453 16439
rect 20453 16405 20487 16439
rect 20487 16405 20496 16439
rect 20444 16396 20496 16405
rect 47676 16464 47728 16516
rect 45560 16396 45612 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 14188 16192 14240 16244
rect 15108 16192 15160 16244
rect 18144 16192 18196 16244
rect 19248 16192 19300 16244
rect 19984 16124 20036 16176
rect 2044 16056 2096 16065
rect 14924 16056 14976 16108
rect 18604 16056 18656 16108
rect 19432 16099 19484 16108
rect 19432 16065 19441 16099
rect 19441 16065 19475 16099
rect 19475 16065 19484 16099
rect 19432 16056 19484 16065
rect 20812 16056 20864 16108
rect 47124 16056 47176 16108
rect 13544 16031 13596 16040
rect 12716 15852 12768 15904
rect 13544 15997 13553 16031
rect 13553 15997 13587 16031
rect 13587 15997 13596 16031
rect 13544 15988 13596 15997
rect 17224 16031 17276 16040
rect 17224 15997 17233 16031
rect 17233 15997 17267 16031
rect 17267 15997 17276 16031
rect 17224 15988 17276 15997
rect 18052 15988 18104 16040
rect 18972 15988 19024 16040
rect 28816 15988 28868 16040
rect 14372 15852 14424 15904
rect 46296 15852 46348 15904
rect 47676 15895 47728 15904
rect 47676 15861 47685 15895
rect 47685 15861 47719 15895
rect 47719 15861 47728 15895
rect 47676 15852 47728 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 13544 15648 13596 15700
rect 14924 15691 14976 15700
rect 14924 15657 14933 15691
rect 14933 15657 14967 15691
rect 14967 15657 14976 15691
rect 14924 15648 14976 15657
rect 18604 15648 18656 15700
rect 20812 15648 20864 15700
rect 12716 15580 12768 15632
rect 18880 15580 18932 15632
rect 18144 15512 18196 15564
rect 46296 15555 46348 15564
rect 46296 15521 46305 15555
rect 46305 15521 46339 15555
rect 46339 15521 46348 15555
rect 46296 15512 46348 15521
rect 47676 15512 47728 15564
rect 48136 15555 48188 15564
rect 48136 15521 48145 15555
rect 48145 15521 48179 15555
rect 48179 15521 48188 15555
rect 48136 15512 48188 15521
rect 1768 15444 1820 15496
rect 14280 15487 14332 15496
rect 14280 15453 14289 15487
rect 14289 15453 14323 15487
rect 14323 15453 14332 15487
rect 14280 15444 14332 15453
rect 14832 15487 14884 15496
rect 14832 15453 14841 15487
rect 14841 15453 14875 15487
rect 14875 15453 14884 15487
rect 14832 15444 14884 15453
rect 19248 15487 19300 15496
rect 19248 15453 19257 15487
rect 19257 15453 19291 15487
rect 19291 15453 19300 15487
rect 19248 15444 19300 15453
rect 20168 15444 20220 15496
rect 18144 15376 18196 15428
rect 16304 15308 16356 15360
rect 18972 15308 19024 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 17224 15104 17276 15156
rect 18052 15147 18104 15156
rect 18052 15113 18061 15147
rect 18061 15113 18095 15147
rect 18095 15113 18104 15147
rect 18052 15104 18104 15113
rect 17868 15036 17920 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 14832 15011 14884 15020
rect 14832 14977 14841 15011
rect 14841 14977 14875 15011
rect 14875 14977 14884 15011
rect 14832 14968 14884 14977
rect 17776 14968 17828 15020
rect 17960 15011 18012 15020
rect 17960 14977 17969 15011
rect 17969 14977 18003 15011
rect 18003 14977 18012 15011
rect 17960 14968 18012 14977
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 15016 14764 15068 14816
rect 17224 14764 17276 14816
rect 17592 14764 17644 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 17316 14560 17368 14612
rect 17224 14492 17276 14544
rect 2688 14356 2740 14408
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 14372 14356 14424 14408
rect 17776 14424 17828 14476
rect 16028 14356 16080 14408
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 20444 14424 20496 14476
rect 19248 14399 19300 14408
rect 19248 14365 19257 14399
rect 19257 14365 19291 14399
rect 19291 14365 19300 14399
rect 19248 14356 19300 14365
rect 17224 14331 17276 14340
rect 17224 14297 17233 14331
rect 17233 14297 17267 14331
rect 17267 14297 17276 14331
rect 17224 14288 17276 14297
rect 17868 14288 17920 14340
rect 14280 14220 14332 14272
rect 15200 14263 15252 14272
rect 15200 14229 15209 14263
rect 15209 14229 15243 14263
rect 15243 14229 15252 14263
rect 15200 14220 15252 14229
rect 15844 14220 15896 14272
rect 17960 14220 18012 14272
rect 19432 14220 19484 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 16028 14059 16080 14068
rect 16028 14025 16037 14059
rect 16037 14025 16071 14059
rect 16071 14025 16080 14059
rect 16028 14016 16080 14025
rect 17684 14016 17736 14068
rect 15016 13948 15068 14000
rect 17316 13948 17368 14000
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 17868 13812 17920 13864
rect 20076 13948 20128 14000
rect 47124 13880 47176 13932
rect 19340 13812 19392 13864
rect 3976 13676 4028 13728
rect 4620 13676 4672 13728
rect 15200 13676 15252 13728
rect 17224 13719 17276 13728
rect 17224 13685 17233 13719
rect 17233 13685 17267 13719
rect 17267 13685 17276 13719
rect 17224 13676 17276 13685
rect 47676 13719 47728 13728
rect 47676 13685 47685 13719
rect 47685 13685 47719 13719
rect 47719 13685 47728 13719
rect 47676 13676 47728 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 12440 13472 12492 13524
rect 16028 13404 16080 13456
rect 15844 13379 15896 13388
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 19340 13472 19392 13524
rect 20076 13472 20128 13524
rect 19248 13404 19300 13456
rect 17408 13336 17460 13388
rect 17224 13268 17276 13320
rect 18236 13268 18288 13320
rect 47676 13336 47728 13388
rect 46296 13311 46348 13320
rect 16856 13200 16908 13252
rect 46296 13277 46305 13311
rect 46305 13277 46339 13311
rect 46339 13277 46348 13311
rect 46296 13268 46348 13277
rect 20444 13200 20496 13252
rect 48136 13243 48188 13252
rect 48136 13209 48145 13243
rect 48145 13209 48179 13243
rect 48179 13209 48188 13243
rect 48136 13200 48188 13209
rect 18144 13132 18196 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 17408 12971 17460 12980
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 17868 12928 17920 12980
rect 18236 12928 18288 12980
rect 18144 12903 18196 12912
rect 18144 12869 18153 12903
rect 18153 12869 18187 12903
rect 18187 12869 18196 12903
rect 18144 12860 18196 12869
rect 19432 12860 19484 12912
rect 17316 12792 17368 12844
rect 17868 12835 17920 12844
rect 17868 12801 17877 12835
rect 17877 12801 17911 12835
rect 17911 12801 17920 12835
rect 17868 12792 17920 12801
rect 46296 12792 46348 12844
rect 25596 12724 25648 12776
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 41604 12180 41656 12232
rect 46480 12044 46532 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 17960 11840 18012 11892
rect 20628 11840 20680 11892
rect 16580 11772 16632 11824
rect 17960 11704 18012 11756
rect 17316 11636 17368 11688
rect 27620 11636 27672 11688
rect 17040 11500 17092 11552
rect 46296 11500 46348 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 14832 11228 14884 11280
rect 16856 11203 16908 11212
rect 16856 11169 16865 11203
rect 16865 11169 16899 11203
rect 16899 11169 16908 11203
rect 16856 11160 16908 11169
rect 17040 11203 17092 11212
rect 17040 11169 17049 11203
rect 17049 11169 17083 11203
rect 17083 11169 17092 11203
rect 17040 11160 17092 11169
rect 46296 11203 46348 11212
rect 46296 11169 46305 11203
rect 46305 11169 46339 11203
rect 46339 11169 46348 11203
rect 46296 11160 46348 11169
rect 46480 11203 46532 11212
rect 46480 11169 46489 11203
rect 46489 11169 46523 11203
rect 46523 11169 46532 11203
rect 46480 11160 46532 11169
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 2780 10956 2832 11008
rect 4896 10956 4948 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 18512 10684 18564 10736
rect 46112 10727 46164 10736
rect 46112 10693 46121 10727
rect 46121 10693 46155 10727
rect 46155 10693 46164 10727
rect 46112 10684 46164 10693
rect 18144 10548 18196 10600
rect 46020 10591 46072 10600
rect 3516 10480 3568 10532
rect 46020 10557 46029 10591
rect 46029 10557 46063 10591
rect 46063 10557 46072 10591
rect 46020 10548 46072 10557
rect 45928 10480 45980 10532
rect 46296 10412 46348 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 17960 10004 18012 10056
rect 47676 9936 47728 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 46112 9664 46164 9716
rect 47676 9639 47728 9648
rect 47676 9605 47685 9639
rect 47685 9605 47719 9639
rect 47719 9605 47728 9639
rect 47676 9596 47728 9605
rect 46848 9528 46900 9580
rect 47492 9528 47544 9580
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 47308 8959 47360 8968
rect 47308 8925 47317 8959
rect 47317 8925 47351 8959
rect 47351 8925 47360 8959
rect 47308 8916 47360 8925
rect 47400 8916 47452 8968
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 47676 8483 47728 8492
rect 47676 8449 47685 8483
rect 47685 8449 47719 8483
rect 47719 8449 47728 8483
rect 47676 8440 47728 8449
rect 24952 8372 25004 8424
rect 3424 8236 3476 8288
rect 12440 8236 12492 8288
rect 17500 8236 17552 8288
rect 45560 8236 45612 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 47860 7964 47912 8016
rect 47400 7896 47452 7948
rect 47676 7939 47728 7948
rect 47676 7905 47685 7939
rect 47685 7905 47719 7939
rect 47719 7905 47728 7939
rect 47676 7896 47728 7905
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 48136 7395 48188 7404
rect 48136 7361 48145 7395
rect 48145 7361 48179 7395
rect 48179 7361 48188 7395
rect 48136 7352 48188 7361
rect 47032 7148 47084 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3516 6808 3568 6860
rect 18144 6808 18196 6860
rect 47032 6851 47084 6860
rect 47032 6817 47041 6851
rect 47041 6817 47075 6851
rect 47075 6817 47084 6851
rect 47032 6808 47084 6817
rect 48044 6851 48096 6860
rect 48044 6817 48053 6851
rect 48053 6817 48087 6851
rect 48087 6817 48096 6851
rect 48044 6808 48096 6817
rect 1676 6672 1728 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 46572 6264 46624 6316
rect 48136 6307 48188 6316
rect 48136 6273 48145 6307
rect 48145 6273 48179 6307
rect 48179 6273 48188 6307
rect 48136 6264 48188 6273
rect 46204 6239 46256 6248
rect 46204 6205 46213 6239
rect 46213 6205 46247 6239
rect 46247 6205 46256 6239
rect 46204 6196 46256 6205
rect 47952 6103 48004 6112
rect 47952 6069 47961 6103
rect 47961 6069 47995 6103
rect 47995 6069 48004 6103
rect 47952 6060 48004 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 44364 5720 44416 5772
rect 47676 5763 47728 5772
rect 47676 5729 47685 5763
rect 47685 5729 47719 5763
rect 47719 5729 47728 5763
rect 47676 5720 47728 5729
rect 27712 5652 27764 5704
rect 46480 5627 46532 5636
rect 46480 5593 46489 5627
rect 46489 5593 46523 5627
rect 46523 5593 46532 5627
rect 46480 5584 46532 5593
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 46020 5287 46072 5296
rect 46020 5253 46029 5287
rect 46029 5253 46063 5287
rect 46063 5253 46072 5287
rect 46020 5244 46072 5253
rect 47952 5244 48004 5296
rect 47768 5176 47820 5228
rect 48044 5108 48096 5160
rect 47676 5015 47728 5024
rect 47676 4981 47685 5015
rect 47685 4981 47719 5015
rect 47719 4981 47728 5015
rect 47676 4972 47728 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 43536 4632 43588 4684
rect 46020 4632 46072 4684
rect 46572 4675 46624 4684
rect 46572 4641 46581 4675
rect 46581 4641 46615 4675
rect 46615 4641 46624 4675
rect 46572 4632 46624 4641
rect 7656 4564 7708 4616
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 20260 4564 20312 4616
rect 20812 4564 20864 4616
rect 20996 4607 21048 4616
rect 20996 4573 21005 4607
rect 21005 4573 21039 4607
rect 21039 4573 21048 4607
rect 20996 4564 21048 4573
rect 20904 4496 20956 4548
rect 23572 4564 23624 4616
rect 42892 4607 42944 4616
rect 42892 4573 42901 4607
rect 42901 4573 42935 4607
rect 42935 4573 42944 4607
rect 42892 4564 42944 4573
rect 45652 4607 45704 4616
rect 45652 4573 45661 4607
rect 45661 4573 45695 4607
rect 45695 4573 45704 4607
rect 45652 4564 45704 4573
rect 22744 4496 22796 4548
rect 46296 4539 46348 4548
rect 46296 4505 46305 4539
rect 46305 4505 46339 4539
rect 46339 4505 46348 4539
rect 46296 4496 46348 4505
rect 19432 4428 19484 4480
rect 20720 4428 20772 4480
rect 21364 4428 21416 4480
rect 22836 4428 22888 4480
rect 23020 4471 23072 4480
rect 23020 4437 23029 4471
rect 23029 4437 23063 4471
rect 23063 4437 23072 4471
rect 23020 4428 23072 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 20260 4224 20312 4276
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 18972 4088 19024 4140
rect 19524 4088 19576 4140
rect 19708 4131 19760 4140
rect 19708 4097 19717 4131
rect 19717 4097 19751 4131
rect 19751 4097 19760 4131
rect 19708 4088 19760 4097
rect 14096 4020 14148 4072
rect 18420 4020 18472 4072
rect 20904 4088 20956 4140
rect 20812 4020 20864 4072
rect 22376 4088 22428 4140
rect 22836 4131 22888 4140
rect 22836 4097 22845 4131
rect 22845 4097 22879 4131
rect 22879 4097 22888 4131
rect 22836 4088 22888 4097
rect 23480 4131 23532 4140
rect 22468 4020 22520 4072
rect 22560 4020 22612 4072
rect 23480 4097 23489 4131
rect 23489 4097 23523 4131
rect 23523 4097 23532 4131
rect 23480 4088 23532 4097
rect 23572 4131 23624 4140
rect 23572 4097 23581 4131
rect 23581 4097 23615 4131
rect 23615 4097 23624 4131
rect 23572 4088 23624 4097
rect 23204 4020 23256 4072
rect 26240 4088 26292 4140
rect 24400 4020 24452 4072
rect 28540 4020 28592 4072
rect 29460 4063 29512 4072
rect 29460 4029 29469 4063
rect 29469 4029 29503 4063
rect 29503 4029 29512 4063
rect 29460 4020 29512 4029
rect 30012 4020 30064 4072
rect 45744 4156 45796 4208
rect 46572 4156 46624 4208
rect 47768 4199 47820 4208
rect 47768 4165 47777 4199
rect 47777 4165 47811 4199
rect 47811 4165 47820 4199
rect 47768 4156 47820 4165
rect 39212 4088 39264 4140
rect 43444 4088 43496 4140
rect 46480 4131 46532 4140
rect 46480 4097 46489 4131
rect 46489 4097 46523 4131
rect 46523 4097 46532 4131
rect 46480 4088 46532 4097
rect 41328 4020 41380 4072
rect 43536 4063 43588 4072
rect 43536 4029 43545 4063
rect 43545 4029 43579 4063
rect 43579 4029 43588 4063
rect 43536 4020 43588 4029
rect 43720 4063 43772 4072
rect 43720 4029 43729 4063
rect 43729 4029 43763 4063
rect 43763 4029 43772 4063
rect 43720 4020 43772 4029
rect 43812 4020 43864 4072
rect 48320 4020 48372 4072
rect 19984 3952 20036 4004
rect 23112 3952 23164 4004
rect 1584 3884 1636 3936
rect 2780 3884 2832 3936
rect 6736 3927 6788 3936
rect 6736 3893 6745 3927
rect 6745 3893 6779 3927
rect 6779 3893 6788 3927
rect 6736 3884 6788 3893
rect 7472 3927 7524 3936
rect 7472 3893 7481 3927
rect 7481 3893 7515 3927
rect 7515 3893 7524 3927
rect 7472 3884 7524 3893
rect 7840 3884 7892 3936
rect 9220 3884 9272 3936
rect 11520 3884 11572 3936
rect 19064 3884 19116 3936
rect 20260 3884 20312 3936
rect 20536 3884 20588 3936
rect 21732 3884 21784 3936
rect 22376 3884 22428 3936
rect 24676 3884 24728 3936
rect 26884 3952 26936 4004
rect 33968 3952 34020 4004
rect 40040 3927 40092 3936
rect 40040 3893 40049 3927
rect 40049 3893 40083 3927
rect 40083 3893 40092 3927
rect 40040 3884 40092 3893
rect 42800 3884 42852 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 6920 3680 6972 3732
rect 15292 3680 15344 3732
rect 19524 3723 19576 3732
rect 19524 3689 19533 3723
rect 19533 3689 19567 3723
rect 19567 3689 19576 3723
rect 19524 3680 19576 3689
rect 19708 3680 19760 3732
rect 20996 3680 21048 3732
rect 9036 3612 9088 3664
rect 1768 3544 1820 3596
rect 6736 3587 6788 3596
rect 6736 3553 6745 3587
rect 6745 3553 6779 3587
rect 6779 3553 6788 3587
rect 6736 3544 6788 3553
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 9220 3587 9272 3596
rect 9220 3553 9229 3587
rect 9229 3553 9263 3587
rect 9263 3553 9272 3587
rect 9220 3544 9272 3553
rect 9956 3612 10008 3664
rect 19892 3612 19944 3664
rect 22560 3680 22612 3732
rect 22744 3680 22796 3732
rect 23388 3680 23440 3732
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 19248 3544 19300 3596
rect 13820 3476 13872 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 17960 3476 18012 3528
rect 18604 3476 18656 3528
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 22192 3612 22244 3664
rect 28540 3680 28592 3732
rect 20168 3544 20220 3596
rect 21456 3544 21508 3596
rect 21548 3544 21600 3596
rect 1308 3408 1360 3460
rect 1952 3340 2004 3392
rect 10048 3408 10100 3460
rect 15476 3451 15528 3460
rect 11704 3340 11756 3392
rect 14004 3340 14056 3392
rect 15476 3417 15485 3451
rect 15485 3417 15519 3451
rect 15519 3417 15528 3451
rect 15476 3408 15528 3417
rect 17132 3451 17184 3460
rect 17132 3417 17141 3451
rect 17141 3417 17175 3451
rect 17175 3417 17184 3451
rect 17132 3408 17184 3417
rect 20260 3476 20312 3528
rect 20720 3519 20772 3528
rect 20720 3485 20729 3519
rect 20729 3485 20763 3519
rect 20763 3485 20772 3519
rect 20720 3476 20772 3485
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 22100 3476 22152 3528
rect 22836 3519 22888 3528
rect 22836 3485 22845 3519
rect 22845 3485 22879 3519
rect 22879 3485 22888 3519
rect 22836 3476 22888 3485
rect 20168 3408 20220 3460
rect 24584 3408 24636 3460
rect 33048 3612 33100 3664
rect 33968 3680 34020 3732
rect 29552 3587 29604 3596
rect 29552 3553 29561 3587
rect 29561 3553 29595 3587
rect 29595 3553 29604 3587
rect 29552 3544 29604 3553
rect 33048 3519 33100 3528
rect 33048 3485 33057 3519
rect 33057 3485 33091 3519
rect 33091 3485 33100 3519
rect 33048 3476 33100 3485
rect 18328 3340 18380 3392
rect 19156 3340 19208 3392
rect 19248 3340 19300 3392
rect 20536 3340 20588 3392
rect 20628 3340 20680 3392
rect 21732 3340 21784 3392
rect 23388 3340 23440 3392
rect 23664 3340 23716 3392
rect 24768 3383 24820 3392
rect 24768 3349 24777 3383
rect 24777 3349 24811 3383
rect 24811 3349 24820 3383
rect 24768 3340 24820 3349
rect 24860 3340 24912 3392
rect 31300 3340 31352 3392
rect 32956 3408 33008 3460
rect 32864 3340 32916 3392
rect 33140 3383 33192 3392
rect 33140 3349 33149 3383
rect 33149 3349 33183 3383
rect 33183 3349 33192 3383
rect 33140 3340 33192 3349
rect 35440 3612 35492 3664
rect 42524 3612 42576 3664
rect 42892 3612 42944 3664
rect 43444 3680 43496 3732
rect 46664 3680 46716 3732
rect 47216 3612 47268 3664
rect 35900 3519 35952 3528
rect 35900 3485 35909 3519
rect 35909 3485 35943 3519
rect 35943 3485 35952 3519
rect 35900 3476 35952 3485
rect 39120 3519 39172 3528
rect 39120 3485 39129 3519
rect 39129 3485 39163 3519
rect 39163 3485 39172 3519
rect 39120 3476 39172 3485
rect 39948 3476 40000 3528
rect 41328 3519 41380 3528
rect 36176 3408 36228 3460
rect 37924 3340 37976 3392
rect 39856 3408 39908 3460
rect 41328 3485 41337 3519
rect 41337 3485 41371 3519
rect 41371 3485 41380 3519
rect 41328 3476 41380 3485
rect 41512 3519 41564 3528
rect 41512 3485 41521 3519
rect 41521 3485 41555 3519
rect 41555 3485 41564 3519
rect 41512 3476 41564 3485
rect 42800 3587 42852 3596
rect 42800 3553 42809 3587
rect 42809 3553 42843 3587
rect 42843 3553 42852 3587
rect 42800 3544 42852 3553
rect 43168 3587 43220 3596
rect 43168 3553 43177 3587
rect 43177 3553 43211 3587
rect 43211 3553 43220 3587
rect 43168 3544 43220 3553
rect 47676 3544 47728 3596
rect 44272 3408 44324 3460
rect 47492 3408 47544 3460
rect 48964 3408 49016 3460
rect 40132 3340 40184 3392
rect 42432 3340 42484 3392
rect 45376 3340 45428 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3884 3136 3936 3188
rect 17960 3179 18012 3188
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 7840 3111 7892 3120
rect 7840 3077 7849 3111
rect 7849 3077 7883 3111
rect 7883 3077 7892 3111
rect 7840 3068 7892 3077
rect 10048 3111 10100 3120
rect 10048 3077 10057 3111
rect 10057 3077 10091 3111
rect 10091 3077 10100 3111
rect 10048 3068 10100 3077
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 14004 3111 14056 3120
rect 14004 3077 14013 3111
rect 14013 3077 14047 3111
rect 14047 3077 14056 3111
rect 14004 3068 14056 3077
rect 17960 3145 17969 3179
rect 17969 3145 18003 3179
rect 18003 3145 18012 3179
rect 17960 3136 18012 3145
rect 18604 3179 18656 3188
rect 18604 3145 18613 3179
rect 18613 3145 18647 3179
rect 18647 3145 18656 3179
rect 18604 3136 18656 3145
rect 18972 3136 19024 3188
rect 20168 3136 20220 3188
rect 20720 3179 20772 3188
rect 20720 3145 20729 3179
rect 20729 3145 20763 3179
rect 20763 3145 20772 3179
rect 20720 3136 20772 3145
rect 36176 3179 36228 3188
rect 22376 3068 22428 3120
rect 22468 3068 22520 3120
rect 24768 3111 24820 3120
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 9956 3043 10008 3052
rect 9956 3009 9965 3043
rect 9965 3009 9999 3043
rect 9999 3009 10008 3043
rect 9956 3000 10008 3009
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 17316 3000 17368 3052
rect 664 2932 716 2984
rect 10968 2932 11020 2984
rect 14188 2932 14240 2984
rect 15200 2932 15252 2984
rect 18328 3000 18380 3052
rect 19156 3043 19208 3052
rect 19156 3009 19165 3043
rect 19165 3009 19199 3043
rect 19199 3009 19208 3043
rect 19156 3000 19208 3009
rect 19984 3043 20036 3052
rect 19984 3009 19993 3043
rect 19993 3009 20027 3043
rect 20027 3009 20036 3043
rect 19984 3000 20036 3009
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 17684 2932 17736 2984
rect 21548 2932 21600 2984
rect 22100 2975 22152 2984
rect 22100 2941 22114 2975
rect 22114 2941 22148 2975
rect 22148 2941 22152 2975
rect 22100 2932 22152 2941
rect 7748 2864 7800 2916
rect 14096 2864 14148 2916
rect 22468 2864 22520 2916
rect 22560 2864 22612 2916
rect 24768 3077 24777 3111
rect 24777 3077 24811 3111
rect 24811 3077 24820 3111
rect 24768 3068 24820 3077
rect 27988 3068 28040 3120
rect 33140 3111 33192 3120
rect 33140 3077 33149 3111
rect 33149 3077 33183 3111
rect 33183 3077 33192 3111
rect 33140 3068 33192 3077
rect 36176 3145 36185 3179
rect 36185 3145 36219 3179
rect 36219 3145 36228 3179
rect 36176 3136 36228 3145
rect 38568 3136 38620 3188
rect 41236 3136 41288 3188
rect 45284 3136 45336 3188
rect 41512 3068 41564 3120
rect 24584 3043 24636 3052
rect 24584 3009 24593 3043
rect 24593 3009 24627 3043
rect 24627 3009 24636 3043
rect 24584 3000 24636 3009
rect 27068 3000 27120 3052
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 32220 3000 32272 3052
rect 32956 3043 33008 3052
rect 32956 3009 32965 3043
rect 32965 3009 32999 3043
rect 32999 3009 33008 3043
rect 32956 3000 33008 3009
rect 36084 3000 36136 3052
rect 37924 3043 37976 3052
rect 37924 3009 37933 3043
rect 37933 3009 37967 3043
rect 37967 3009 37976 3043
rect 37924 3000 37976 3009
rect 42432 3043 42484 3052
rect 42432 3009 42441 3043
rect 42441 3009 42475 3043
rect 42475 3009 42484 3043
rect 42432 3000 42484 3009
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 35900 2932 35952 2984
rect 38568 2975 38620 2984
rect 38568 2941 38577 2975
rect 38577 2941 38611 2975
rect 38611 2941 38620 2975
rect 38568 2932 38620 2941
rect 39856 2975 39908 2984
rect 39856 2941 39865 2975
rect 39865 2941 39899 2975
rect 39899 2941 39908 2975
rect 39856 2932 39908 2941
rect 29092 2864 29144 2916
rect 39028 2864 39080 2916
rect 39212 2907 39264 2916
rect 39212 2873 39221 2907
rect 39221 2873 39255 2907
rect 39255 2873 39264 2907
rect 39212 2864 39264 2873
rect 6828 2839 6880 2848
rect 6828 2805 6837 2839
rect 6837 2805 6871 2839
rect 6871 2805 6880 2839
rect 6828 2796 6880 2805
rect 17408 2796 17460 2848
rect 19892 2796 19944 2848
rect 19984 2796 20036 2848
rect 21180 2796 21232 2848
rect 21272 2796 21324 2848
rect 26884 2796 26936 2848
rect 27620 2796 27672 2848
rect 30932 2796 30984 2848
rect 32864 2796 32916 2848
rect 44364 3068 44416 3120
rect 45376 3111 45428 3120
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 47768 3043 47820 3052
rect 47768 3009 47777 3043
rect 47777 3009 47811 3043
rect 47811 3009 47820 3043
rect 47768 3000 47820 3009
rect 45652 2932 45704 2984
rect 47676 2932 47728 2984
rect 40132 2796 40184 2848
rect 44364 2796 44416 2848
rect 47860 2839 47912 2848
rect 47860 2805 47869 2839
rect 47869 2805 47903 2839
rect 47903 2805 47912 2839
rect 47860 2796 47912 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3240 2592 3292 2644
rect 10416 2592 10468 2644
rect 15476 2592 15528 2644
rect 16948 2592 17000 2644
rect 18512 2592 18564 2644
rect 19892 2592 19944 2644
rect 21272 2592 21324 2644
rect 23480 2592 23532 2644
rect 23848 2592 23900 2644
rect 28632 2635 28684 2644
rect 2780 2524 2832 2576
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2872 2499 2924 2508
rect 2872 2465 2881 2499
rect 2881 2465 2915 2499
rect 2915 2465 2924 2499
rect 2872 2456 2924 2465
rect 15200 2524 15252 2576
rect 22652 2524 22704 2576
rect 24400 2524 24452 2576
rect 6828 2456 6880 2508
rect 6920 2456 6972 2508
rect 2596 2320 2648 2372
rect 5172 2388 5224 2440
rect 15476 2388 15528 2440
rect 21640 2456 21692 2508
rect 25412 2524 25464 2576
rect 28632 2601 28641 2635
rect 28641 2601 28675 2635
rect 28675 2601 28684 2635
rect 28632 2592 28684 2601
rect 38292 2635 38344 2644
rect 38292 2601 38301 2635
rect 38301 2601 38335 2635
rect 38335 2601 38344 2635
rect 38292 2592 38344 2601
rect 39120 2592 39172 2644
rect 39304 2592 39356 2644
rect 43720 2592 43772 2644
rect 44364 2635 44416 2644
rect 44364 2601 44373 2635
rect 44373 2601 44407 2635
rect 44407 2601 44416 2635
rect 44364 2592 44416 2601
rect 24676 2499 24728 2508
rect 24676 2465 24685 2499
rect 24685 2465 24719 2499
rect 24719 2465 24728 2499
rect 24676 2456 24728 2465
rect 7472 2320 7524 2372
rect 8392 2320 8444 2372
rect 16120 2320 16172 2372
rect 19064 2388 19116 2440
rect 23020 2431 23072 2440
rect 23020 2397 23029 2431
rect 23029 2397 23063 2431
rect 23063 2397 23072 2431
rect 23020 2388 23072 2397
rect 23664 2431 23716 2440
rect 23664 2397 23673 2431
rect 23673 2397 23707 2431
rect 23707 2397 23716 2431
rect 23664 2388 23716 2397
rect 20628 2320 20680 2372
rect 25688 2499 25740 2508
rect 25688 2465 25697 2499
rect 25697 2465 25731 2499
rect 25731 2465 25740 2499
rect 25688 2456 25740 2465
rect 27160 2456 27212 2508
rect 30012 2499 30064 2508
rect 25596 2388 25648 2440
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 9680 2252 9732 2261
rect 21916 2252 21968 2304
rect 24492 2252 24544 2304
rect 26424 2388 26476 2440
rect 29644 2388 29696 2440
rect 30012 2465 30021 2499
rect 30021 2465 30055 2499
rect 30055 2465 30064 2499
rect 30012 2456 30064 2465
rect 41512 2456 41564 2508
rect 46112 2456 46164 2508
rect 47032 2456 47084 2508
rect 35440 2388 35492 2440
rect 38016 2388 38068 2440
rect 40040 2388 40092 2440
rect 41236 2388 41288 2440
rect 43812 2388 43864 2440
rect 44180 2431 44232 2440
rect 44180 2397 44189 2431
rect 44189 2397 44223 2431
rect 44223 2397 44232 2431
rect 44180 2388 44232 2397
rect 46296 2388 46348 2440
rect 28356 2320 28408 2372
rect 39304 2320 39356 2372
rect 40592 2320 40644 2372
rect 31576 2252 31628 2304
rect 46388 2320 46440 2372
rect 47952 2320 48004 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 9680 2048 9732 2100
rect 25044 2048 25096 2100
rect 44180 484 44232 536
rect 46848 484 46900 536
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4844 49314
rect 4498 49200 4610 49286
rect 32 20874 60 49200
rect 1398 47696 1454 47705
rect 1398 47631 1454 47640
rect 1412 46578 1440 47631
rect 1964 47054 1992 49200
rect 2608 47054 2636 49200
rect 3252 47054 3280 49200
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2596 47048 2648 47054
rect 2596 46990 2648 46996
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3422 47016 3478 47025
rect 3422 46951 3478 46960
rect 2136 46912 2188 46918
rect 2136 46854 2188 46860
rect 2872 46912 2924 46918
rect 2872 46854 2924 46860
rect 1400 46572 1452 46578
rect 1400 46514 1452 46520
rect 1676 46368 1728 46374
rect 1676 46310 1728 46316
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1584 43104 1636 43110
rect 1584 43046 1636 43052
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1596 42158 1624 43046
rect 1584 42152 1636 42158
rect 1584 42094 1636 42100
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1584 41540 1636 41546
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1688 35894 1716 46310
rect 2148 43246 2176 46854
rect 2884 46646 2912 46854
rect 2872 46640 2924 46646
rect 2872 46582 2924 46588
rect 2320 46368 2372 46374
rect 2320 46310 2372 46316
rect 2778 46336 2834 46345
rect 2332 46034 2360 46310
rect 2778 46271 2834 46280
rect 2792 46034 2820 46271
rect 2320 46028 2372 46034
rect 2320 45970 2372 45976
rect 2780 46028 2832 46034
rect 2780 45970 2832 45976
rect 2320 45892 2372 45898
rect 2320 45834 2372 45840
rect 2332 45626 2360 45834
rect 2320 45620 2372 45626
rect 2320 45562 2372 45568
rect 2320 45484 2372 45490
rect 2320 45426 2372 45432
rect 2136 43240 2188 43246
rect 2136 43182 2188 43188
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 2044 40452 2096 40458
rect 2044 40394 2096 40400
rect 1872 40225 1900 40394
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 2056 37398 2084 40394
rect 2044 37392 2096 37398
rect 2044 37334 2096 37340
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1780 36786 1808 37198
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 2228 36712 2280 36718
rect 2228 36654 2280 36660
rect 2240 36378 2268 36654
rect 2228 36372 2280 36378
rect 2228 36314 2280 36320
rect 2136 36168 2188 36174
rect 2136 36110 2188 36116
rect 1688 35866 1808 35894
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1492 35488 1544 35494
rect 1596 35465 1624 35634
rect 1492 35430 1544 35436
rect 1582 35456 1638 35465
rect 1308 33992 1360 33998
rect 1308 33934 1360 33940
rect 1320 32745 1348 33934
rect 1400 33448 1452 33454
rect 1398 33416 1400 33425
rect 1452 33416 1454 33425
rect 1398 33351 1454 33360
rect 1504 33046 1532 35430
rect 1582 35391 1638 35400
rect 1584 33856 1636 33862
rect 1584 33798 1636 33804
rect 1492 33040 1544 33046
rect 1492 32982 1544 32988
rect 1596 32978 1624 33798
rect 1676 33448 1728 33454
rect 1676 33390 1728 33396
rect 1584 32972 1636 32978
rect 1584 32914 1636 32920
rect 1306 32736 1362 32745
rect 1306 32671 1362 32680
rect 1688 32502 1716 33390
rect 1676 32496 1728 32502
rect 1676 32438 1728 32444
rect 1400 32224 1452 32230
rect 1400 32166 1452 32172
rect 1412 31890 1440 32166
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1596 31482 1624 31690
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 1780 27130 1808 35866
rect 1858 32056 1914 32065
rect 1858 31991 1914 32000
rect 1872 31890 1900 31991
rect 1860 31884 1912 31890
rect 1860 31826 1912 31832
rect 1768 27124 1820 27130
rect 1768 27066 1820 27072
rect 1400 25288 1452 25294
rect 1398 25256 1400 25265
rect 1452 25256 1454 25265
rect 1398 25191 1454 25200
rect 1676 25220 1728 25226
rect 1676 25162 1728 25168
rect 20 20868 72 20874
rect 20 20810 72 20816
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1688 6730 1716 25162
rect 1952 24268 2004 24274
rect 1952 24210 2004 24216
rect 1964 23866 1992 24210
rect 1952 23860 2004 23866
rect 1952 23802 2004 23808
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 23225 1900 23666
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2148 18766 2176 36110
rect 2332 31346 2360 45426
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36718 2820 36751
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 3240 32836 3292 32842
rect 3240 32778 3292 32784
rect 3252 32366 3280 32778
rect 2412 32360 2464 32366
rect 2412 32302 2464 32308
rect 3240 32360 3292 32366
rect 3240 32302 3292 32308
rect 2320 31340 2372 31346
rect 2320 31282 2372 31288
rect 2424 19514 2452 32302
rect 3252 20330 3280 32302
rect 3436 23866 3464 46951
rect 3896 46102 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4816 47054 4844 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49200 7186 50000
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49314 13626 50000
rect 13514 49286 13768 49314
rect 13514 49200 13626 49286
rect 5828 47054 5856 49200
rect 7116 47054 7144 49200
rect 4804 47048 4856 47054
rect 4804 46990 4856 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7104 47048 7156 47054
rect 7104 46990 7156 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 7840 46980 7892 46986
rect 7840 46922 7892 46928
rect 3884 46096 3936 46102
rect 3884 46038 3936 46044
rect 3514 44976 3570 44985
rect 3514 44911 3570 44920
rect 3528 44334 3556 44911
rect 3516 44328 3568 44334
rect 3516 44270 3568 44276
rect 3698 43616 3754 43625
rect 3698 43551 3754 43560
rect 3514 39536 3570 39545
rect 3514 39471 3570 39480
rect 3528 24682 3556 39471
rect 3712 28626 3740 43551
rect 3882 31376 3938 31385
rect 3882 31311 3938 31320
rect 3700 28620 3752 28626
rect 3700 28562 3752 28568
rect 3516 24676 3568 24682
rect 3516 24618 3568 24624
rect 3896 24342 3924 31311
rect 3974 28656 4030 28665
rect 3974 28591 4030 28600
rect 3988 27878 4016 28591
rect 3976 27872 4028 27878
rect 3976 27814 4028 27820
rect 3884 24336 3936 24342
rect 3884 24278 3936 24284
rect 3424 23860 3476 23866
rect 3424 23802 3476 23808
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3240 20324 3292 20330
rect 3240 20266 3292 20272
rect 3988 19825 4016 20538
rect 3974 19816 4030 19825
rect 3974 19751 4030 19760
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2148 18358 2176 18702
rect 3330 18456 3386 18465
rect 3330 18391 3386 18400
rect 2136 18352 2188 18358
rect 2136 18294 2188 18300
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1872 17785 1900 18226
rect 1858 17776 1914 17785
rect 1858 17711 1914 17720
rect 3344 16794 3372 18391
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3988 17105 4016 17682
rect 3974 17096 4030 17105
rect 3974 17031 4030 17040
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1872 16425 1900 16594
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 2148 16250 2176 16458
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 2056 4146 2084 16050
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1320 800 1348 3402
rect 1596 2514 1624 3878
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 3058 1808 3538
rect 2700 3534 2728 14350
rect 3976 13728 4028 13734
rect 3974 13696 3976 13705
rect 4028 13696 4030 13705
rect 3974 13631 4030 13640
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10305 2820 10950
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7585 3464 8230
rect 3422 7576 3478 7585
rect 3422 7511 3478 7520
rect 3528 7426 3556 10474
rect 3436 7398 3556 7426
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1964 3126 1992 3334
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2792 2582 2820 3878
rect 3436 3505 3464 7398
rect 4080 6914 4108 46922
rect 4896 46912 4948 46918
rect 4896 46854 4948 46860
rect 6920 46912 6972 46918
rect 6920 46854 6972 46860
rect 4620 46368 4672 46374
rect 4620 46310 4672 46316
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4632 46034 4660 46310
rect 4620 46028 4672 46034
rect 4620 45970 4672 45976
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4632 13734 4660 21626
rect 4908 18970 4936 46854
rect 5080 45892 5132 45898
rect 5080 45834 5132 45840
rect 5092 45626 5120 45834
rect 5080 45620 5132 45626
rect 5080 45562 5132 45568
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4908 11014 4936 18770
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3514 6896 3570 6905
rect 3514 6831 3516 6840
rect 3568 6831 3570 6840
rect 3988 6886 4108 6914
rect 3516 6802 3568 6808
rect 3988 4049 4016 6886
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 6656 4146 6684 18294
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 3974 4040 4030 4049
rect 3974 3975 4030 3984
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 6748 3602 6776 3878
rect 6932 3738 6960 46854
rect 7852 29238 7880 46922
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9496 46980 9548 46986
rect 9496 46922 9548 46928
rect 8312 45526 8432 45554
rect 8312 30802 8340 45526
rect 9508 37466 9536 46922
rect 10416 46368 10468 46374
rect 10416 46310 10468 46316
rect 10428 46034 10456 46310
rect 10980 46034 11008 49200
rect 11624 47122 11652 49200
rect 11612 47116 11664 47122
rect 11612 47058 11664 47064
rect 11980 47048 12032 47054
rect 11980 46990 12032 46996
rect 10416 46028 10468 46034
rect 10416 45970 10468 45976
rect 10968 46028 11020 46034
rect 10968 45970 11020 45976
rect 10600 45892 10652 45898
rect 10600 45834 10652 45840
rect 10612 45626 10640 45834
rect 10600 45620 10652 45626
rect 10600 45562 10652 45568
rect 11992 38282 12020 46990
rect 12268 46578 12296 49200
rect 12912 47054 12940 49200
rect 13740 47138 13768 49286
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49314 16202 50000
rect 16090 49286 16528 49314
rect 16090 49200 16202 49286
rect 14200 47954 14228 49200
rect 14200 47926 14320 47954
rect 13740 47110 13860 47138
rect 13832 47054 13860 47110
rect 12900 47048 12952 47054
rect 12900 46990 12952 46996
rect 13820 47048 13872 47054
rect 13820 46990 13872 46996
rect 12256 46572 12308 46578
rect 12256 46514 12308 46520
rect 14292 46510 14320 47926
rect 14648 46980 14700 46986
rect 14648 46922 14700 46928
rect 13544 46504 13596 46510
rect 13544 46446 13596 46452
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 12532 46368 12584 46374
rect 12532 46310 12584 46316
rect 11980 38276 12032 38282
rect 11980 38218 12032 38224
rect 9496 37460 9548 37466
rect 9496 37402 9548 37408
rect 12544 32978 12572 46310
rect 13556 46170 13584 46446
rect 14200 46170 14228 46446
rect 13544 46164 13596 46170
rect 13544 46106 13596 46112
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 14096 45960 14148 45966
rect 14096 45902 14148 45908
rect 14108 41138 14136 45902
rect 14096 41132 14148 41138
rect 14096 41074 14148 41080
rect 12532 32972 12584 32978
rect 12532 32914 12584 32920
rect 14660 30802 14688 46922
rect 15488 45554 15516 49200
rect 16500 47054 16528 49286
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49200 27150 50000
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49314 31014 50000
rect 30760 49286 31014 49314
rect 17420 47410 17448 49200
rect 16592 47382 17448 47410
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 15488 45526 16160 45554
rect 15660 36168 15712 36174
rect 15660 36110 15712 36116
rect 15672 33998 15700 36110
rect 15660 33992 15712 33998
rect 15660 33934 15712 33940
rect 15672 32434 15700 33934
rect 16028 33924 16080 33930
rect 16028 33866 16080 33872
rect 16040 33658 16068 33866
rect 16028 33652 16080 33658
rect 16028 33594 16080 33600
rect 15660 32428 15712 32434
rect 15660 32370 15712 32376
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 14648 30796 14700 30802
rect 14648 30738 14700 30744
rect 14004 30728 14056 30734
rect 14004 30670 14056 30676
rect 13636 30252 13688 30258
rect 13636 30194 13688 30200
rect 13648 29646 13676 30194
rect 13912 30184 13964 30190
rect 13912 30126 13964 30132
rect 13636 29640 13688 29646
rect 13636 29582 13688 29588
rect 7840 29232 7892 29238
rect 7840 29174 7892 29180
rect 13924 29170 13952 30126
rect 10876 29164 10928 29170
rect 10876 29106 10928 29112
rect 13544 29164 13596 29170
rect 13544 29106 13596 29112
rect 13912 29164 13964 29170
rect 13912 29106 13964 29112
rect 10048 28484 10100 28490
rect 10048 28426 10100 28432
rect 9956 28416 10008 28422
rect 9956 28358 10008 28364
rect 9772 27532 9824 27538
rect 9772 27474 9824 27480
rect 9128 27328 9180 27334
rect 9128 27270 9180 27276
rect 9140 26994 9168 27270
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9416 26586 9444 26862
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 9784 24818 9812 27474
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9876 24954 9904 25230
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9588 24200 9640 24206
rect 9784 24188 9812 24754
rect 9640 24160 9812 24188
rect 9588 24142 9640 24148
rect 8208 24064 8260 24070
rect 8208 24006 8260 24012
rect 8220 23730 8248 24006
rect 8208 23724 8260 23730
rect 8208 23666 8260 23672
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 8496 23322 8524 23598
rect 9692 23594 9720 24160
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9784 23798 9812 24006
rect 9772 23792 9824 23798
rect 9772 23734 9824 23740
rect 9968 23662 9996 28358
rect 10060 28218 10088 28426
rect 10048 28212 10100 28218
rect 10048 28154 10100 28160
rect 10888 28082 10916 29106
rect 12072 28552 12124 28558
rect 12072 28494 12124 28500
rect 13084 28552 13136 28558
rect 13084 28494 13136 28500
rect 13176 28552 13228 28558
rect 13176 28494 13228 28500
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11808 28150 11836 28358
rect 11796 28144 11848 28150
rect 11796 28086 11848 28092
rect 10876 28076 10928 28082
rect 10876 28018 10928 28024
rect 10888 27538 10916 28018
rect 12084 27674 12112 28494
rect 12072 27668 12124 27674
rect 12072 27610 12124 27616
rect 13096 27606 13124 28494
rect 13188 27674 13216 28494
rect 13268 27872 13320 27878
rect 13268 27814 13320 27820
rect 13176 27668 13228 27674
rect 13176 27610 13228 27616
rect 13084 27600 13136 27606
rect 13084 27542 13136 27548
rect 10876 27532 10928 27538
rect 10876 27474 10928 27480
rect 10600 27464 10652 27470
rect 10600 27406 10652 27412
rect 10416 27056 10468 27062
rect 10416 26998 10468 27004
rect 10428 26042 10456 26998
rect 10612 26858 10640 27406
rect 11980 27396 12032 27402
rect 11980 27338 12032 27344
rect 10876 27328 10928 27334
rect 10876 27270 10928 27276
rect 10600 26852 10652 26858
rect 10600 26794 10652 26800
rect 10612 26450 10640 26794
rect 10888 26790 10916 27270
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10600 26444 10652 26450
rect 10600 26386 10652 26392
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 10152 24954 10180 25162
rect 10140 24948 10192 24954
rect 10140 24890 10192 24896
rect 10244 24750 10272 25842
rect 10612 24818 10640 26386
rect 10888 26382 10916 26726
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 11428 25220 11480 25226
rect 11428 25162 11480 25168
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 9956 23656 10008 23662
rect 9956 23598 10008 23604
rect 9680 23588 9732 23594
rect 9680 23530 9732 23536
rect 9968 23322 9996 23598
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9784 22778 9812 23054
rect 9968 23050 9996 23258
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 10048 22976 10100 22982
rect 10152 22964 10180 24142
rect 10244 24138 10272 24686
rect 10428 24410 10456 24754
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 11072 24206 11100 25094
rect 11440 24750 11468 25162
rect 11704 24948 11756 24954
rect 11704 24890 11756 24896
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 10232 24132 10284 24138
rect 10232 24074 10284 24080
rect 10244 24018 10272 24074
rect 10508 24064 10560 24070
rect 10244 23990 10456 24018
rect 10508 24006 10560 24012
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 10100 22936 10180 22964
rect 10048 22918 10100 22924
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9496 22500 9548 22506
rect 9496 22442 9548 22448
rect 9508 22234 9536 22442
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9692 21978 9720 22646
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9784 22098 9812 22374
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9876 21978 9904 22374
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 9692 21962 9812 21978
rect 9692 21956 9824 21962
rect 9692 21950 9772 21956
rect 9876 21950 9996 21978
rect 9772 21898 9824 21904
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8220 21622 8248 21830
rect 8208 21616 8260 21622
rect 8208 21558 8260 21564
rect 9784 21486 9812 21898
rect 9968 21894 9996 21950
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 10060 21690 10088 22034
rect 10152 21962 10180 22936
rect 10244 22710 10272 23258
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10232 22704 10284 22710
rect 10232 22646 10284 22652
rect 10336 22438 10364 22918
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10140 21616 10192 21622
rect 10140 21558 10192 21564
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9140 21146 9168 21422
rect 10152 21146 10180 21558
rect 10428 21350 10456 23990
rect 10520 23526 10548 24006
rect 11072 23798 11100 24142
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 11060 23792 11112 23798
rect 11060 23734 11112 23740
rect 10600 23588 10652 23594
rect 10600 23530 10652 23536
rect 10508 23520 10560 23526
rect 10508 23462 10560 23468
rect 10520 23322 10548 23462
rect 10508 23316 10560 23322
rect 10508 23258 10560 23264
rect 10612 23186 10640 23530
rect 11256 23322 11284 24074
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 10692 23248 10744 23254
rect 10692 23190 10744 23196
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10704 22710 10732 23190
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10704 22030 10732 22646
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 10428 20942 10456 21286
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 9416 20534 9444 20878
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 10428 20466 10456 20878
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 8944 20256 8996 20262
rect 8944 20198 8996 20204
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 8956 19922 8984 20198
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 9968 19786 9996 20198
rect 10612 20058 10640 21830
rect 11072 20942 11100 23054
rect 11716 22030 11744 24890
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11900 22098 11928 22374
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 9956 19780 10008 19786
rect 9956 19722 10008 19728
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7576 18426 7604 19110
rect 8864 18766 8892 19314
rect 9232 19310 9260 19722
rect 10612 19378 10640 19994
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 8220 17202 8248 18702
rect 11072 17202 11100 20878
rect 11440 19854 11468 21898
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11532 19922 11560 20878
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11256 19446 11284 19654
rect 11244 19440 11296 19446
rect 11244 19382 11296 19388
rect 11348 19378 11376 19654
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11440 19242 11468 19790
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11716 17338 11744 17546
rect 11992 17542 12020 27338
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12992 26988 13044 26994
rect 13096 26976 13124 27542
rect 13280 27470 13308 27814
rect 13268 27464 13320 27470
rect 13268 27406 13320 27412
rect 13556 27402 13584 29106
rect 13820 28960 13872 28966
rect 13820 28902 13872 28908
rect 13832 28626 13860 28902
rect 13820 28620 13872 28626
rect 13820 28562 13872 28568
rect 13924 27402 13952 29106
rect 14016 27606 14044 30670
rect 14280 30660 14332 30666
rect 14280 30602 14332 30608
rect 14292 30326 14320 30602
rect 16132 30326 16160 45526
rect 16304 37800 16356 37806
rect 16304 37742 16356 37748
rect 16316 36174 16344 37742
rect 16304 36168 16356 36174
rect 16304 36110 16356 36116
rect 14280 30320 14332 30326
rect 14280 30262 14332 30268
rect 16120 30320 16172 30326
rect 16120 30262 16172 30268
rect 14648 30184 14700 30190
rect 14648 30126 14700 30132
rect 14660 29850 14688 30126
rect 14648 29844 14700 29850
rect 14648 29786 14700 29792
rect 15844 29096 15896 29102
rect 15844 29038 15896 29044
rect 14096 29028 14148 29034
rect 14096 28970 14148 28976
rect 14108 28626 14136 28970
rect 15856 28762 15884 29038
rect 16592 29034 16620 47382
rect 17776 47184 17828 47190
rect 17776 47126 17828 47132
rect 16672 45892 16724 45898
rect 16672 45834 16724 45840
rect 16684 45490 16712 45834
rect 16672 45484 16724 45490
rect 16672 45426 16724 45432
rect 16684 39370 16712 45426
rect 16672 39364 16724 39370
rect 16672 39306 16724 39312
rect 17592 39364 17644 39370
rect 17592 39306 17644 39312
rect 17132 38208 17184 38214
rect 17132 38150 17184 38156
rect 17144 37942 17172 38150
rect 17132 37936 17184 37942
rect 17132 37878 17184 37884
rect 17316 36100 17368 36106
rect 17316 36042 17368 36048
rect 17328 35834 17356 36042
rect 17316 35828 17368 35834
rect 17316 35770 17368 35776
rect 16672 35692 16724 35698
rect 16672 35634 16724 35640
rect 16684 33522 16712 35634
rect 17500 34672 17552 34678
rect 17500 34614 17552 34620
rect 17132 34604 17184 34610
rect 17132 34546 17184 34552
rect 16948 34400 17000 34406
rect 16948 34342 17000 34348
rect 16960 34066 16988 34342
rect 16948 34060 17000 34066
rect 16948 34002 17000 34008
rect 17144 33658 17172 34546
rect 17132 33652 17184 33658
rect 17132 33594 17184 33600
rect 16672 33516 16724 33522
rect 16672 33458 16724 33464
rect 17316 33516 17368 33522
rect 17368 33476 17448 33504
rect 17316 33458 17368 33464
rect 16684 33046 16712 33458
rect 17040 33448 17092 33454
rect 17040 33390 17092 33396
rect 16672 33040 16724 33046
rect 16672 32982 16724 32988
rect 16856 32768 16908 32774
rect 16856 32710 16908 32716
rect 16868 32502 16896 32710
rect 16856 32496 16908 32502
rect 16856 32438 16908 32444
rect 16948 32360 17000 32366
rect 16948 32302 17000 32308
rect 16960 32026 16988 32302
rect 16948 32020 17000 32026
rect 16948 31962 17000 31968
rect 16856 31680 16908 31686
rect 16856 31622 16908 31628
rect 16868 31414 16896 31622
rect 16856 31408 16908 31414
rect 16856 31350 16908 31356
rect 16856 29096 16908 29102
rect 16856 29038 16908 29044
rect 16580 29028 16632 29034
rect 16580 28970 16632 28976
rect 15844 28756 15896 28762
rect 15844 28698 15896 28704
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 14832 28484 14884 28490
rect 14832 28426 14884 28432
rect 14844 28218 14872 28426
rect 14832 28212 14884 28218
rect 14832 28154 14884 28160
rect 14096 28076 14148 28082
rect 14096 28018 14148 28024
rect 14004 27600 14056 27606
rect 14004 27542 14056 27548
rect 13544 27396 13596 27402
rect 13544 27338 13596 27344
rect 13912 27396 13964 27402
rect 13912 27338 13964 27344
rect 13556 26994 13584 27338
rect 13044 26948 13124 26976
rect 13544 26988 13596 26994
rect 12992 26930 13044 26936
rect 13820 26988 13872 26994
rect 13596 26948 13820 26976
rect 13544 26930 13596 26936
rect 13820 26930 13872 26936
rect 12072 26784 12124 26790
rect 12072 26726 12124 26732
rect 12084 26450 12112 26726
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12728 26042 12756 26182
rect 12716 26036 12768 26042
rect 12716 25978 12768 25984
rect 12820 25362 12848 26930
rect 14016 26926 14044 27542
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 14016 26586 14044 26862
rect 14004 26580 14056 26586
rect 14004 26522 14056 26528
rect 14108 26382 14136 28018
rect 15856 27674 15884 28698
rect 16868 28218 16896 29038
rect 16856 28212 16908 28218
rect 16856 28154 16908 28160
rect 16028 28008 16080 28014
rect 16028 27950 16080 27956
rect 16672 28008 16724 28014
rect 16672 27950 16724 27956
rect 16856 28008 16908 28014
rect 16856 27950 16908 27956
rect 15844 27668 15896 27674
rect 15844 27610 15896 27616
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 14648 27328 14700 27334
rect 14648 27270 14700 27276
rect 14660 27062 14688 27270
rect 14648 27056 14700 27062
rect 14648 26998 14700 27004
rect 15200 27056 15252 27062
rect 15200 26998 15252 27004
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12360 24954 12388 25230
rect 12992 25152 13044 25158
rect 12992 25094 13044 25100
rect 12348 24948 12400 24954
rect 12348 24890 12400 24896
rect 13004 24886 13032 25094
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 12532 24676 12584 24682
rect 12532 24618 12584 24624
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12452 24274 12480 24550
rect 12544 24274 12572 24618
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 12716 24200 12768 24206
rect 12716 24142 12768 24148
rect 12728 22778 12756 24142
rect 13464 24138 13492 25842
rect 13544 24880 13596 24886
rect 14108 24834 14136 26318
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 13544 24822 13596 24828
rect 13556 24342 13584 24822
rect 14016 24806 14136 24834
rect 13544 24336 13596 24342
rect 13544 24278 13596 24284
rect 14016 24206 14044 24806
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 14108 24342 14136 24686
rect 14096 24336 14148 24342
rect 14096 24278 14148 24284
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 13452 24132 13504 24138
rect 13452 24074 13504 24080
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 13004 23050 13032 23666
rect 13464 23526 13492 24074
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 13452 23520 13504 23526
rect 13504 23468 13584 23474
rect 13452 23462 13584 23468
rect 13464 23446 13584 23462
rect 12992 23044 13044 23050
rect 12992 22986 13044 22992
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 13004 20466 13032 22986
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 13372 22098 13400 22714
rect 13452 22568 13504 22574
rect 13452 22510 13504 22516
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13464 21962 13492 22510
rect 13556 22030 13584 23446
rect 14568 23322 14596 23734
rect 15120 23594 15148 25774
rect 15212 24818 15240 26998
rect 15660 26852 15712 26858
rect 15660 26794 15712 26800
rect 15672 26382 15700 26794
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15764 26042 15792 27406
rect 15936 27328 15988 27334
rect 15936 27270 15988 27276
rect 15948 26994 15976 27270
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 16040 26874 16068 27950
rect 16120 27056 16172 27062
rect 16120 26998 16172 27004
rect 15948 26846 16068 26874
rect 15752 26036 15804 26042
rect 15752 25978 15804 25984
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15580 25770 15608 25842
rect 15568 25764 15620 25770
rect 15568 25706 15620 25712
rect 15580 25378 15608 25706
rect 15396 25350 15608 25378
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15212 24138 15240 24754
rect 15304 24342 15332 24890
rect 15292 24336 15344 24342
rect 15292 24278 15344 24284
rect 15200 24132 15252 24138
rect 15200 24074 15252 24080
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15108 23588 15160 23594
rect 15108 23530 15160 23536
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 14108 22234 14136 22510
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13452 21956 13504 21962
rect 13452 21898 13504 21904
rect 13464 21554 13492 21898
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13372 20942 13400 21286
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 13096 20262 13124 20470
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13096 19718 13124 20198
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12544 18970 12572 19382
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 13096 18766 13124 19654
rect 13188 19514 13216 19926
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 13372 18834 13400 20878
rect 14188 20528 14240 20534
rect 14188 20470 14240 20476
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 13924 20058 13952 20334
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 14200 19990 14228 20470
rect 14568 20058 14596 23258
rect 15304 23050 15332 23666
rect 15292 23044 15344 23050
rect 15292 22986 15344 22992
rect 15396 22982 15424 25350
rect 15476 25288 15528 25294
rect 15476 25230 15528 25236
rect 15488 24886 15516 25230
rect 15568 25152 15620 25158
rect 15568 25094 15620 25100
rect 15660 25152 15712 25158
rect 15660 25094 15712 25100
rect 15476 24880 15528 24886
rect 15476 24822 15528 24828
rect 15580 24274 15608 25094
rect 15672 24886 15700 25094
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15488 23662 15516 24006
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 14648 20800 14700 20806
rect 14648 20742 14700 20748
rect 14660 20534 14688 20742
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14188 19984 14240 19990
rect 14188 19926 14240 19932
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13740 19310 13768 19722
rect 13924 19446 13952 19790
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 14108 19378 14136 19654
rect 14200 19378 14228 19722
rect 14280 19440 14332 19446
rect 14280 19382 14332 19388
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 18290 12940 18566
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 13372 17202 13400 18770
rect 14108 18698 14136 19314
rect 14200 18970 14228 19314
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 13924 17338 13952 18294
rect 14200 17542 14228 18906
rect 14292 18630 14320 19382
rect 14476 18970 14504 19858
rect 15212 18970 15240 22918
rect 15384 22704 15436 22710
rect 15384 22646 15436 22652
rect 15396 22098 15424 22646
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14280 18624 14332 18630
rect 14332 18584 14412 18612
rect 14280 18566 14332 18572
rect 14384 17678 14412 18584
rect 14476 18358 14504 18906
rect 15212 18834 15240 18906
rect 15488 18850 15516 23598
rect 15672 23118 15700 24822
rect 15764 24206 15792 25978
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 15856 24070 15884 25230
rect 15948 24138 15976 26846
rect 16028 26444 16080 26450
rect 16028 26386 16080 26392
rect 16040 25974 16068 26386
rect 16028 25968 16080 25974
rect 16028 25910 16080 25916
rect 15936 24132 15988 24138
rect 15936 24074 15988 24080
rect 15844 24064 15896 24070
rect 15844 24006 15896 24012
rect 15856 23254 15884 24006
rect 15844 23248 15896 23254
rect 15844 23190 15896 23196
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15764 22778 15792 23122
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 15948 22506 15976 24074
rect 16132 23730 16160 26998
rect 16580 26988 16632 26994
rect 16580 26930 16632 26936
rect 16396 26784 16448 26790
rect 16396 26726 16448 26732
rect 16408 26450 16436 26726
rect 16592 26586 16620 26930
rect 16580 26580 16632 26586
rect 16580 26522 16632 26528
rect 16684 26466 16712 27950
rect 16868 27674 16896 27950
rect 16856 27668 16908 27674
rect 16856 27610 16908 27616
rect 16764 26852 16816 26858
rect 16764 26794 16816 26800
rect 16396 26444 16448 26450
rect 16396 26386 16448 26392
rect 16592 26438 16712 26466
rect 16592 25974 16620 26438
rect 16776 26330 16804 26794
rect 16672 26308 16724 26314
rect 16776 26302 16896 26330
rect 16672 26250 16724 26256
rect 16580 25968 16632 25974
rect 16580 25910 16632 25916
rect 16684 25498 16712 26250
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16776 26042 16804 26182
rect 16764 26036 16816 26042
rect 16764 25978 16816 25984
rect 16672 25492 16724 25498
rect 16672 25434 16724 25440
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 16592 24274 16620 25230
rect 16776 24954 16804 25978
rect 16764 24948 16816 24954
rect 16764 24890 16816 24896
rect 16672 24744 16724 24750
rect 16672 24686 16724 24692
rect 16580 24268 16632 24274
rect 16580 24210 16632 24216
rect 16592 23730 16620 24210
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16580 23724 16632 23730
rect 16580 23666 16632 23672
rect 16684 23594 16712 24686
rect 16776 24070 16804 24890
rect 16868 24206 16896 26302
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 16960 24342 16988 24686
rect 16948 24336 17000 24342
rect 16948 24278 17000 24284
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 16672 23588 16724 23594
rect 16672 23530 16724 23536
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 15936 22500 15988 22506
rect 15936 22442 15988 22448
rect 15948 21554 15976 22442
rect 16132 22438 16160 23054
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15856 21010 15884 21286
rect 15948 21146 15976 21490
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15672 20602 15700 20878
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15672 19854 15700 20538
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15396 18822 15516 18850
rect 15396 18766 15424 18822
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14660 18086 14688 18634
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14660 17746 14688 18022
rect 15120 17882 15148 18226
rect 15396 18086 15424 18702
rect 15672 18290 15700 19654
rect 16132 18290 16160 22374
rect 16684 21622 16712 22578
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 16868 21622 16896 22374
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16960 21690 16988 21898
rect 16948 21684 17000 21690
rect 16948 21626 17000 21632
rect 16672 21616 16724 21622
rect 16672 21558 16724 21564
rect 16856 21616 16908 21622
rect 16856 21558 16908 21564
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 8220 17066 8248 17138
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 3422 3496 3478 3505
rect 3422 3431 3478 3440
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2608 800 2636 2314
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 2884 785 2912 2450
rect 3252 1465 3280 2586
rect 3238 1456 3294 1465
rect 3238 1391 3294 1400
rect 3896 800 3924 3130
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 6840 2514 6868 2790
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 5172 2440 5224 2446
rect 3974 2408 4030 2417
rect 5172 2382 5224 2388
rect 3974 2343 4030 2352
rect 3988 2310 4016 2343
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 5184 800 5212 2382
rect 6932 1442 6960 2450
rect 6472 1414 6960 1442
rect 6472 800 6500 1414
rect 7116 800 7144 3538
rect 7484 2378 7512 3878
rect 7668 3058 7696 4558
rect 8220 4146 8248 17002
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 7852 3126 7880 3878
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 7760 800 7788 2858
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8404 800 8432 2314
rect 9048 800 9076 3606
rect 9232 3602 9260 3878
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9968 3058 9996 3606
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10060 3126 10088 3402
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10428 2650 10456 17070
rect 11624 16998 11652 17138
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 14200 16250 14228 17478
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12728 15638 12756 15846
rect 13556 15706 13584 15982
rect 14384 15910 14412 17614
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15212 17338 15240 17546
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15672 17202 15700 18226
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14292 14414 14320 15438
rect 14384 14414 14412 15846
rect 14844 15502 14872 17138
rect 15672 16998 15700 17138
rect 16592 17134 16620 19382
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15764 16658 15792 16934
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15120 16250 15148 16526
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14936 15706 14964 16050
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14844 15026 14872 15438
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 13938 14320 14214
rect 15028 14006 15056 14758
rect 16316 14414 16344 15302
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 15212 13734 15240 14214
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12452 8294 12480 13466
rect 15856 13394 15884 14214
rect 16040 14074 16068 14350
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 16040 13462 16068 14010
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 16592 11830 16620 17070
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11532 3058 11560 3878
rect 14108 3534 14136 4014
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11716 3126 11744 3334
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 13832 3058 13860 3470
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 14016 3126 14044 3334
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 2106 9720 2246
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 10980 800 11008 2926
rect 14108 2922 14136 3470
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14096 2916 14148 2922
rect 14096 2858 14148 2864
rect 14200 800 14228 2926
rect 14844 800 14872 11222
rect 16868 11218 16896 13194
rect 17052 12434 17080 33390
rect 17316 31884 17368 31890
rect 17316 31826 17368 31832
rect 17328 31793 17356 31826
rect 17314 31784 17370 31793
rect 17314 31719 17370 31728
rect 17420 30394 17448 33476
rect 17512 33114 17540 34614
rect 17500 33108 17552 33114
rect 17500 33050 17552 33056
rect 17512 31822 17540 33050
rect 17500 31816 17552 31822
rect 17500 31758 17552 31764
rect 17408 30388 17460 30394
rect 17408 30330 17460 30336
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17512 25498 17540 26318
rect 17500 25492 17552 25498
rect 17500 25434 17552 25440
rect 17500 25288 17552 25294
rect 17500 25230 17552 25236
rect 17512 24206 17540 25230
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17604 23730 17632 39306
rect 17788 36786 17816 47126
rect 18708 47054 18736 49200
rect 19996 48226 20024 49200
rect 19996 48198 20116 48226
rect 20088 47122 20116 48198
rect 20260 47184 20312 47190
rect 20260 47126 20312 47132
rect 20076 47116 20128 47122
rect 20076 47058 20128 47064
rect 18696 47048 18748 47054
rect 18696 46990 18748 46996
rect 19984 47048 20036 47054
rect 19984 46990 20036 46996
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19616 46504 19668 46510
rect 19616 46446 19668 46452
rect 19628 46170 19656 46446
rect 19616 46164 19668 46170
rect 19616 46106 19668 46112
rect 18788 45960 18840 45966
rect 18788 45902 18840 45908
rect 18328 45552 18380 45558
rect 18328 45494 18380 45500
rect 18340 39506 18368 45494
rect 18420 40044 18472 40050
rect 18420 39986 18472 39992
rect 18328 39500 18380 39506
rect 18328 39442 18380 39448
rect 18432 39438 18460 39986
rect 18420 39432 18472 39438
rect 18420 39374 18472 39380
rect 18432 38962 18460 39374
rect 18420 38956 18472 38962
rect 18420 38898 18472 38904
rect 18432 38554 18460 38898
rect 18420 38548 18472 38554
rect 18420 38490 18472 38496
rect 18696 38208 18748 38214
rect 18696 38150 18748 38156
rect 18144 37936 18196 37942
rect 18144 37878 18196 37884
rect 18156 36922 18184 37878
rect 18604 37664 18656 37670
rect 18604 37606 18656 37612
rect 18616 37346 18644 37606
rect 18708 37398 18736 38150
rect 18236 37324 18288 37330
rect 18236 37266 18288 37272
rect 18524 37318 18644 37346
rect 18696 37392 18748 37398
rect 18696 37334 18748 37340
rect 18144 36916 18196 36922
rect 18144 36858 18196 36864
rect 17684 36780 17736 36786
rect 17684 36722 17736 36728
rect 17776 36780 17828 36786
rect 17776 36722 17828 36728
rect 17696 35698 17724 36722
rect 17684 35692 17736 35698
rect 17684 35634 17736 35640
rect 17788 27554 17816 36722
rect 18052 36032 18104 36038
rect 18052 35974 18104 35980
rect 18064 35698 18092 35974
rect 17868 35692 17920 35698
rect 17868 35634 17920 35640
rect 18052 35692 18104 35698
rect 18052 35634 18104 35640
rect 17880 35086 17908 35634
rect 18064 35154 18092 35634
rect 18248 35442 18276 37266
rect 18524 37262 18552 37318
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 18156 35414 18276 35442
rect 18328 35488 18380 35494
rect 18328 35430 18380 35436
rect 18052 35148 18104 35154
rect 18052 35090 18104 35096
rect 17868 35080 17920 35086
rect 17868 35022 17920 35028
rect 18052 35012 18104 35018
rect 18052 34954 18104 34960
rect 17960 34604 18012 34610
rect 17960 34546 18012 34552
rect 17972 34202 18000 34546
rect 18064 34474 18092 34954
rect 18052 34468 18104 34474
rect 18052 34410 18104 34416
rect 17960 34196 18012 34202
rect 17960 34138 18012 34144
rect 18156 34134 18184 35414
rect 18236 35284 18288 35290
rect 18236 35226 18288 35232
rect 18144 34128 18196 34134
rect 18144 34070 18196 34076
rect 18156 33998 18184 34070
rect 18248 33998 18276 35226
rect 18340 34610 18368 35430
rect 18420 35148 18472 35154
rect 18420 35090 18472 35096
rect 18328 34604 18380 34610
rect 18328 34546 18380 34552
rect 18432 34490 18460 35090
rect 18524 35086 18552 37198
rect 18696 36780 18748 36786
rect 18696 36722 18748 36728
rect 18512 35080 18564 35086
rect 18512 35022 18564 35028
rect 18604 35080 18656 35086
rect 18604 35022 18656 35028
rect 18616 34746 18644 35022
rect 18604 34740 18656 34746
rect 18604 34682 18656 34688
rect 18340 34462 18460 34490
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 18236 33992 18288 33998
rect 18236 33934 18288 33940
rect 18248 33590 18276 33934
rect 18144 33584 18196 33590
rect 18144 33526 18196 33532
rect 18236 33584 18288 33590
rect 18236 33526 18288 33532
rect 17960 32836 18012 32842
rect 17960 32778 18012 32784
rect 17972 31822 18000 32778
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 17972 31142 18000 31622
rect 18064 31346 18092 32710
rect 18052 31340 18104 31346
rect 18052 31282 18104 31288
rect 17960 31136 18012 31142
rect 17960 31078 18012 31084
rect 17868 30660 17920 30666
rect 17868 30602 17920 30608
rect 17880 30394 17908 30602
rect 17868 30388 17920 30394
rect 17868 30330 17920 30336
rect 17972 28626 18000 31078
rect 18156 30666 18184 33526
rect 18248 33386 18276 33526
rect 18236 33380 18288 33386
rect 18236 33322 18288 33328
rect 18236 32904 18288 32910
rect 18236 32846 18288 32852
rect 18248 32502 18276 32846
rect 18236 32496 18288 32502
rect 18236 32438 18288 32444
rect 18340 31754 18368 34462
rect 18420 34400 18472 34406
rect 18420 34342 18472 34348
rect 18432 33402 18460 34342
rect 18616 33998 18644 34682
rect 18708 34678 18736 36722
rect 18696 34672 18748 34678
rect 18696 34614 18748 34620
rect 18604 33992 18656 33998
rect 18524 33940 18604 33946
rect 18524 33934 18656 33940
rect 18524 33918 18644 33934
rect 18524 33522 18552 33918
rect 18604 33856 18656 33862
rect 18604 33798 18656 33804
rect 18616 33658 18644 33798
rect 18604 33652 18656 33658
rect 18604 33594 18656 33600
rect 18512 33516 18564 33522
rect 18512 33458 18564 33464
rect 18432 33374 18644 33402
rect 18512 33312 18564 33318
rect 18512 33254 18564 33260
rect 18418 33008 18474 33017
rect 18418 32943 18420 32952
rect 18472 32943 18474 32952
rect 18420 32914 18472 32920
rect 18524 32910 18552 33254
rect 18616 32910 18644 33374
rect 18708 33318 18736 34614
rect 18696 33312 18748 33318
rect 18696 33254 18748 33260
rect 18512 32904 18564 32910
rect 18512 32846 18564 32852
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18340 31726 18460 31754
rect 18144 30660 18196 30666
rect 18144 30602 18196 30608
rect 18052 30592 18104 30598
rect 18052 30534 18104 30540
rect 18236 30592 18288 30598
rect 18236 30534 18288 30540
rect 18064 30138 18092 30534
rect 18248 30258 18276 30534
rect 18236 30252 18288 30258
rect 18236 30194 18288 30200
rect 18064 30110 18184 30138
rect 18052 30048 18104 30054
rect 18052 29990 18104 29996
rect 17960 28620 18012 28626
rect 17960 28562 18012 28568
rect 18064 28422 18092 29990
rect 18156 29646 18184 30110
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 18156 28744 18184 29582
rect 18328 29572 18380 29578
rect 18328 29514 18380 29520
rect 18236 28756 18288 28762
rect 18156 28716 18236 28744
rect 18236 28698 18288 28704
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 17788 27526 17908 27554
rect 17776 27464 17828 27470
rect 17776 27406 17828 27412
rect 17684 24880 17736 24886
rect 17684 24822 17736 24828
rect 17696 24342 17724 24822
rect 17684 24336 17736 24342
rect 17684 24278 17736 24284
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 17684 23656 17736 23662
rect 17684 23598 17736 23604
rect 17696 22574 17724 23598
rect 17684 22568 17736 22574
rect 17684 22510 17736 22516
rect 17788 20602 17816 27406
rect 17880 26330 17908 27526
rect 18340 26382 18368 29514
rect 18328 26376 18380 26382
rect 17880 26302 18000 26330
rect 18328 26318 18380 26324
rect 17868 26240 17920 26246
rect 17868 26182 17920 26188
rect 17880 25974 17908 26182
rect 17868 25968 17920 25974
rect 17868 25910 17920 25916
rect 17972 25786 18000 26302
rect 18340 25922 18368 26318
rect 17880 25758 18000 25786
rect 18248 25894 18368 25922
rect 17880 23662 17908 25758
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 18248 23322 18276 25894
rect 18328 25832 18380 25838
rect 18328 25774 18380 25780
rect 18340 25362 18368 25774
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 18340 24954 18368 25298
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 18432 24614 18460 31726
rect 18616 31482 18644 32846
rect 18696 31816 18748 31822
rect 18696 31758 18748 31764
rect 18708 31482 18736 31758
rect 18604 31476 18656 31482
rect 18604 31418 18656 31424
rect 18696 31476 18748 31482
rect 18696 31418 18748 31424
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18524 29850 18552 30194
rect 18512 29844 18564 29850
rect 18512 29786 18564 29792
rect 18604 28076 18656 28082
rect 18604 28018 18656 28024
rect 18512 26240 18564 26246
rect 18512 26182 18564 26188
rect 18524 25974 18552 26182
rect 18512 25968 18564 25974
rect 18512 25910 18564 25916
rect 18616 25294 18644 28018
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 18616 24274 18644 25230
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18616 23594 18644 24210
rect 18604 23588 18656 23594
rect 18604 23530 18656 23536
rect 18236 23316 18288 23322
rect 18236 23258 18288 23264
rect 18248 22642 18276 23258
rect 18800 22642 18828 45902
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 18972 40112 19024 40118
rect 18972 40054 19024 40060
rect 18880 34604 18932 34610
rect 18880 34546 18932 34552
rect 18892 32910 18920 34546
rect 18984 34490 19012 40054
rect 19156 40044 19208 40050
rect 19156 39986 19208 39992
rect 19168 38894 19196 39986
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19156 38888 19208 38894
rect 19156 38830 19208 38836
rect 19064 36032 19116 36038
rect 19064 35974 19116 35980
rect 19076 35766 19104 35974
rect 19064 35760 19116 35766
rect 19064 35702 19116 35708
rect 19064 35624 19116 35630
rect 19064 35566 19116 35572
rect 19076 35154 19104 35566
rect 19064 35148 19116 35154
rect 19064 35090 19116 35096
rect 19064 34944 19116 34950
rect 19064 34886 19116 34892
rect 19076 34678 19104 34886
rect 19064 34672 19116 34678
rect 19064 34614 19116 34620
rect 18984 34462 19104 34490
rect 18972 33516 19024 33522
rect 18972 33458 19024 33464
rect 18880 32904 18932 32910
rect 18880 32846 18932 32852
rect 18892 32570 18920 32846
rect 18984 32774 19012 33458
rect 18972 32768 19024 32774
rect 19076 32745 19104 34462
rect 18972 32710 19024 32716
rect 19062 32736 19118 32745
rect 18880 32564 18932 32570
rect 18880 32506 18932 32512
rect 18880 32224 18932 32230
rect 18880 32166 18932 32172
rect 18892 31890 18920 32166
rect 18984 31890 19012 32710
rect 19062 32671 19118 32680
rect 19064 32564 19116 32570
rect 19064 32506 19116 32512
rect 18880 31884 18932 31890
rect 18880 31826 18932 31832
rect 18972 31884 19024 31890
rect 18972 31826 19024 31832
rect 18970 31784 19026 31793
rect 18970 31719 19026 31728
rect 18880 28484 18932 28490
rect 18880 28426 18932 28432
rect 18892 28218 18920 28426
rect 18880 28212 18932 28218
rect 18880 28154 18932 28160
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 17868 22500 17920 22506
rect 17868 22442 17920 22448
rect 17880 20942 17908 22442
rect 17960 22092 18012 22098
rect 18800 22094 18828 22578
rect 18800 22066 18920 22094
rect 17960 22034 18012 22040
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17236 19854 17264 20402
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17236 19378 17264 19790
rect 17696 19786 17724 20334
rect 17788 19922 17816 20538
rect 17880 20466 17908 20878
rect 17972 20534 18000 22034
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 17960 20528 18012 20534
rect 17960 20470 18012 20476
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 18064 19922 18092 20334
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 17684 19780 17736 19786
rect 17604 19740 17684 19768
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17328 18698 17356 19110
rect 17316 18692 17368 18698
rect 17316 18634 17368 18640
rect 17328 18358 17356 18634
rect 17316 18352 17368 18358
rect 17316 18294 17368 18300
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17236 16590 17264 17546
rect 17328 17270 17356 18294
rect 17316 17264 17368 17270
rect 17316 17206 17368 17212
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17500 16516 17552 16522
rect 17500 16458 17552 16464
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17236 15162 17264 15982
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17236 14550 17264 14758
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17236 13734 17264 14282
rect 17328 14006 17356 14554
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 13326 17264 13670
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17328 12850 17356 13942
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17420 12986 17448 13330
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 16960 12406 17080 12434
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15304 3534 15332 3674
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15212 2582 15240 2926
rect 15488 2650 15516 3402
rect 16960 2650 16988 12406
rect 17328 11694 17356 12786
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17052 11218 17080 11494
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 17512 8294 17540 16458
rect 17604 14822 17632 19740
rect 17684 19722 17736 19728
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17604 6914 17632 14758
rect 17696 14074 17724 18566
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17788 17270 17816 17546
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17880 15094 17908 17682
rect 18064 16726 18092 19858
rect 18236 18692 18288 18698
rect 18236 18634 18288 18640
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 18156 17542 18184 18022
rect 18248 17678 18276 18634
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 18156 16522 18184 17206
rect 18248 17066 18276 17614
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 18340 16946 18368 21422
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18432 19378 18460 19654
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18524 19366 18828 19394
rect 18524 19258 18552 19366
rect 18800 19310 18828 19366
rect 18432 19242 18552 19258
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18420 19236 18552 19242
rect 18472 19230 18552 19236
rect 18420 19178 18472 19184
rect 18708 18970 18736 19246
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18512 16992 18564 16998
rect 18340 16918 18460 16946
rect 18512 16934 18564 16940
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18144 16516 18196 16522
rect 18144 16458 18196 16464
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17788 14482 17816 14962
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17880 14346 17908 15030
rect 17972 15026 18000 16390
rect 18156 16250 18184 16458
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 18064 15162 18092 15982
rect 18156 15570 18184 16186
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17868 14340 17920 14346
rect 17868 14282 17920 14288
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17880 13870 17908 14282
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17880 12986 17908 13806
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17972 12866 18000 14214
rect 18156 13954 18184 15370
rect 17880 12850 18000 12866
rect 17868 12844 18000 12850
rect 17920 12838 18000 12844
rect 18064 13926 18184 13954
rect 17868 12786 17920 12792
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17972 11762 18000 11834
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17972 10062 18000 11698
rect 18064 10146 18092 13926
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18156 12918 18184 13126
rect 18248 12986 18276 13262
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18156 10266 18184 10542
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18064 10118 18184 10146
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17604 6886 17724 6914
rect 17130 3496 17186 3505
rect 17130 3431 17132 3440
rect 17184 3431 17186 3440
rect 17132 3402 17184 3408
rect 17314 3088 17370 3097
rect 17314 3023 17316 3032
rect 17368 3023 17370 3032
rect 17316 2994 17368 3000
rect 17696 2990 17724 6886
rect 18156 6866 18184 10118
rect 18340 6914 18368 16662
rect 18248 6886 18368 6914
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17972 3194 18000 3470
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18248 3097 18276 6886
rect 18432 4078 18460 16918
rect 18524 16590 18552 16934
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18524 16454 18552 16526
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18524 10742 18552 16390
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18616 15706 18644 16050
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18800 6914 18828 18158
rect 18892 15638 18920 22066
rect 18984 16046 19012 31719
rect 19076 19310 19104 32506
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 19076 17338 19104 18226
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18984 15366 19012 15982
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18708 6886 18828 6914
rect 19168 6914 19196 38830
rect 19996 38350 20024 46990
rect 20076 46368 20128 46374
rect 20076 46310 20128 46316
rect 20088 46034 20116 46310
rect 20076 46028 20128 46034
rect 20076 45970 20128 45976
rect 19984 38344 20036 38350
rect 19984 38286 20036 38292
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19984 37392 20036 37398
rect 20036 37352 20208 37380
rect 19984 37334 20036 37340
rect 20180 37262 20208 37352
rect 19800 37256 19852 37262
rect 20168 37256 20220 37262
rect 19852 37216 20024 37244
rect 19800 37198 19852 37204
rect 19340 37188 19392 37194
rect 19340 37130 19392 37136
rect 19248 36236 19300 36242
rect 19248 36178 19300 36184
rect 19260 35834 19288 36178
rect 19248 35828 19300 35834
rect 19248 35770 19300 35776
rect 19352 35766 19380 37130
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19996 36922 20024 37216
rect 20168 37198 20220 37204
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19340 35760 19392 35766
rect 19340 35702 19392 35708
rect 19800 35556 19852 35562
rect 19800 35498 19852 35504
rect 19812 35290 19840 35498
rect 19800 35284 19852 35290
rect 19800 35226 19852 35232
rect 19984 34944 20036 34950
rect 19984 34886 20036 34892
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19996 34678 20024 34886
rect 19984 34672 20036 34678
rect 19984 34614 20036 34620
rect 19248 34468 19300 34474
rect 19248 34410 19300 34416
rect 19260 33658 19288 34410
rect 19340 33924 19392 33930
rect 19340 33866 19392 33872
rect 19352 33674 19380 33866
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19248 33652 19300 33658
rect 19352 33646 19472 33674
rect 19248 33594 19300 33600
rect 19260 32230 19288 33594
rect 19340 33516 19392 33522
rect 19340 33458 19392 33464
rect 19352 32842 19380 33458
rect 19444 33386 19472 33646
rect 19432 33380 19484 33386
rect 19432 33322 19484 33328
rect 19340 32836 19392 32842
rect 19340 32778 19392 32784
rect 19444 32502 19472 33322
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 19524 32360 19576 32366
rect 19522 32328 19524 32337
rect 19576 32328 19578 32337
rect 19522 32263 19578 32272
rect 19248 32224 19300 32230
rect 19248 32166 19300 32172
rect 19708 32224 19760 32230
rect 20168 32224 20220 32230
rect 19708 32166 19760 32172
rect 20166 32192 20168 32201
rect 20220 32192 20222 32201
rect 19720 32065 19748 32166
rect 20166 32127 20222 32136
rect 19706 32056 19762 32065
rect 19706 31991 19762 32000
rect 19720 31822 19748 31991
rect 20180 31890 20208 32127
rect 20168 31884 20220 31890
rect 20168 31826 20220 31832
rect 19708 31816 19760 31822
rect 19708 31758 19760 31764
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19340 31272 19392 31278
rect 19338 31240 19340 31249
rect 19392 31240 19394 31249
rect 19338 31175 19394 31184
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19984 29572 20036 29578
rect 19984 29514 20036 29520
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19996 29102 20024 29514
rect 20168 29164 20220 29170
rect 20168 29106 20220 29112
rect 19984 29096 20036 29102
rect 19984 29038 20036 29044
rect 20180 29034 20208 29106
rect 20168 29028 20220 29034
rect 20168 28970 20220 28976
rect 19248 28552 19300 28558
rect 19248 28494 19300 28500
rect 19260 25294 19288 28494
rect 19984 28484 20036 28490
rect 19984 28426 20036 28432
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19996 28218 20024 28426
rect 19984 28212 20036 28218
rect 19984 28154 20036 28160
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 20272 26908 20300 47126
rect 20444 47048 20496 47054
rect 20444 46990 20496 46996
rect 20352 37256 20404 37262
rect 20352 37198 20404 37204
rect 20364 36310 20392 37198
rect 20352 36304 20404 36310
rect 20352 36246 20404 36252
rect 20364 35698 20392 36246
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 20352 35012 20404 35018
rect 20352 34954 20404 34960
rect 20364 34610 20392 34954
rect 20352 34604 20404 34610
rect 20352 34546 20404 34552
rect 20456 31414 20484 46990
rect 20640 46510 20668 49200
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 21284 46034 21312 49200
rect 22928 46980 22980 46986
rect 22928 46922 22980 46928
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 22744 39500 22796 39506
rect 22744 39442 22796 39448
rect 20628 39364 20680 39370
rect 20628 39306 20680 39312
rect 20536 38208 20588 38214
rect 20536 38150 20588 38156
rect 20548 37942 20576 38150
rect 20536 37936 20588 37942
rect 20536 37878 20588 37884
rect 20536 37800 20588 37806
rect 20536 37742 20588 37748
rect 20548 37398 20576 37742
rect 20536 37392 20588 37398
rect 20536 37334 20588 37340
rect 20536 31680 20588 31686
rect 20536 31622 20588 31628
rect 20444 31408 20496 31414
rect 20444 31350 20496 31356
rect 20548 30666 20576 31622
rect 20536 30660 20588 30666
rect 20536 30602 20588 30608
rect 20536 29300 20588 29306
rect 20536 29242 20588 29248
rect 20548 29102 20576 29242
rect 20536 29096 20588 29102
rect 20536 29038 20588 29044
rect 20272 26880 20392 26908
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19260 24750 19288 25230
rect 19444 25226 19472 26182
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19352 23032 19380 23462
rect 19444 23186 19472 24142
rect 20076 24132 20128 24138
rect 20076 24074 20128 24080
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 20088 23594 20116 24074
rect 20076 23588 20128 23594
rect 20076 23530 20128 23536
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19432 23044 19484 23050
rect 19352 23004 19432 23032
rect 19432 22986 19484 22992
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19996 22642 20024 22918
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 19260 21622 19288 21966
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19904 20890 19932 21490
rect 19996 21146 20024 21966
rect 20088 21894 20116 23530
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20088 21010 20116 21830
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20398 19380 20742
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19444 19854 19472 20878
rect 19904 20862 20116 20890
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19984 20324 20036 20330
rect 19984 20266 20036 20272
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19260 18834 19288 19246
rect 19444 18834 19472 19790
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19996 19514 20024 20266
rect 20088 20262 20116 20862
rect 20180 20534 20208 23462
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 20272 22642 20300 23258
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20168 20528 20220 20534
rect 20168 20470 20220 20476
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 20088 19990 20116 20198
rect 20076 19984 20128 19990
rect 20076 19926 20128 19932
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19340 18760 19392 18766
rect 19260 18708 19340 18714
rect 19260 18702 19392 18708
rect 19260 18686 19380 18702
rect 19432 18692 19484 18698
rect 19260 18290 19288 18686
rect 19432 18634 19484 18640
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19260 17610 19288 18226
rect 19352 18086 19380 18294
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19444 17882 19472 18634
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19536 17746 19564 18022
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19524 17740 19576 17746
rect 19524 17682 19576 17688
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19352 16658 19380 17682
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19996 17338 20024 18770
rect 20088 18358 20116 19382
rect 20076 18352 20128 18358
rect 20076 18294 20128 18300
rect 20180 18290 20208 19654
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19996 17202 20024 17274
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19260 16250 19288 16526
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19444 16114 19472 16934
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19996 16182 20024 16594
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 20180 15502 20208 18226
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 19260 14414 19288 15438
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19260 13462 19288 14350
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19352 13530 19380 13806
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 19444 12918 19472 14214
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 20088 13530 20116 13942
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 20272 12434 20300 22578
rect 20364 20058 20392 26880
rect 20444 24880 20496 24886
rect 20444 24822 20496 24828
rect 20456 24342 20484 24822
rect 20444 24336 20496 24342
rect 20444 24278 20496 24284
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20456 20942 20484 21626
rect 20444 20936 20496 20942
rect 20444 20878 20496 20884
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20456 19922 20484 20470
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 20364 19446 20392 19722
rect 20352 19440 20404 19446
rect 20352 19382 20404 19388
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 20548 17814 20576 18566
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 14482 20484 16390
rect 20444 14476 20496 14482
rect 20444 14418 20496 14424
rect 20456 13258 20484 14418
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 20272 12406 20392 12434
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 20364 6914 20392 12406
rect 20640 11898 20668 39306
rect 22192 39296 22244 39302
rect 22192 39238 22244 39244
rect 22468 39296 22520 39302
rect 22468 39238 22520 39244
rect 22652 39296 22704 39302
rect 22652 39238 22704 39244
rect 21824 38888 21876 38894
rect 21824 38830 21876 38836
rect 22100 38888 22152 38894
rect 22100 38830 22152 38836
rect 21836 38486 21864 38830
rect 21088 38480 21140 38486
rect 21088 38422 21140 38428
rect 21824 38480 21876 38486
rect 21824 38422 21876 38428
rect 20904 38412 20956 38418
rect 20904 38354 20956 38360
rect 20916 37738 20944 38354
rect 20904 37732 20956 37738
rect 20904 37674 20956 37680
rect 21100 37670 21128 38422
rect 21180 38344 21232 38350
rect 21180 38286 21232 38292
rect 21192 37874 21220 38286
rect 22112 38214 22140 38830
rect 22204 38350 22232 39238
rect 22480 39098 22508 39238
rect 22468 39092 22520 39098
rect 22468 39034 22520 39040
rect 22192 38344 22244 38350
rect 22192 38286 22244 38292
rect 22100 38208 22152 38214
rect 22100 38150 22152 38156
rect 22480 37874 22508 39034
rect 22560 39024 22612 39030
rect 22560 38966 22612 38972
rect 22572 38010 22600 38966
rect 22664 38554 22692 39238
rect 22652 38548 22704 38554
rect 22652 38490 22704 38496
rect 22560 38004 22612 38010
rect 22560 37946 22612 37952
rect 21180 37868 21232 37874
rect 21180 37810 21232 37816
rect 22468 37868 22520 37874
rect 22468 37810 22520 37816
rect 22652 37868 22704 37874
rect 22652 37810 22704 37816
rect 20812 37664 20864 37670
rect 20812 37606 20864 37612
rect 21088 37664 21140 37670
rect 21088 37606 21140 37612
rect 20824 36258 20852 37606
rect 20732 36230 20852 36258
rect 20732 35630 20760 36230
rect 20720 35624 20772 35630
rect 20720 35566 20772 35572
rect 20732 35154 20760 35566
rect 20720 35148 20772 35154
rect 20720 35090 20772 35096
rect 21088 35148 21140 35154
rect 21088 35090 21140 35096
rect 20996 35012 21048 35018
rect 20996 34954 21048 34960
rect 21008 34202 21036 34954
rect 21100 34746 21128 35090
rect 21088 34740 21140 34746
rect 21088 34682 21140 34688
rect 21088 34604 21140 34610
rect 21192 34592 21220 37810
rect 22100 37800 22152 37806
rect 22100 37742 22152 37748
rect 21272 37664 21324 37670
rect 21272 37606 21324 37612
rect 21284 37330 21312 37606
rect 22112 37398 22140 37742
rect 22664 37398 22692 37810
rect 22100 37392 22152 37398
rect 22100 37334 22152 37340
rect 22652 37392 22704 37398
rect 22652 37334 22704 37340
rect 21272 37324 21324 37330
rect 21272 37266 21324 37272
rect 22284 37324 22336 37330
rect 22284 37266 22336 37272
rect 22296 37194 22324 37266
rect 22664 37194 22692 37334
rect 22756 37194 22784 39442
rect 22284 37188 22336 37194
rect 22284 37130 22336 37136
rect 22652 37188 22704 37194
rect 22652 37130 22704 37136
rect 22744 37188 22796 37194
rect 22744 37130 22796 37136
rect 21732 37120 21784 37126
rect 21732 37062 21784 37068
rect 21744 36786 21772 37062
rect 21732 36780 21784 36786
rect 21732 36722 21784 36728
rect 22756 36174 22784 37130
rect 22940 36242 22968 46922
rect 24952 46504 25004 46510
rect 24952 46446 25004 46452
rect 24964 46170 24992 46446
rect 24952 46164 25004 46170
rect 24952 46106 25004 46112
rect 25148 46102 25176 49200
rect 25688 47048 25740 47054
rect 25688 46990 25740 46996
rect 25412 46164 25464 46170
rect 25412 46106 25464 46112
rect 25136 46096 25188 46102
rect 25136 46038 25188 46044
rect 25424 45558 25452 46106
rect 25700 46034 25728 46990
rect 25792 46510 25820 49200
rect 27080 46918 27108 49200
rect 28368 47054 28396 49200
rect 29368 47252 29420 47258
rect 29368 47194 29420 47200
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 27068 46912 27120 46918
rect 27068 46854 27120 46860
rect 27620 46912 27672 46918
rect 27620 46854 27672 46860
rect 28264 46912 28316 46918
rect 28264 46854 28316 46860
rect 25780 46504 25832 46510
rect 25780 46446 25832 46452
rect 25688 46028 25740 46034
rect 25688 45970 25740 45976
rect 27068 45892 27120 45898
rect 27068 45834 27120 45840
rect 27080 45558 27108 45834
rect 25412 45552 25464 45558
rect 25412 45494 25464 45500
rect 27068 45552 27120 45558
rect 27068 45494 27120 45500
rect 25320 45484 25372 45490
rect 25320 45426 25372 45432
rect 26516 45484 26568 45490
rect 26516 45426 26568 45432
rect 25332 45354 25360 45426
rect 25320 45348 25372 45354
rect 25320 45290 25372 45296
rect 25332 40050 25360 45290
rect 25596 43308 25648 43314
rect 25596 43250 25648 43256
rect 25320 40044 25372 40050
rect 25320 39986 25372 39992
rect 24860 38752 24912 38758
rect 24860 38694 24912 38700
rect 24492 38548 24544 38554
rect 24492 38490 24544 38496
rect 23480 38412 23532 38418
rect 23480 38354 23532 38360
rect 23296 38208 23348 38214
rect 23296 38150 23348 38156
rect 23308 38010 23336 38150
rect 23296 38004 23348 38010
rect 23296 37946 23348 37952
rect 23492 37874 23520 38354
rect 24504 38010 24532 38490
rect 24872 38282 24900 38694
rect 25412 38412 25464 38418
rect 25412 38354 25464 38360
rect 24860 38276 24912 38282
rect 24860 38218 24912 38224
rect 25320 38276 25372 38282
rect 25320 38218 25372 38224
rect 25332 38010 25360 38218
rect 24492 38004 24544 38010
rect 24492 37946 24544 37952
rect 25320 38004 25372 38010
rect 25320 37946 25372 37952
rect 23480 37868 23532 37874
rect 23480 37810 23532 37816
rect 24504 37738 24532 37946
rect 24584 37868 24636 37874
rect 24584 37810 24636 37816
rect 24676 37868 24728 37874
rect 24676 37810 24728 37816
rect 24308 37732 24360 37738
rect 24308 37674 24360 37680
rect 24492 37732 24544 37738
rect 24492 37674 24544 37680
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 22928 36236 22980 36242
rect 22928 36178 22980 36184
rect 22468 36168 22520 36174
rect 22468 36110 22520 36116
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 22480 35698 22508 36110
rect 22928 36032 22980 36038
rect 22928 35974 22980 35980
rect 22468 35692 22520 35698
rect 22468 35634 22520 35640
rect 22560 35692 22612 35698
rect 22560 35634 22612 35640
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22376 35624 22428 35630
rect 22376 35566 22428 35572
rect 22284 35488 22336 35494
rect 22284 35430 22336 35436
rect 22192 35284 22244 35290
rect 22192 35226 22244 35232
rect 21456 35012 21508 35018
rect 21456 34954 21508 34960
rect 21468 34746 21496 34954
rect 21456 34740 21508 34746
rect 21456 34682 21508 34688
rect 21140 34564 21220 34592
rect 22100 34604 22152 34610
rect 21088 34546 21140 34552
rect 22100 34546 22152 34552
rect 20996 34196 21048 34202
rect 20996 34138 21048 34144
rect 21100 34082 21128 34546
rect 21732 34400 21784 34406
rect 21732 34342 21784 34348
rect 21744 34202 21772 34342
rect 21732 34196 21784 34202
rect 21732 34138 21784 34144
rect 21008 34054 21128 34082
rect 20812 32972 20864 32978
rect 20812 32914 20864 32920
rect 20720 31748 20772 31754
rect 20720 31690 20772 31696
rect 20732 30734 20760 31690
rect 20824 31210 20852 32914
rect 21008 32774 21036 34054
rect 21088 33924 21140 33930
rect 21088 33866 21140 33872
rect 20996 32768 21048 32774
rect 20996 32710 21048 32716
rect 21008 32570 21036 32710
rect 20996 32564 21048 32570
rect 20996 32506 21048 32512
rect 20996 32020 21048 32026
rect 20996 31962 21048 31968
rect 21100 32008 21128 33866
rect 21546 33008 21602 33017
rect 21546 32943 21548 32952
rect 21600 32943 21602 32952
rect 21548 32914 21600 32920
rect 22112 32298 22140 34546
rect 22204 32366 22232 35226
rect 22296 34066 22324 35430
rect 22388 34202 22416 35566
rect 22572 35290 22600 35634
rect 22560 35284 22612 35290
rect 22560 35226 22612 35232
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22480 34542 22508 34886
rect 22572 34678 22600 35226
rect 22560 34672 22612 34678
rect 22560 34614 22612 34620
rect 22468 34536 22520 34542
rect 22468 34478 22520 34484
rect 22376 34196 22428 34202
rect 22376 34138 22428 34144
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22388 33522 22416 34138
rect 22480 33946 22508 34478
rect 22848 34202 22876 35634
rect 22836 34196 22888 34202
rect 22836 34138 22888 34144
rect 22480 33918 22692 33946
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22376 33516 22428 33522
rect 22376 33458 22428 33464
rect 22284 33312 22336 33318
rect 22284 33254 22336 33260
rect 22296 33114 22324 33254
rect 22284 33108 22336 33114
rect 22284 33050 22336 33056
rect 22296 32978 22324 33050
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22376 32768 22428 32774
rect 22376 32710 22428 32716
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 22192 32360 22244 32366
rect 22190 32328 22192 32337
rect 22244 32328 22246 32337
rect 22100 32292 22152 32298
rect 22190 32263 22246 32272
rect 22100 32234 22152 32240
rect 21180 32020 21232 32026
rect 21100 31980 21180 32008
rect 21008 31754 21036 31962
rect 20916 31726 21036 31754
rect 20812 31204 20864 31210
rect 20812 31146 20864 31152
rect 20720 30728 20772 30734
rect 20720 30670 20772 30676
rect 20824 30569 20852 31146
rect 20916 30818 20944 31726
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 21008 30920 21036 31282
rect 21100 31210 21128 31980
rect 21180 31962 21232 31968
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 21088 31204 21140 31210
rect 21088 31146 21140 31152
rect 22020 31142 22048 31282
rect 22008 31136 22060 31142
rect 22008 31078 22060 31084
rect 21008 30892 21220 30920
rect 20916 30790 21128 30818
rect 20810 30560 20866 30569
rect 20810 30495 20866 30504
rect 20720 29640 20772 29646
rect 20904 29640 20956 29646
rect 20720 29582 20772 29588
rect 20824 29600 20904 29628
rect 20732 29306 20760 29582
rect 20720 29300 20772 29306
rect 20720 29242 20772 29248
rect 20732 28762 20760 29242
rect 20720 28756 20772 28762
rect 20720 28698 20772 28704
rect 20732 28150 20760 28698
rect 20824 28694 20852 29600
rect 20904 29582 20956 29588
rect 20904 28960 20956 28966
rect 20904 28902 20956 28908
rect 20812 28688 20864 28694
rect 20812 28630 20864 28636
rect 20720 28144 20772 28150
rect 20720 28086 20772 28092
rect 20824 28082 20852 28630
rect 20916 28626 20944 28902
rect 20904 28620 20956 28626
rect 20904 28562 20956 28568
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 21100 28014 21128 30790
rect 21192 30598 21220 30892
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 21272 30660 21324 30666
rect 21272 30602 21324 30608
rect 21180 30592 21232 30598
rect 21180 30534 21232 30540
rect 21284 30054 21312 30602
rect 21928 30258 21956 30670
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 22112 30054 22140 32234
rect 22296 31890 22324 32506
rect 22388 32298 22416 32710
rect 22376 32292 22428 32298
rect 22376 32234 22428 32240
rect 22284 31884 22336 31890
rect 22284 31826 22336 31832
rect 22296 30666 22324 31826
rect 22480 31385 22508 33798
rect 22560 32360 22612 32366
rect 22560 32302 22612 32308
rect 22466 31376 22522 31385
rect 22466 31311 22522 31320
rect 22468 31272 22520 31278
rect 22468 31214 22520 31220
rect 22376 30932 22428 30938
rect 22376 30874 22428 30880
rect 22388 30841 22416 30874
rect 22374 30832 22430 30841
rect 22374 30767 22430 30776
rect 22480 30682 22508 31214
rect 22284 30660 22336 30666
rect 22284 30602 22336 30608
rect 22388 30654 22508 30682
rect 22190 30424 22246 30433
rect 22190 30359 22246 30368
rect 21272 30048 21324 30054
rect 21272 29990 21324 29996
rect 22100 30048 22152 30054
rect 22100 29990 22152 29996
rect 22204 29714 22232 30359
rect 22192 29708 22244 29714
rect 22192 29650 22244 29656
rect 22100 29640 22152 29646
rect 22100 29582 22152 29588
rect 21548 29504 21600 29510
rect 21548 29446 21600 29452
rect 21560 28762 21588 29446
rect 22112 29306 22140 29582
rect 22192 29572 22244 29578
rect 22192 29514 22244 29520
rect 22100 29300 22152 29306
rect 22100 29242 22152 29248
rect 22204 29238 22232 29514
rect 22192 29232 22244 29238
rect 22192 29174 22244 29180
rect 22296 29170 22324 30602
rect 22388 30190 22416 30654
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22376 30184 22428 30190
rect 22376 30126 22428 30132
rect 22284 29164 22336 29170
rect 22284 29106 22336 29112
rect 22388 29050 22416 30126
rect 22480 29850 22508 30194
rect 22468 29844 22520 29850
rect 22468 29786 22520 29792
rect 22468 29640 22520 29646
rect 22468 29582 22520 29588
rect 22008 29028 22060 29034
rect 22008 28970 22060 28976
rect 22100 29028 22152 29034
rect 22100 28970 22152 28976
rect 22296 29022 22416 29050
rect 22480 29034 22508 29582
rect 22468 29028 22520 29034
rect 22020 28762 22048 28970
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 22008 28756 22060 28762
rect 22008 28698 22060 28704
rect 22112 28626 22140 28970
rect 22296 28966 22324 29022
rect 22468 28970 22520 28976
rect 22284 28960 22336 28966
rect 22284 28902 22336 28908
rect 22376 28960 22428 28966
rect 22376 28902 22428 28908
rect 22388 28762 22416 28902
rect 22376 28756 22428 28762
rect 22376 28698 22428 28704
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20732 26042 20760 26930
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 20824 22574 20852 26726
rect 20996 26240 21048 26246
rect 20996 26182 21048 26188
rect 21008 25498 21036 26182
rect 20996 25492 21048 25498
rect 20996 25434 21048 25440
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20824 19378 20852 22374
rect 20916 22098 20944 22578
rect 21100 22438 21128 27950
rect 22112 26858 22140 28154
rect 22204 27878 22232 28494
rect 22192 27872 22244 27878
rect 22192 27814 22244 27820
rect 22204 27538 22232 27814
rect 22388 27674 22416 28698
rect 22468 28416 22520 28422
rect 22468 28358 22520 28364
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22192 27532 22244 27538
rect 22192 27474 22244 27480
rect 22204 26858 22232 27474
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22296 26994 22324 27270
rect 22388 27062 22416 27610
rect 22376 27056 22428 27062
rect 22376 26998 22428 27004
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 22100 26852 22152 26858
rect 22100 26794 22152 26800
rect 22192 26852 22244 26858
rect 22192 26794 22244 26800
rect 22112 26382 22140 26794
rect 22296 26586 22324 26930
rect 22284 26580 22336 26586
rect 22284 26522 22336 26528
rect 21640 26376 21692 26382
rect 21640 26318 21692 26324
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 21284 25838 21312 26250
rect 21272 25832 21324 25838
rect 21272 25774 21324 25780
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 21192 25158 21220 25638
rect 21284 25294 21312 25774
rect 21272 25288 21324 25294
rect 21272 25230 21324 25236
rect 21180 25152 21232 25158
rect 21180 25094 21232 25100
rect 21284 24954 21312 25230
rect 21272 24948 21324 24954
rect 21272 24890 21324 24896
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 20904 22092 20956 22098
rect 20904 22034 20956 22040
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 21008 21146 21036 21898
rect 21088 21344 21140 21350
rect 21088 21286 21140 21292
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 21100 20602 21128 21286
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 20824 19258 20852 19314
rect 20732 19230 20852 19258
rect 20732 18834 20760 19230
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20824 18222 20852 19110
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20916 18290 20944 18702
rect 21008 18630 21036 19314
rect 21088 19236 21140 19242
rect 21088 19178 21140 19184
rect 21100 18834 21128 19178
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20824 17746 20852 18158
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20824 15706 20852 16050
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 19168 6886 19288 6914
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18234 3088 18290 3097
rect 18340 3058 18368 3334
rect 18234 3023 18290 3032
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 17684 2984 17736 2990
rect 17684 2926 17736 2932
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15488 800 15516 2382
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16132 800 16160 2314
rect 17420 800 17448 2790
rect 18524 2650 18552 4558
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18616 3194 18644 3470
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18708 800 18736 6886
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18984 3194 19012 4082
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 19076 2446 19104 3878
rect 19260 3602 19288 6886
rect 19996 6886 20392 6914
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19260 3398 19288 3538
rect 19444 3534 19472 4422
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19708 4140 19760 4146
rect 19996 4128 20024 6886
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 20272 4282 20300 4558
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 19708 4082 19760 4088
rect 19904 4100 20024 4128
rect 19536 3738 19564 4082
rect 19720 3738 19748 4082
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19708 3732 19760 3738
rect 19708 3674 19760 3680
rect 19904 3670 19932 4100
rect 19984 4004 20036 4010
rect 19984 3946 20036 3952
rect 19892 3664 19944 3670
rect 19892 3606 19944 3612
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19168 3058 19196 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19996 3058 20024 3946
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20088 3602 20208 3618
rect 20088 3596 20220 3602
rect 20088 3590 20168 3596
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 20088 2938 20116 3590
rect 20168 3538 20220 3544
rect 20272 3534 20300 3878
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 20180 3194 20208 3402
rect 20548 3398 20576 3878
rect 20732 3534 20760 4422
rect 20824 4078 20852 4558
rect 20904 4548 20956 4554
rect 20904 4490 20956 4496
rect 20916 4146 20944 4490
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 21008 3738 21036 4558
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 20640 3058 20668 3334
rect 20718 3224 20774 3233
rect 20718 3159 20720 3168
rect 20772 3159 20774 3168
rect 20720 3130 20772 3136
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 19352 2910 20116 2938
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 19352 800 19380 2910
rect 21192 2854 21220 22986
rect 21272 22432 21324 22438
rect 21272 22374 21324 22380
rect 21284 22234 21312 22374
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21456 19984 21508 19990
rect 21456 19926 21508 19932
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21376 17882 21404 19314
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21376 3534 21404 4422
rect 21468 3602 21496 19926
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 21548 3596 21600 3602
rect 21548 3538 21600 3544
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21560 2990 21588 3538
rect 21548 2984 21600 2990
rect 21548 2926 21600 2932
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 19904 2650 19932 2790
rect 19892 2644 19944 2650
rect 19892 2586 19944 2592
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2790
rect 21284 2650 21312 2790
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21652 2514 21680 26318
rect 21824 26308 21876 26314
rect 21824 26250 21876 26256
rect 21836 25906 21864 26250
rect 21732 25900 21784 25906
rect 21732 25842 21784 25848
rect 21824 25900 21876 25906
rect 21824 25842 21876 25848
rect 21744 25430 21772 25842
rect 21732 25424 21784 25430
rect 21732 25366 21784 25372
rect 21732 25288 21784 25294
rect 21836 25276 21864 25842
rect 22480 25838 22508 28358
rect 22572 26874 22600 32302
rect 22664 31770 22692 33918
rect 22848 33658 22876 34138
rect 22836 33652 22888 33658
rect 22836 33594 22888 33600
rect 22848 32434 22876 33594
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22744 32224 22796 32230
rect 22744 32166 22796 32172
rect 22756 31890 22784 32166
rect 22834 31920 22890 31929
rect 22744 31884 22796 31890
rect 22834 31855 22890 31864
rect 22744 31826 22796 31832
rect 22664 31742 22784 31770
rect 22652 31136 22704 31142
rect 22652 31078 22704 31084
rect 22664 30666 22692 31078
rect 22652 30660 22704 30666
rect 22652 30602 22704 30608
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22664 28558 22692 29990
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22664 27334 22692 28018
rect 22756 27402 22784 31742
rect 22848 30433 22876 31855
rect 22834 30424 22890 30433
rect 22834 30359 22890 30368
rect 22836 30252 22888 30258
rect 22836 30194 22888 30200
rect 22848 29714 22876 30194
rect 22836 29708 22888 29714
rect 22836 29650 22888 29656
rect 22848 29238 22876 29650
rect 22940 29510 22968 35974
rect 23112 35080 23164 35086
rect 23112 35022 23164 35028
rect 23124 34610 23152 35022
rect 23216 35018 23244 37062
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 23388 36644 23440 36650
rect 23388 36586 23440 36592
rect 23296 36168 23348 36174
rect 23296 36110 23348 36116
rect 23308 36038 23336 36110
rect 23296 36032 23348 36038
rect 23296 35974 23348 35980
rect 23308 35737 23336 35974
rect 23294 35728 23350 35737
rect 23294 35663 23350 35672
rect 23400 35086 23428 36586
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 23204 35012 23256 35018
rect 23204 34954 23256 34960
rect 23112 34604 23164 34610
rect 23112 34546 23164 34552
rect 23112 33448 23164 33454
rect 23112 33390 23164 33396
rect 23020 33108 23072 33114
rect 23124 33096 23152 33390
rect 23072 33068 23152 33096
rect 23020 33050 23072 33056
rect 23216 33046 23244 34954
rect 23296 33924 23348 33930
rect 23296 33866 23348 33872
rect 23204 33040 23256 33046
rect 23204 32982 23256 32988
rect 23112 32496 23164 32502
rect 23112 32438 23164 32444
rect 23020 32224 23072 32230
rect 23020 32166 23072 32172
rect 23032 31822 23060 32166
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 23124 31754 23152 32438
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 23216 32026 23244 32370
rect 23308 32366 23336 33866
rect 23296 32360 23348 32366
rect 23296 32302 23348 32308
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23204 31816 23256 31822
rect 23204 31758 23256 31764
rect 23112 31748 23164 31754
rect 23112 31690 23164 31696
rect 23216 31482 23244 31758
rect 23204 31476 23256 31482
rect 23204 31418 23256 31424
rect 23202 31376 23258 31385
rect 23112 31340 23164 31346
rect 23202 31311 23258 31320
rect 23112 31282 23164 31288
rect 23124 31249 23152 31282
rect 23110 31240 23166 31249
rect 23110 31175 23166 31184
rect 23020 30592 23072 30598
rect 23020 30534 23072 30540
rect 23112 30592 23164 30598
rect 23112 30534 23164 30540
rect 23032 30258 23060 30534
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 23124 30190 23152 30534
rect 23112 30184 23164 30190
rect 23112 30126 23164 30132
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 22836 29232 22888 29238
rect 22836 29174 22888 29180
rect 23216 28218 23244 31311
rect 23308 30326 23336 32302
rect 23400 31929 23428 35022
rect 23492 33998 23520 36518
rect 23584 36242 23796 36258
rect 23572 36236 23796 36242
rect 23624 36230 23796 36236
rect 23572 36178 23624 36184
rect 23572 36100 23624 36106
rect 23572 36042 23624 36048
rect 23584 35222 23612 36042
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23676 35766 23704 35974
rect 23768 35834 23796 36230
rect 23756 35828 23808 35834
rect 23756 35770 23808 35776
rect 23664 35760 23716 35766
rect 23664 35702 23716 35708
rect 23572 35216 23624 35222
rect 23572 35158 23624 35164
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23756 33856 23808 33862
rect 23756 33798 23808 33804
rect 23768 33590 23796 33798
rect 23756 33584 23808 33590
rect 23756 33526 23808 33532
rect 23756 33312 23808 33318
rect 23756 33254 23808 33260
rect 23480 33040 23532 33046
rect 23480 32982 23532 32988
rect 23386 31920 23442 31929
rect 23386 31855 23442 31864
rect 23492 31770 23520 32982
rect 23400 31742 23520 31770
rect 23400 30802 23428 31742
rect 23664 31476 23716 31482
rect 23664 31418 23716 31424
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23388 30796 23440 30802
rect 23388 30738 23440 30744
rect 23296 30320 23348 30326
rect 23296 30262 23348 30268
rect 23584 30258 23612 31282
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23308 29510 23336 29582
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 23296 29164 23348 29170
rect 23296 29106 23348 29112
rect 23308 28558 23336 29106
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23204 28212 23256 28218
rect 23204 28154 23256 28160
rect 22744 27396 22796 27402
rect 22744 27338 22796 27344
rect 22652 27328 22704 27334
rect 22652 27270 22704 27276
rect 22756 26994 22784 27338
rect 23388 27328 23440 27334
rect 23388 27270 23440 27276
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22572 26846 22692 26874
rect 22468 25832 22520 25838
rect 22468 25774 22520 25780
rect 22100 25764 22152 25770
rect 22100 25706 22152 25712
rect 22112 25430 22140 25706
rect 22284 25696 22336 25702
rect 22284 25638 22336 25644
rect 22296 25498 22324 25638
rect 22284 25492 22336 25498
rect 22284 25434 22336 25440
rect 22100 25424 22152 25430
rect 22100 25366 22152 25372
rect 22560 25424 22612 25430
rect 22560 25366 22612 25372
rect 21784 25248 21864 25276
rect 21732 25230 21784 25236
rect 22572 24818 22600 25366
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21928 23798 21956 24006
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 22284 23044 22336 23050
rect 22284 22986 22336 22992
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21732 22094 21784 22098
rect 21836 22094 21864 22374
rect 22296 22234 22324 22986
rect 22376 22636 22428 22642
rect 22376 22578 22428 22584
rect 22388 22234 22416 22578
rect 22284 22228 22336 22234
rect 22284 22170 22336 22176
rect 22376 22228 22428 22234
rect 22376 22170 22428 22176
rect 21732 22092 21864 22094
rect 21784 22066 21864 22092
rect 21732 22034 21784 22040
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 21824 21888 21876 21894
rect 21824 21830 21876 21836
rect 21836 20942 21864 21830
rect 22572 21690 22600 21966
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22284 21616 22336 21622
rect 22468 21616 22520 21622
rect 22336 21564 22468 21570
rect 22284 21558 22520 21564
rect 22192 21548 22244 21554
rect 22296 21542 22508 21558
rect 22572 21554 22600 21626
rect 22560 21548 22612 21554
rect 22192 21490 22244 21496
rect 22560 21490 22612 21496
rect 22100 21412 22152 21418
rect 22100 21354 22152 21360
rect 22112 21010 22140 21354
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 22204 20806 22232 21490
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22388 21010 22416 21286
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21836 17202 21864 20538
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 21928 19922 21956 20198
rect 21916 19916 21968 19922
rect 21916 19858 21968 19864
rect 22204 19786 22232 20742
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22020 17338 22048 18702
rect 22204 17610 22232 19450
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22296 17746 22324 18566
rect 22284 17740 22336 17746
rect 22284 17682 22336 17688
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 22008 17332 22060 17338
rect 22008 17274 22060 17280
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21836 16522 21864 17138
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 22388 4146 22416 20402
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 22480 18290 22508 18566
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 21744 3398 21772 3878
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 21732 3392 21784 3398
rect 21732 3334 21784 3340
rect 22112 2990 22140 3470
rect 22204 3097 22232 3606
rect 22388 3126 22416 3878
rect 22480 3126 22508 4014
rect 22572 3738 22600 4014
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 22376 3120 22428 3126
rect 22190 3088 22246 3097
rect 22376 3062 22428 3068
rect 22468 3120 22520 3126
rect 22468 3062 22520 3068
rect 22190 3023 22246 3032
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 22466 2952 22522 2961
rect 22466 2887 22468 2896
rect 22520 2887 22522 2896
rect 22560 2916 22612 2922
rect 22468 2858 22520 2864
rect 22560 2858 22612 2864
rect 21640 2508 21692 2514
rect 21640 2450 21692 2456
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20640 800 20668 2314
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 21928 800 21956 2246
rect 22572 800 22600 2858
rect 22664 2582 22692 26846
rect 23400 26450 23428 27270
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 23400 25770 23428 26386
rect 23388 25764 23440 25770
rect 23388 25706 23440 25712
rect 22744 25696 22796 25702
rect 22744 25638 22796 25644
rect 22756 25294 22784 25638
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22836 25220 22888 25226
rect 22836 25162 22888 25168
rect 22848 24954 22876 25162
rect 22836 24948 22888 24954
rect 22836 24890 22888 24896
rect 23112 24812 23164 24818
rect 23112 24754 23164 24760
rect 23020 23520 23072 23526
rect 23020 23462 23072 23468
rect 23032 23050 23060 23462
rect 23020 23044 23072 23050
rect 23020 22986 23072 22992
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 22940 22658 22968 22714
rect 22940 22630 23060 22658
rect 22940 22522 22968 22630
rect 22848 22506 22968 22522
rect 22836 22500 22968 22506
rect 22888 22494 22968 22500
rect 22836 22442 22888 22448
rect 23032 22438 23060 22630
rect 23020 22432 23072 22438
rect 23020 22374 23072 22380
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 23032 20262 23060 20402
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 22744 4548 22796 4554
rect 22744 4490 22796 4496
rect 22756 3738 22784 4490
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 23020 4480 23072 4486
rect 23020 4422 23072 4428
rect 22848 4146 22876 4422
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22848 3233 22876 3470
rect 22834 3224 22890 3233
rect 22834 3159 22890 3168
rect 22652 2576 22704 2582
rect 22652 2518 22704 2524
rect 23032 2446 23060 4422
rect 23124 4010 23152 24754
rect 23584 24562 23612 29582
rect 23676 26518 23704 31418
rect 23768 28150 23796 33254
rect 23860 32434 23888 36858
rect 23940 32904 23992 32910
rect 23940 32846 23992 32852
rect 23848 32428 23900 32434
rect 23848 32370 23900 32376
rect 23860 30734 23888 32370
rect 23848 30728 23900 30734
rect 23848 30670 23900 30676
rect 23952 29646 23980 32846
rect 24320 31482 24348 37674
rect 24400 36576 24452 36582
rect 24400 36518 24452 36524
rect 24412 35766 24440 36518
rect 24400 35760 24452 35766
rect 24400 35702 24452 35708
rect 24596 33930 24624 37810
rect 24688 36786 24716 37810
rect 24676 36780 24728 36786
rect 24676 36722 24728 36728
rect 25424 36242 25452 38354
rect 25412 36236 25464 36242
rect 25412 36178 25464 36184
rect 24676 35828 24728 35834
rect 24676 35770 24728 35776
rect 24688 35086 24716 35770
rect 24952 35284 25004 35290
rect 24952 35226 25004 35232
rect 24676 35080 24728 35086
rect 24676 35022 24728 35028
rect 24688 34610 24716 35022
rect 24964 34746 24992 35226
rect 25320 35012 25372 35018
rect 25320 34954 25372 34960
rect 24952 34740 25004 34746
rect 24952 34682 25004 34688
rect 25332 34610 25360 34954
rect 24676 34604 24728 34610
rect 24676 34546 24728 34552
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 24584 33924 24636 33930
rect 24584 33866 24636 33872
rect 24596 31754 24624 33866
rect 25608 33522 25636 43250
rect 26528 41414 26556 45426
rect 26976 43784 27028 43790
rect 26976 43726 27028 43732
rect 26988 43246 27016 43726
rect 27632 43722 27660 46854
rect 28276 46578 28304 46854
rect 28264 46572 28316 46578
rect 28264 46514 28316 46520
rect 28080 44736 28132 44742
rect 28080 44678 28132 44684
rect 28092 44470 28120 44678
rect 28080 44464 28132 44470
rect 28080 44406 28132 44412
rect 27712 44328 27764 44334
rect 27712 44270 27764 44276
rect 27620 43716 27672 43722
rect 27620 43658 27672 43664
rect 26976 43240 27028 43246
rect 26976 43182 27028 43188
rect 26700 42152 26752 42158
rect 26700 42094 26752 42100
rect 26528 41386 26648 41414
rect 26148 38208 26200 38214
rect 26148 38150 26200 38156
rect 26332 38208 26384 38214
rect 26332 38150 26384 38156
rect 26424 38208 26476 38214
rect 26424 38150 26476 38156
rect 26160 38010 26188 38150
rect 26148 38004 26200 38010
rect 26148 37946 26200 37952
rect 26344 37874 26372 38150
rect 26332 37868 26384 37874
rect 26332 37810 26384 37816
rect 26436 37806 26464 38150
rect 26424 37800 26476 37806
rect 26424 37742 26476 37748
rect 26332 37732 26384 37738
rect 26332 37674 26384 37680
rect 26148 37664 26200 37670
rect 26148 37606 26200 37612
rect 25964 35148 26016 35154
rect 25964 35090 26016 35096
rect 25780 34944 25832 34950
rect 25780 34886 25832 34892
rect 24952 33516 25004 33522
rect 24952 33458 25004 33464
rect 25596 33516 25648 33522
rect 25596 33458 25648 33464
rect 24676 33040 24728 33046
rect 24676 32982 24728 32988
rect 24688 32434 24716 32982
rect 24964 32434 24992 33458
rect 25044 33448 25096 33454
rect 25044 33390 25096 33396
rect 25056 32978 25084 33390
rect 25228 33312 25280 33318
rect 25228 33254 25280 33260
rect 25240 33114 25268 33254
rect 25228 33108 25280 33114
rect 25228 33050 25280 33056
rect 25044 32972 25096 32978
rect 25044 32914 25096 32920
rect 25504 32904 25556 32910
rect 25504 32846 25556 32852
rect 25228 32564 25280 32570
rect 25228 32506 25280 32512
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 24860 32428 24912 32434
rect 24860 32370 24912 32376
rect 24952 32428 25004 32434
rect 24952 32370 25004 32376
rect 24504 31726 24624 31754
rect 24308 31476 24360 31482
rect 24308 31418 24360 31424
rect 23940 29640 23992 29646
rect 23940 29582 23992 29588
rect 24504 29306 24532 31726
rect 24872 31498 24900 32370
rect 24964 32201 24992 32370
rect 24950 32192 25006 32201
rect 25240 32178 25268 32506
rect 25516 32434 25544 32846
rect 25596 32496 25648 32502
rect 25596 32438 25648 32444
rect 25504 32428 25556 32434
rect 25504 32370 25556 32376
rect 24950 32127 25006 32136
rect 25056 32150 25268 32178
rect 24780 31482 24900 31498
rect 24768 31476 24900 31482
rect 24820 31470 24900 31476
rect 24768 31418 24820 31424
rect 24780 31278 24808 31418
rect 24964 31414 24992 32127
rect 24860 31408 24912 31414
rect 24860 31350 24912 31356
rect 24952 31408 25004 31414
rect 24952 31350 25004 31356
rect 24768 31272 24820 31278
rect 24768 31214 24820 31220
rect 24872 30938 24900 31350
rect 24952 31272 25004 31278
rect 24952 31214 25004 31220
rect 24860 30932 24912 30938
rect 24860 30874 24912 30880
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24596 30258 24624 30670
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24492 29300 24544 29306
rect 24492 29242 24544 29248
rect 23756 28144 23808 28150
rect 23756 28086 23808 28092
rect 23768 27470 23796 28086
rect 24504 27946 24532 29242
rect 24492 27940 24544 27946
rect 24492 27882 24544 27888
rect 24216 27872 24268 27878
rect 24216 27814 24268 27820
rect 24228 27470 24256 27814
rect 23756 27464 23808 27470
rect 23756 27406 23808 27412
rect 24216 27464 24268 27470
rect 24216 27406 24268 27412
rect 24228 27130 24256 27406
rect 24216 27124 24268 27130
rect 24216 27066 24268 27072
rect 24676 27124 24728 27130
rect 24676 27066 24728 27072
rect 23756 26784 23808 26790
rect 23756 26726 23808 26732
rect 23664 26512 23716 26518
rect 23664 26454 23716 26460
rect 23768 24750 23796 26726
rect 24688 26518 24716 27066
rect 24872 27062 24900 30874
rect 24964 29170 24992 31214
rect 24952 29164 25004 29170
rect 24952 29106 25004 29112
rect 24860 27056 24912 27062
rect 24860 26998 24912 27004
rect 24676 26512 24728 26518
rect 24676 26454 24728 26460
rect 24032 25764 24084 25770
rect 24032 25706 24084 25712
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 23584 24534 23796 24562
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23388 23656 23440 23662
rect 23388 23598 23440 23604
rect 23204 23588 23256 23594
rect 23204 23530 23256 23536
rect 23216 20466 23244 23530
rect 23400 22506 23428 23598
rect 23492 22574 23520 23666
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23584 23186 23612 23462
rect 23572 23180 23624 23186
rect 23572 23122 23624 23128
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23388 22500 23440 22506
rect 23388 22442 23440 22448
rect 23400 21978 23428 22442
rect 23664 22024 23716 22030
rect 23400 21972 23664 21978
rect 23400 21966 23716 21972
rect 23400 21950 23704 21966
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23308 21690 23336 21830
rect 23296 21684 23348 21690
rect 23296 21626 23348 21632
rect 23400 21486 23428 21950
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 20874 23704 21286
rect 23664 20868 23716 20874
rect 23664 20810 23716 20816
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 23216 19718 23244 20402
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23400 20058 23428 20198
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23584 17610 23612 18566
rect 23572 17604 23624 17610
rect 23572 17546 23624 17552
rect 23768 12434 23796 24534
rect 23848 23656 23900 23662
rect 23848 23598 23900 23604
rect 23860 22642 23888 23598
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23860 22166 23888 22578
rect 23848 22160 23900 22166
rect 23848 22102 23900 22108
rect 23952 21894 23980 22578
rect 23940 21888 23992 21894
rect 23940 21830 23992 21836
rect 23952 20806 23980 21830
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 24044 19310 24072 25706
rect 24872 25226 24900 26998
rect 24964 26586 24992 29106
rect 25056 26874 25084 32150
rect 25516 32065 25544 32370
rect 25502 32056 25558 32065
rect 25502 31991 25558 32000
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25136 30048 25188 30054
rect 25136 29990 25188 29996
rect 25148 29578 25176 29990
rect 25136 29572 25188 29578
rect 25136 29514 25188 29520
rect 25056 26846 25176 26874
rect 24952 26580 25004 26586
rect 24952 26522 25004 26528
rect 24860 25220 24912 25226
rect 24860 25162 24912 25168
rect 24492 24880 24544 24886
rect 24492 24822 24544 24828
rect 24504 24410 24532 24822
rect 24492 24404 24544 24410
rect 24492 24346 24544 24352
rect 24124 23180 24176 23186
rect 24124 23122 24176 23128
rect 24136 22778 24164 23122
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 24676 21956 24728 21962
rect 24676 21898 24728 21904
rect 24860 21956 24912 21962
rect 24860 21898 24912 21904
rect 24688 21554 24716 21898
rect 24872 21690 24900 21898
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24584 20324 24636 20330
rect 24584 20266 24636 20272
rect 24596 19922 24624 20266
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 24596 19378 24624 19858
rect 24584 19372 24636 19378
rect 24584 19314 24636 19320
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 24044 17882 24072 19246
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24504 18358 24532 18566
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24596 12434 24624 19314
rect 23768 12406 23888 12434
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23584 4146 23612 4558
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23112 4004 23164 4010
rect 23112 3946 23164 3952
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 23216 800 23244 4014
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 23400 3398 23428 3674
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23492 2650 23520 4082
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 23676 2446 23704 3334
rect 23860 2650 23888 12406
rect 24412 12406 24624 12434
rect 24412 4078 24440 12406
rect 24964 8430 24992 26522
rect 25044 24812 25096 24818
rect 25044 24754 25096 24760
rect 25056 24206 25084 24754
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 25056 20330 25084 24142
rect 25044 20324 25096 20330
rect 25044 20266 25096 20272
rect 25056 18766 25084 20266
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 25148 12434 25176 26846
rect 25240 24750 25268 31758
rect 25608 31754 25636 32438
rect 25792 32298 25820 34886
rect 25976 34678 26004 35090
rect 25964 34672 26016 34678
rect 25964 34614 26016 34620
rect 26160 34610 26188 37606
rect 26148 34604 26200 34610
rect 26148 34546 26200 34552
rect 26160 34406 26188 34546
rect 26148 34400 26200 34406
rect 26148 34342 26200 34348
rect 26148 33856 26200 33862
rect 26148 33798 26200 33804
rect 26160 33658 26188 33798
rect 26344 33658 26372 37674
rect 26516 37188 26568 37194
rect 26516 37130 26568 37136
rect 26424 36236 26476 36242
rect 26424 36178 26476 36184
rect 26436 35290 26464 36178
rect 26424 35284 26476 35290
rect 26424 35226 26476 35232
rect 26528 33930 26556 37130
rect 26516 33924 26568 33930
rect 26516 33866 26568 33872
rect 26148 33652 26200 33658
rect 26148 33594 26200 33600
rect 26332 33652 26384 33658
rect 26332 33594 26384 33600
rect 25872 33516 25924 33522
rect 25872 33458 25924 33464
rect 25780 32292 25832 32298
rect 25780 32234 25832 32240
rect 25596 31748 25648 31754
rect 25596 31690 25648 31696
rect 25412 31340 25464 31346
rect 25412 31282 25464 31288
rect 25424 30734 25452 31282
rect 25504 31204 25556 31210
rect 25504 31146 25556 31152
rect 25412 30728 25464 30734
rect 25412 30670 25464 30676
rect 25516 30258 25544 31146
rect 25504 30252 25556 30258
rect 25504 30194 25556 30200
rect 25608 28150 25636 31690
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 25688 30116 25740 30122
rect 25688 30058 25740 30064
rect 25700 29782 25728 30058
rect 25688 29776 25740 29782
rect 25688 29718 25740 29724
rect 25596 28144 25648 28150
rect 25596 28086 25648 28092
rect 25608 27606 25636 28086
rect 25596 27600 25648 27606
rect 25596 27542 25648 27548
rect 25700 27334 25728 29718
rect 25688 27328 25740 27334
rect 25688 27270 25740 27276
rect 25792 26994 25820 30194
rect 25884 28150 25912 33458
rect 26148 33312 26200 33318
rect 26148 33254 26200 33260
rect 26160 32502 26188 33254
rect 26344 33114 26372 33594
rect 26528 33504 26556 33866
rect 26436 33476 26556 33504
rect 26332 33108 26384 33114
rect 26332 33050 26384 33056
rect 26436 33046 26464 33476
rect 26516 33312 26568 33318
rect 26516 33254 26568 33260
rect 26424 33040 26476 33046
rect 26424 32982 26476 32988
rect 26528 32910 26556 33254
rect 26516 32904 26568 32910
rect 26516 32846 26568 32852
rect 26148 32496 26200 32502
rect 26148 32438 26200 32444
rect 26424 32360 26476 32366
rect 26422 32328 26424 32337
rect 26476 32328 26478 32337
rect 26422 32263 26478 32272
rect 26516 32020 26568 32026
rect 26516 31962 26568 31968
rect 26528 31822 26556 31962
rect 26516 31816 26568 31822
rect 26516 31758 26568 31764
rect 26148 31748 26200 31754
rect 26148 31690 26200 31696
rect 26160 31346 26188 31690
rect 26148 31340 26200 31346
rect 26148 31282 26200 31288
rect 26240 30728 26292 30734
rect 26240 30670 26292 30676
rect 26252 30326 26280 30670
rect 26240 30320 26292 30326
rect 26240 30262 26292 30268
rect 25964 29028 26016 29034
rect 25964 28970 26016 28976
rect 25976 28626 26004 28970
rect 25964 28620 26016 28626
rect 25964 28562 26016 28568
rect 25976 28150 26004 28562
rect 25872 28144 25924 28150
rect 25872 28086 25924 28092
rect 25964 28144 26016 28150
rect 25964 28086 26016 28092
rect 25872 27328 25924 27334
rect 25872 27270 25924 27276
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25332 26450 25360 26862
rect 25688 26784 25740 26790
rect 25688 26726 25740 26732
rect 25320 26444 25372 26450
rect 25320 26386 25372 26392
rect 25332 24954 25360 26386
rect 25700 26382 25728 26726
rect 25792 26382 25820 26930
rect 25688 26376 25740 26382
rect 25688 26318 25740 26324
rect 25780 26376 25832 26382
rect 25780 26318 25832 26324
rect 25884 26314 25912 27270
rect 26620 26586 26648 41386
rect 26608 26580 26660 26586
rect 26608 26522 26660 26528
rect 25872 26308 25924 26314
rect 25872 26250 25924 26256
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 26252 25362 26280 26182
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25412 25152 25464 25158
rect 25412 25094 25464 25100
rect 25320 24948 25372 24954
rect 25320 24890 25372 24896
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25424 24138 25452 25094
rect 25412 24132 25464 24138
rect 25412 24074 25464 24080
rect 25228 22432 25280 22438
rect 25228 22374 25280 22380
rect 25240 21554 25268 22374
rect 25228 21548 25280 21554
rect 25228 21490 25280 21496
rect 25608 12782 25636 25230
rect 26424 24608 26476 24614
rect 26424 24550 26476 24556
rect 26436 24138 26464 24550
rect 26424 24132 26476 24138
rect 26424 24074 26476 24080
rect 26424 23656 26476 23662
rect 26424 23598 26476 23604
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25700 22098 25728 22374
rect 25688 22092 25740 22098
rect 25688 22034 25740 22040
rect 25976 21418 26004 22578
rect 26240 22432 26292 22438
rect 26240 22374 26292 22380
rect 26252 22234 26280 22374
rect 26436 22234 26464 23598
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26424 22228 26476 22234
rect 26424 22170 26476 22176
rect 26240 21956 26292 21962
rect 26240 21898 26292 21904
rect 26252 21690 26280 21898
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 25964 21412 26016 21418
rect 25964 21354 26016 21360
rect 25976 20942 26004 21354
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 25976 19854 26004 20334
rect 26056 19916 26108 19922
rect 26056 19858 26108 19864
rect 25964 19848 26016 19854
rect 25964 19790 26016 19796
rect 25976 19378 26004 19790
rect 25964 19372 26016 19378
rect 25964 19314 26016 19320
rect 26068 18766 26096 19858
rect 26252 19718 26280 20402
rect 26712 20330 26740 42094
rect 26988 39914 27016 43182
rect 26976 39908 27028 39914
rect 26976 39850 27028 39856
rect 26976 38956 27028 38962
rect 26976 38898 27028 38904
rect 26988 38554 27016 38898
rect 26976 38548 27028 38554
rect 26976 38490 27028 38496
rect 26884 37868 26936 37874
rect 26884 37810 26936 37816
rect 26896 37194 26924 37810
rect 27528 37800 27580 37806
rect 27528 37742 27580 37748
rect 27160 37664 27212 37670
rect 27160 37606 27212 37612
rect 27172 37330 27200 37606
rect 27160 37324 27212 37330
rect 27160 37266 27212 37272
rect 26884 37188 26936 37194
rect 26884 37130 26936 37136
rect 26976 37120 27028 37126
rect 26976 37062 27028 37068
rect 26988 36650 27016 37062
rect 26976 36644 27028 36650
rect 26976 36586 27028 36592
rect 26988 35698 27016 36586
rect 27068 36100 27120 36106
rect 27068 36042 27120 36048
rect 27080 35834 27108 36042
rect 27160 36032 27212 36038
rect 27160 35974 27212 35980
rect 27068 35828 27120 35834
rect 27068 35770 27120 35776
rect 26976 35692 27028 35698
rect 26896 35652 26976 35680
rect 26792 33992 26844 33998
rect 26792 33934 26844 33940
rect 26804 33114 26832 33934
rect 26896 33454 26924 35652
rect 26976 35634 27028 35640
rect 27172 35290 27200 35974
rect 27160 35284 27212 35290
rect 27160 35226 27212 35232
rect 27068 35216 27120 35222
rect 27068 35158 27120 35164
rect 26976 33584 27028 33590
rect 26976 33526 27028 33532
rect 26884 33448 26936 33454
rect 26884 33390 26936 33396
rect 26792 33108 26844 33114
rect 26792 33050 26844 33056
rect 26988 32434 27016 33526
rect 26976 32428 27028 32434
rect 26976 32370 27028 32376
rect 26792 32292 26844 32298
rect 26792 32234 26844 32240
rect 26804 32026 26832 32234
rect 26792 32020 26844 32026
rect 26792 31962 26844 31968
rect 26976 30932 27028 30938
rect 26976 30874 27028 30880
rect 26792 30728 26844 30734
rect 26792 30670 26844 30676
rect 26804 28762 26832 30670
rect 26988 30054 27016 30874
rect 27080 30054 27108 35158
rect 27172 35154 27200 35226
rect 27160 35148 27212 35154
rect 27160 35090 27212 35096
rect 27344 35148 27396 35154
rect 27344 35090 27396 35096
rect 27172 34610 27200 35090
rect 27252 35012 27304 35018
rect 27252 34954 27304 34960
rect 27160 34604 27212 34610
rect 27160 34546 27212 34552
rect 27160 34400 27212 34406
rect 27160 34342 27212 34348
rect 27172 33810 27200 34342
rect 27264 33998 27292 34954
rect 27356 34678 27384 35090
rect 27540 35086 27568 37742
rect 27620 35624 27672 35630
rect 27620 35566 27672 35572
rect 27436 35080 27488 35086
rect 27436 35022 27488 35028
rect 27528 35080 27580 35086
rect 27528 35022 27580 35028
rect 27448 34746 27476 35022
rect 27436 34740 27488 34746
rect 27436 34682 27488 34688
rect 27632 34678 27660 35566
rect 27344 34672 27396 34678
rect 27344 34614 27396 34620
rect 27620 34672 27672 34678
rect 27620 34614 27672 34620
rect 27436 34400 27488 34406
rect 27436 34342 27488 34348
rect 27448 34066 27476 34342
rect 27436 34060 27488 34066
rect 27436 34002 27488 34008
rect 27252 33992 27304 33998
rect 27252 33934 27304 33940
rect 27172 33782 27292 33810
rect 27160 33516 27212 33522
rect 27160 33458 27212 33464
rect 27172 32842 27200 33458
rect 27160 32836 27212 32842
rect 27160 32778 27212 32784
rect 27172 32434 27200 32778
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 27172 32298 27200 32370
rect 27160 32292 27212 32298
rect 27160 32234 27212 32240
rect 27160 30660 27212 30666
rect 27160 30602 27212 30608
rect 26976 30048 27028 30054
rect 26976 29990 27028 29996
rect 27068 30048 27120 30054
rect 27068 29990 27120 29996
rect 27080 29646 27108 29990
rect 27068 29640 27120 29646
rect 27068 29582 27120 29588
rect 27172 29102 27200 30602
rect 27264 29850 27292 33782
rect 27448 33590 27476 34002
rect 27620 33992 27672 33998
rect 27620 33934 27672 33940
rect 27528 33924 27580 33930
rect 27528 33866 27580 33872
rect 27436 33584 27488 33590
rect 27436 33526 27488 33532
rect 27540 33318 27568 33866
rect 27528 33312 27580 33318
rect 27528 33254 27580 33260
rect 27632 32994 27660 33934
rect 27540 32966 27660 32994
rect 27540 32502 27568 32966
rect 27620 32836 27672 32842
rect 27620 32778 27672 32784
rect 27632 32570 27660 32778
rect 27620 32564 27672 32570
rect 27620 32506 27672 32512
rect 27528 32496 27580 32502
rect 27528 32438 27580 32444
rect 27724 31754 27752 44270
rect 28816 43240 28868 43246
rect 28816 43182 28868 43188
rect 28828 42158 28856 43182
rect 28816 42152 28868 42158
rect 28816 42094 28868 42100
rect 28172 37800 28224 37806
rect 28172 37742 28224 37748
rect 28184 36786 28212 37742
rect 28264 37664 28316 37670
rect 28316 37624 28396 37652
rect 28264 37606 28316 37612
rect 28368 37262 28396 37624
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 28724 37256 28776 37262
rect 28724 37198 28776 37204
rect 28172 36780 28224 36786
rect 28172 36722 28224 36728
rect 27896 36100 27948 36106
rect 27896 36042 27948 36048
rect 27804 35692 27856 35698
rect 27804 35634 27856 35640
rect 27816 35562 27844 35634
rect 27804 35556 27856 35562
rect 27804 35498 27856 35504
rect 27816 35222 27844 35498
rect 27804 35216 27856 35222
rect 27804 35158 27856 35164
rect 27908 35068 27936 36042
rect 28080 36032 28132 36038
rect 28080 35974 28132 35980
rect 27988 35692 28040 35698
rect 28092 35680 28120 35974
rect 28264 35760 28316 35766
rect 28264 35702 28316 35708
rect 28040 35652 28120 35680
rect 27988 35634 28040 35640
rect 28276 35442 28304 35702
rect 27816 35040 27936 35068
rect 28000 35414 28304 35442
rect 27816 34202 27844 35040
rect 27896 34604 27948 34610
rect 27896 34546 27948 34552
rect 27908 34406 27936 34546
rect 27896 34400 27948 34406
rect 27896 34342 27948 34348
rect 27804 34196 27856 34202
rect 27804 34138 27856 34144
rect 27896 34060 27948 34066
rect 28000 34048 28028 35414
rect 28368 35329 28396 37198
rect 28540 36780 28592 36786
rect 28540 36722 28592 36728
rect 28354 35320 28410 35329
rect 28264 35284 28316 35290
rect 28354 35255 28410 35264
rect 28264 35226 28316 35232
rect 28080 34128 28132 34134
rect 28080 34070 28132 34076
rect 27948 34020 28028 34048
rect 27896 34002 27948 34008
rect 27908 32502 27936 34002
rect 27988 33856 28040 33862
rect 27988 33798 28040 33804
rect 27896 32496 27948 32502
rect 27896 32438 27948 32444
rect 27804 32428 27856 32434
rect 27804 32370 27856 32376
rect 27528 31748 27580 31754
rect 27528 31690 27580 31696
rect 27632 31726 27752 31754
rect 27540 30666 27568 31690
rect 27528 30660 27580 30666
rect 27528 30602 27580 30608
rect 27436 30252 27488 30258
rect 27436 30194 27488 30200
rect 27252 29844 27304 29850
rect 27252 29786 27304 29792
rect 27160 29096 27212 29102
rect 27160 29038 27212 29044
rect 26792 28756 26844 28762
rect 26792 28698 26844 28704
rect 26804 28082 26832 28698
rect 26792 28076 26844 28082
rect 26792 28018 26844 28024
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 27080 27674 27108 27814
rect 27068 27668 27120 27674
rect 27068 27610 27120 27616
rect 26792 27464 26844 27470
rect 26976 27464 27028 27470
rect 26792 27406 26844 27412
rect 26896 27424 26976 27452
rect 26804 27062 26832 27406
rect 26792 27056 26844 27062
rect 26792 26998 26844 27004
rect 26896 26994 26924 27424
rect 26976 27406 27028 27412
rect 26884 26988 26936 26994
rect 26884 26930 26936 26936
rect 26976 26988 27028 26994
rect 26976 26930 27028 26936
rect 26896 26790 26924 26930
rect 26884 26784 26936 26790
rect 26884 26726 26936 26732
rect 26896 26314 26924 26726
rect 26988 26450 27016 26930
rect 27172 26518 27200 29038
rect 27448 28490 27476 30194
rect 27436 28484 27488 28490
rect 27436 28426 27488 28432
rect 27344 28076 27396 28082
rect 27344 28018 27396 28024
rect 27252 27532 27304 27538
rect 27252 27474 27304 27480
rect 27264 26858 27292 27474
rect 27252 26852 27304 26858
rect 27252 26794 27304 26800
rect 27160 26512 27212 26518
rect 27160 26454 27212 26460
rect 26976 26444 27028 26450
rect 26976 26386 27028 26392
rect 26884 26308 26936 26314
rect 26884 26250 26936 26256
rect 26896 24342 26924 26250
rect 26988 25974 27016 26386
rect 27264 26382 27292 26794
rect 27252 26376 27304 26382
rect 27252 26318 27304 26324
rect 27264 25974 27292 26318
rect 26976 25968 27028 25974
rect 26976 25910 27028 25916
rect 27252 25968 27304 25974
rect 27252 25910 27304 25916
rect 27252 25288 27304 25294
rect 27356 25276 27384 28018
rect 27448 26858 27476 28426
rect 27436 26852 27488 26858
rect 27436 26794 27488 26800
rect 27436 26512 27488 26518
rect 27436 26454 27488 26460
rect 27448 26382 27476 26454
rect 27436 26376 27488 26382
rect 27436 26318 27488 26324
rect 27528 25696 27580 25702
rect 27528 25638 27580 25644
rect 27304 25248 27384 25276
rect 27252 25230 27304 25236
rect 26884 24336 26936 24342
rect 26884 24278 26936 24284
rect 27264 24274 27292 25230
rect 27540 25226 27568 25638
rect 27528 25220 27580 25226
rect 27528 25162 27580 25168
rect 27252 24268 27304 24274
rect 27252 24210 27304 24216
rect 26884 22024 26936 22030
rect 26884 21966 26936 21972
rect 26896 21078 26924 21966
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27356 21554 27384 21830
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 26884 21072 26936 21078
rect 26884 21014 26936 21020
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 26700 20324 26752 20330
rect 26700 20266 26752 20272
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 26516 19984 26568 19990
rect 26516 19926 26568 19932
rect 26424 19848 26476 19854
rect 26424 19790 26476 19796
rect 26240 19712 26292 19718
rect 26240 19654 26292 19660
rect 26436 19378 26464 19790
rect 26528 19514 26556 19926
rect 27356 19854 27384 20198
rect 27448 20058 27476 20402
rect 27436 20052 27488 20058
rect 27436 19994 27488 20000
rect 26608 19848 26660 19854
rect 26608 19790 26660 19796
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27344 19848 27396 19854
rect 27344 19790 27396 19796
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 26620 19514 26648 19790
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 26056 18760 26108 18766
rect 26056 18702 26108 18708
rect 26068 18290 26096 18702
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26252 18290 26280 18566
rect 26620 18358 26648 19450
rect 27172 19378 27200 19790
rect 27344 19712 27396 19718
rect 27344 19654 27396 19660
rect 27356 19514 27384 19654
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 27540 19446 27568 19790
rect 27528 19440 27580 19446
rect 27528 19382 27580 19388
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 26988 19258 27016 19314
rect 26988 19230 27108 19258
rect 26884 19168 26936 19174
rect 26884 19110 26936 19116
rect 26896 18766 26924 19110
rect 26884 18760 26936 18766
rect 26884 18702 26936 18708
rect 26896 18358 26924 18702
rect 26608 18352 26660 18358
rect 26608 18294 26660 18300
rect 26884 18352 26936 18358
rect 26884 18294 26936 18300
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 26068 17610 26096 18226
rect 26252 17610 26280 18226
rect 26424 18216 26476 18222
rect 26424 18158 26476 18164
rect 26436 17882 26464 18158
rect 26424 17876 26476 17882
rect 26424 17818 26476 17824
rect 25688 17604 25740 17610
rect 25688 17546 25740 17552
rect 26056 17604 26108 17610
rect 26056 17546 26108 17552
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 25596 12776 25648 12782
rect 25596 12718 25648 12724
rect 25056 12406 25176 12434
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24400 4072 24452 4078
rect 24400 4014 24452 4020
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 24412 2582 24440 4014
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 24584 3460 24636 3466
rect 24584 3402 24636 3408
rect 24596 3058 24624 3402
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24400 2576 24452 2582
rect 24400 2518 24452 2524
rect 24688 2514 24716 3878
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24780 3126 24808 3334
rect 24768 3120 24820 3126
rect 24768 3062 24820 3068
rect 24872 2961 24900 3334
rect 24858 2952 24914 2961
rect 24858 2887 24914 2896
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24504 800 24532 2246
rect 25056 2106 25084 12406
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 25044 2100 25096 2106
rect 25044 2042 25096 2048
rect 25148 800 25176 2926
rect 25412 2576 25464 2582
rect 25412 2518 25464 2524
rect 25424 2428 25452 2518
rect 25700 2514 25728 17546
rect 26252 4146 26280 17546
rect 27080 12434 27108 19230
rect 27172 18970 27200 19314
rect 27160 18964 27212 18970
rect 27160 18906 27212 18912
rect 27632 18766 27660 31726
rect 27816 31482 27844 32370
rect 27908 31958 27936 32438
rect 28000 32434 28028 33798
rect 27988 32428 28040 32434
rect 27988 32370 28040 32376
rect 27896 31952 27948 31958
rect 27896 31894 27948 31900
rect 28092 31754 28120 34070
rect 28172 33108 28224 33114
rect 28172 33050 28224 33056
rect 28184 32298 28212 33050
rect 28276 32366 28304 35226
rect 28552 35154 28580 36722
rect 28736 36106 28764 37198
rect 28724 36100 28776 36106
rect 28724 36042 28776 36048
rect 28828 35737 28856 42094
rect 28908 37800 28960 37806
rect 28908 37742 28960 37748
rect 28920 37466 28948 37742
rect 28908 37460 28960 37466
rect 28908 37402 28960 37408
rect 29184 37188 29236 37194
rect 29184 37130 29236 37136
rect 29000 36032 29052 36038
rect 29000 35974 29052 35980
rect 29012 35737 29040 35974
rect 29090 35864 29146 35873
rect 29090 35799 29146 35808
rect 29104 35766 29132 35799
rect 29092 35760 29144 35766
rect 28814 35728 28870 35737
rect 28814 35663 28870 35672
rect 28998 35728 29054 35737
rect 29092 35702 29144 35708
rect 28998 35663 29000 35672
rect 29052 35663 29054 35672
rect 29000 35634 29052 35640
rect 29090 35592 29146 35601
rect 29090 35527 29146 35536
rect 29104 35494 29132 35527
rect 29092 35488 29144 35494
rect 28814 35456 28870 35465
rect 29092 35430 29144 35436
rect 28814 35391 28870 35400
rect 28722 35320 28778 35329
rect 28722 35255 28778 35264
rect 28540 35148 28592 35154
rect 28540 35090 28592 35096
rect 28356 34604 28408 34610
rect 28356 34546 28408 34552
rect 28368 34474 28396 34546
rect 28356 34468 28408 34474
rect 28356 34410 28408 34416
rect 28368 34134 28396 34410
rect 28356 34128 28408 34134
rect 28356 34070 28408 34076
rect 28552 33658 28580 35090
rect 28632 34944 28684 34950
rect 28632 34886 28684 34892
rect 28644 34610 28672 34886
rect 28632 34604 28684 34610
rect 28632 34546 28684 34552
rect 28540 33652 28592 33658
rect 28540 33594 28592 33600
rect 28448 33516 28500 33522
rect 28448 33458 28500 33464
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28172 32292 28224 32298
rect 28172 32234 28224 32240
rect 28000 31726 28120 31754
rect 27804 31476 27856 31482
rect 27804 31418 27856 31424
rect 28000 31346 28028 31726
rect 28184 31346 28212 32234
rect 27988 31340 28040 31346
rect 27988 31282 28040 31288
rect 28172 31340 28224 31346
rect 28172 31282 28224 31288
rect 27712 29504 27764 29510
rect 27712 29446 27764 29452
rect 27804 29504 27856 29510
rect 27804 29446 27856 29452
rect 27724 29102 27752 29446
rect 27816 29170 27844 29446
rect 27804 29164 27856 29170
rect 27804 29106 27856 29112
rect 27712 29096 27764 29102
rect 27712 29038 27764 29044
rect 27724 28966 27752 29038
rect 27896 29028 27948 29034
rect 27896 28970 27948 28976
rect 27712 28960 27764 28966
rect 27712 28902 27764 28908
rect 27908 28558 27936 28970
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 27896 28008 27948 28014
rect 27896 27950 27948 27956
rect 27712 22092 27764 22098
rect 27712 22034 27764 22040
rect 27724 21486 27752 22034
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27908 20534 27936 27950
rect 28000 27402 28028 31282
rect 28276 30870 28304 32302
rect 28460 31958 28488 33458
rect 28552 32978 28580 33594
rect 28540 32972 28592 32978
rect 28540 32914 28592 32920
rect 28448 31952 28500 31958
rect 28448 31894 28500 31900
rect 28460 31754 28488 31894
rect 28460 31726 28580 31754
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28264 30864 28316 30870
rect 28264 30806 28316 30812
rect 28368 30274 28396 31282
rect 28276 30246 28396 30274
rect 28448 30252 28500 30258
rect 28080 29776 28132 29782
rect 28080 29718 28132 29724
rect 28092 29170 28120 29718
rect 28172 29640 28224 29646
rect 28172 29582 28224 29588
rect 28080 29164 28132 29170
rect 28080 29106 28132 29112
rect 28080 28688 28132 28694
rect 28080 28630 28132 28636
rect 27988 27396 28040 27402
rect 27988 27338 28040 27344
rect 27988 26240 28040 26246
rect 27988 26182 28040 26188
rect 28000 25906 28028 26182
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 28092 25344 28120 28630
rect 28184 28558 28212 29582
rect 28276 29034 28304 30246
rect 28448 30194 28500 30200
rect 28460 30138 28488 30194
rect 28368 30110 28488 30138
rect 28368 29646 28396 30110
rect 28448 29844 28500 29850
rect 28448 29786 28500 29792
rect 28356 29640 28408 29646
rect 28356 29582 28408 29588
rect 28460 29170 28488 29786
rect 28448 29164 28500 29170
rect 28448 29106 28500 29112
rect 28264 29028 28316 29034
rect 28264 28970 28316 28976
rect 28276 28642 28304 28970
rect 28276 28614 28396 28642
rect 28368 28558 28396 28614
rect 28552 28558 28580 31726
rect 28632 31136 28684 31142
rect 28632 31078 28684 31084
rect 28172 28552 28224 28558
rect 28172 28494 28224 28500
rect 28356 28552 28408 28558
rect 28356 28494 28408 28500
rect 28540 28552 28592 28558
rect 28540 28494 28592 28500
rect 28184 28218 28212 28494
rect 28172 28212 28224 28218
rect 28172 28154 28224 28160
rect 28368 27674 28396 28494
rect 28448 28416 28500 28422
rect 28448 28358 28500 28364
rect 28460 28082 28488 28358
rect 28448 28076 28500 28082
rect 28448 28018 28500 28024
rect 28356 27668 28408 27674
rect 28356 27610 28408 27616
rect 28172 27396 28224 27402
rect 28172 27338 28224 27344
rect 28184 25906 28212 27338
rect 28368 27062 28396 27610
rect 28356 27056 28408 27062
rect 28356 26998 28408 27004
rect 28264 26920 28316 26926
rect 28264 26862 28316 26868
rect 28276 26382 28304 26862
rect 28264 26376 28316 26382
rect 28264 26318 28316 26324
rect 28172 25900 28224 25906
rect 28172 25842 28224 25848
rect 28276 25838 28304 26318
rect 28368 25974 28396 26998
rect 28356 25968 28408 25974
rect 28356 25910 28408 25916
rect 28264 25832 28316 25838
rect 28264 25774 28316 25780
rect 28356 25832 28408 25838
rect 28356 25774 28408 25780
rect 28276 25498 28304 25774
rect 28264 25492 28316 25498
rect 28264 25434 28316 25440
rect 28000 25316 28120 25344
rect 27896 20528 27948 20534
rect 27896 20470 27948 20476
rect 27712 20460 27764 20466
rect 27712 20402 27764 20408
rect 27724 19990 27752 20402
rect 27712 19984 27764 19990
rect 27712 19926 27764 19932
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27172 18358 27200 18702
rect 27804 18692 27856 18698
rect 27804 18634 27856 18640
rect 27160 18352 27212 18358
rect 27160 18294 27212 18300
rect 27816 18222 27844 18634
rect 27804 18216 27856 18222
rect 27804 18158 27856 18164
rect 27436 18148 27488 18154
rect 27436 18090 27488 18096
rect 27448 17678 27476 18090
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27712 17604 27764 17610
rect 27712 17546 27764 17552
rect 27724 17134 27752 17546
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 27080 12406 27200 12434
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 26884 4004 26936 4010
rect 26884 3946 26936 3952
rect 26896 2854 26924 3946
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 26884 2848 26936 2854
rect 26884 2790 26936 2796
rect 25688 2508 25740 2514
rect 25688 2450 25740 2456
rect 25596 2440 25648 2446
rect 25424 2400 25596 2428
rect 25596 2382 25648 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26436 800 26464 2382
rect 27080 800 27108 2994
rect 27172 2514 27200 12406
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27632 2854 27660 11630
rect 27724 5710 27752 17070
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 28000 3126 28028 25316
rect 28080 25220 28132 25226
rect 28080 25162 28132 25168
rect 28092 24818 28120 25162
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28264 22024 28316 22030
rect 28264 21966 28316 21972
rect 28276 21690 28304 21966
rect 28368 21690 28396 25774
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28552 22778 28580 23054
rect 28540 22772 28592 22778
rect 28540 22714 28592 22720
rect 28540 22636 28592 22642
rect 28540 22578 28592 22584
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 28356 21684 28408 21690
rect 28356 21626 28408 21632
rect 28552 20602 28580 22578
rect 28540 20596 28592 20602
rect 28540 20538 28592 20544
rect 28080 18692 28132 18698
rect 28080 18634 28132 18640
rect 28092 18426 28120 18634
rect 28080 18420 28132 18426
rect 28080 18362 28132 18368
rect 28080 18216 28132 18222
rect 28080 18158 28132 18164
rect 28092 17678 28120 18158
rect 28080 17672 28132 17678
rect 28080 17614 28132 17620
rect 28172 17128 28224 17134
rect 28172 17070 28224 17076
rect 28184 16794 28212 17070
rect 28172 16788 28224 16794
rect 28172 16730 28224 16736
rect 28540 4072 28592 4078
rect 28540 4014 28592 4020
rect 28552 3738 28580 4014
rect 28540 3732 28592 3738
rect 28540 3674 28592 3680
rect 27988 3120 28040 3126
rect 27988 3062 28040 3068
rect 27620 2848 27672 2854
rect 27620 2790 27672 2796
rect 28644 2650 28672 31078
rect 28736 29238 28764 35255
rect 28724 29232 28776 29238
rect 28724 29174 28776 29180
rect 28736 28762 28764 29174
rect 28724 28756 28776 28762
rect 28724 28698 28776 28704
rect 28724 28416 28776 28422
rect 28724 28358 28776 28364
rect 28736 28150 28764 28358
rect 28724 28144 28776 28150
rect 28724 28086 28776 28092
rect 28828 28014 28856 35391
rect 29196 35290 29224 37130
rect 29274 35864 29330 35873
rect 29274 35799 29330 35808
rect 29184 35284 29236 35290
rect 29184 35226 29236 35232
rect 29000 34400 29052 34406
rect 29000 34342 29052 34348
rect 28908 32904 28960 32910
rect 28908 32846 28960 32852
rect 28920 32230 28948 32846
rect 28908 32224 28960 32230
rect 28908 32166 28960 32172
rect 28816 28008 28868 28014
rect 28816 27950 28868 27956
rect 28920 27470 28948 32166
rect 29012 31686 29040 34342
rect 29184 33312 29236 33318
rect 29184 33254 29236 33260
rect 29196 32842 29224 33254
rect 29184 32836 29236 32842
rect 29184 32778 29236 32784
rect 29092 32292 29144 32298
rect 29092 32234 29144 32240
rect 29000 31680 29052 31686
rect 29000 31622 29052 31628
rect 29000 30592 29052 30598
rect 29000 30534 29052 30540
rect 29012 29646 29040 30534
rect 29000 29640 29052 29646
rect 29000 29582 29052 29588
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28724 23724 28776 23730
rect 28724 23666 28776 23672
rect 28736 22642 28764 23666
rect 28920 23594 28948 27406
rect 28908 23588 28960 23594
rect 28908 23530 28960 23536
rect 28724 22636 28776 22642
rect 28724 22578 28776 22584
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28724 18080 28776 18086
rect 28724 18022 28776 18028
rect 28736 17270 28764 18022
rect 28724 17264 28776 17270
rect 28724 17206 28776 17212
rect 28828 16046 28856 19790
rect 29012 18154 29040 19790
rect 29000 18148 29052 18154
rect 29000 18090 29052 18096
rect 28816 16040 28868 16046
rect 28816 15982 28868 15988
rect 29104 2922 29132 32234
rect 29288 30938 29316 35799
rect 29276 30932 29328 30938
rect 29276 30874 29328 30880
rect 29276 30796 29328 30802
rect 29276 30738 29328 30744
rect 29184 30660 29236 30666
rect 29184 30602 29236 30608
rect 29196 30258 29224 30602
rect 29184 30252 29236 30258
rect 29184 30194 29236 30200
rect 29288 30054 29316 30738
rect 29276 30048 29328 30054
rect 29276 29990 29328 29996
rect 29276 24744 29328 24750
rect 29276 24686 29328 24692
rect 29184 24200 29236 24206
rect 29184 24142 29236 24148
rect 29196 19922 29224 24142
rect 29288 22642 29316 24686
rect 29276 22636 29328 22642
rect 29276 22578 29328 22584
rect 29184 19916 29236 19922
rect 29184 19858 29236 19864
rect 29380 19514 29408 47194
rect 29656 47054 29684 49200
rect 30760 47122 30788 49286
rect 30902 49200 31014 49286
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49200 40030 50000
rect 40562 49200 40674 50000
rect 41206 49200 41318 50000
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49314 43250 50000
rect 43138 49286 43668 49314
rect 43138 49200 43250 49286
rect 30748 47116 30800 47122
rect 30748 47058 30800 47064
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 31116 47048 31168 47054
rect 31116 46990 31168 46996
rect 29552 44872 29604 44878
rect 29552 44814 29604 44820
rect 29564 44198 29592 44814
rect 29552 44192 29604 44198
rect 29552 44134 29604 44140
rect 29564 43790 29592 44134
rect 29552 43784 29604 43790
rect 29552 43726 29604 43732
rect 30196 38956 30248 38962
rect 30196 38898 30248 38904
rect 29552 37868 29604 37874
rect 29552 37810 29604 37816
rect 29564 37466 29592 37810
rect 29920 37664 29972 37670
rect 29920 37606 29972 37612
rect 29552 37460 29604 37466
rect 29552 37402 29604 37408
rect 29932 37330 29960 37606
rect 29736 37324 29788 37330
rect 29736 37266 29788 37272
rect 29920 37324 29972 37330
rect 29920 37266 29972 37272
rect 29460 36712 29512 36718
rect 29460 36654 29512 36660
rect 29472 35834 29500 36654
rect 29748 36174 29776 37266
rect 29736 36168 29788 36174
rect 29736 36110 29788 36116
rect 29920 36168 29972 36174
rect 29920 36110 29972 36116
rect 30012 36168 30064 36174
rect 30012 36110 30064 36116
rect 29644 36100 29696 36106
rect 29644 36042 29696 36048
rect 29460 35828 29512 35834
rect 29460 35770 29512 35776
rect 29552 35828 29604 35834
rect 29552 35770 29604 35776
rect 29460 35624 29512 35630
rect 29564 35601 29592 35770
rect 29656 35766 29684 36042
rect 29644 35760 29696 35766
rect 29644 35702 29696 35708
rect 29748 35630 29776 36110
rect 29828 36032 29880 36038
rect 29828 35974 29880 35980
rect 29736 35624 29788 35630
rect 29460 35566 29512 35572
rect 29550 35592 29606 35601
rect 29472 32298 29500 35566
rect 29550 35527 29606 35536
rect 29656 35584 29736 35612
rect 29656 35290 29684 35584
rect 29736 35566 29788 35572
rect 29736 35488 29788 35494
rect 29736 35430 29788 35436
rect 29644 35284 29696 35290
rect 29644 35226 29696 35232
rect 29748 35154 29776 35430
rect 29736 35148 29788 35154
rect 29736 35090 29788 35096
rect 29644 35080 29696 35086
rect 29840 35034 29868 35974
rect 29932 35698 29960 36110
rect 29920 35692 29972 35698
rect 29920 35634 29972 35640
rect 30024 35494 30052 36110
rect 30012 35488 30064 35494
rect 30012 35430 30064 35436
rect 29696 35028 29868 35034
rect 29644 35022 29868 35028
rect 29656 35006 29868 35022
rect 30104 35012 30156 35018
rect 30104 34954 30156 34960
rect 30116 34610 30144 34954
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 30104 34604 30156 34610
rect 30104 34546 30156 34552
rect 29932 33998 29960 34546
rect 30116 33998 30144 34546
rect 29920 33992 29972 33998
rect 29920 33934 29972 33940
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30116 33454 30144 33934
rect 30104 33448 30156 33454
rect 30104 33390 30156 33396
rect 30104 33108 30156 33114
rect 30104 33050 30156 33056
rect 30116 32774 30144 33050
rect 30104 32768 30156 32774
rect 30104 32710 30156 32716
rect 29460 32292 29512 32298
rect 29460 32234 29512 32240
rect 30104 31884 30156 31890
rect 30104 31826 30156 31832
rect 29552 31748 29604 31754
rect 29552 31690 29604 31696
rect 29460 31680 29512 31686
rect 29460 31622 29512 31628
rect 29472 31482 29500 31622
rect 29460 31476 29512 31482
rect 29460 31418 29512 31424
rect 29564 31346 29592 31690
rect 30116 31686 30144 31826
rect 30104 31680 30156 31686
rect 30104 31622 30156 31628
rect 29552 31340 29604 31346
rect 29552 31282 29604 31288
rect 29564 29578 29592 31282
rect 30116 31278 30144 31622
rect 30104 31272 30156 31278
rect 30104 31214 30156 31220
rect 29920 31204 29972 31210
rect 29920 31146 29972 31152
rect 29828 30864 29880 30870
rect 29828 30806 29880 30812
rect 29840 30734 29868 30806
rect 29828 30728 29880 30734
rect 29828 30670 29880 30676
rect 29840 30258 29868 30670
rect 29736 30252 29788 30258
rect 29736 30194 29788 30200
rect 29828 30252 29880 30258
rect 29828 30194 29880 30200
rect 29644 30184 29696 30190
rect 29644 30126 29696 30132
rect 29656 29782 29684 30126
rect 29644 29776 29696 29782
rect 29644 29718 29696 29724
rect 29552 29572 29604 29578
rect 29552 29514 29604 29520
rect 29748 29152 29776 30194
rect 29932 29850 29960 31146
rect 30012 31136 30064 31142
rect 30012 31078 30064 31084
rect 30024 30734 30052 31078
rect 30012 30728 30064 30734
rect 30012 30670 30064 30676
rect 29920 29844 29972 29850
rect 29920 29786 29972 29792
rect 29828 29164 29880 29170
rect 29748 29124 29828 29152
rect 29644 29096 29696 29102
rect 29748 29084 29776 29124
rect 29828 29106 29880 29112
rect 29696 29056 29776 29084
rect 29644 29038 29696 29044
rect 29736 28484 29788 28490
rect 29736 28426 29788 28432
rect 29460 27872 29512 27878
rect 29460 27814 29512 27820
rect 29472 27470 29500 27814
rect 29460 27464 29512 27470
rect 29460 27406 29512 27412
rect 29748 26994 29776 28426
rect 30012 27668 30064 27674
rect 30012 27610 30064 27616
rect 30024 27470 30052 27610
rect 30012 27464 30064 27470
rect 30012 27406 30064 27412
rect 29828 27328 29880 27334
rect 29828 27270 29880 27276
rect 30104 27328 30156 27334
rect 30104 27270 30156 27276
rect 29840 27130 29868 27270
rect 29828 27124 29880 27130
rect 29828 27066 29880 27072
rect 30116 27062 30144 27270
rect 30104 27056 30156 27062
rect 30104 26998 30156 27004
rect 29736 26988 29788 26994
rect 29736 26930 29788 26936
rect 29644 24744 29696 24750
rect 29644 24686 29696 24692
rect 29828 24744 29880 24750
rect 29828 24686 29880 24692
rect 29656 24342 29684 24686
rect 29644 24336 29696 24342
rect 29644 24278 29696 24284
rect 29840 23866 29868 24686
rect 30208 24206 30236 38898
rect 30748 37256 30800 37262
rect 30748 37198 30800 37204
rect 30760 36786 30788 37198
rect 30748 36780 30800 36786
rect 30748 36722 30800 36728
rect 30288 36576 30340 36582
rect 30288 36518 30340 36524
rect 30300 35737 30328 36518
rect 30286 35728 30342 35737
rect 30286 35663 30342 35672
rect 30932 35692 30984 35698
rect 30300 35086 30328 35663
rect 30932 35634 30984 35640
rect 30944 35494 30972 35634
rect 30932 35488 30984 35494
rect 30932 35430 30984 35436
rect 30288 35080 30340 35086
rect 30288 35022 30340 35028
rect 30944 34678 30972 35430
rect 31024 35012 31076 35018
rect 31024 34954 31076 34960
rect 30932 34672 30984 34678
rect 30932 34614 30984 34620
rect 30288 34536 30340 34542
rect 30288 34478 30340 34484
rect 30300 34202 30328 34478
rect 31036 34202 31064 34954
rect 30288 34196 30340 34202
rect 30288 34138 30340 34144
rect 31024 34196 31076 34202
rect 31024 34138 31076 34144
rect 30840 33856 30892 33862
rect 30840 33798 30892 33804
rect 30852 33522 30880 33798
rect 30656 33516 30708 33522
rect 30656 33458 30708 33464
rect 30840 33516 30892 33522
rect 30840 33458 30892 33464
rect 30668 32570 30696 33458
rect 30656 32564 30708 32570
rect 30656 32506 30708 32512
rect 30472 32360 30524 32366
rect 30472 32302 30524 32308
rect 30484 32026 30512 32302
rect 30472 32020 30524 32026
rect 30472 31962 30524 31968
rect 31128 31822 31156 46990
rect 31668 46368 31720 46374
rect 31668 46310 31720 46316
rect 31680 46034 31708 46310
rect 32232 46034 32260 49200
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 31668 46028 31720 46034
rect 31668 45970 31720 45976
rect 32220 46028 32272 46034
rect 32220 45970 32272 45976
rect 32220 45892 32272 45898
rect 32220 45834 32272 45840
rect 32232 45626 32260 45834
rect 32220 45620 32272 45626
rect 32220 45562 32272 45568
rect 38028 45554 38056 49200
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 38120 46578 38148 46990
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 38292 46504 38344 46510
rect 38292 46446 38344 46452
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 38304 46170 38332 46446
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38200 45960 38252 45966
rect 38200 45902 38252 45908
rect 37292 45526 38056 45554
rect 31944 45484 31996 45490
rect 31944 45426 31996 45432
rect 31956 44198 31984 45426
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 31944 44192 31996 44198
rect 31944 44134 31996 44140
rect 31852 35692 31904 35698
rect 31852 35634 31904 35640
rect 31760 35624 31812 35630
rect 31760 35566 31812 35572
rect 31300 35556 31352 35562
rect 31300 35498 31352 35504
rect 31208 34400 31260 34406
rect 31208 34342 31260 34348
rect 31220 33998 31248 34342
rect 31312 34202 31340 35498
rect 31772 34746 31800 35566
rect 31760 34740 31812 34746
rect 31760 34682 31812 34688
rect 31300 34196 31352 34202
rect 31300 34138 31352 34144
rect 31208 33992 31260 33998
rect 31208 33934 31260 33940
rect 31864 33522 31892 35634
rect 31208 33516 31260 33522
rect 31208 33458 31260 33464
rect 31852 33516 31904 33522
rect 31852 33458 31904 33464
rect 30656 31816 30708 31822
rect 30656 31758 30708 31764
rect 31116 31816 31168 31822
rect 31116 31758 31168 31764
rect 30564 31748 30616 31754
rect 30564 31690 30616 31696
rect 30576 31346 30604 31690
rect 30564 31340 30616 31346
rect 30564 31282 30616 31288
rect 30288 30728 30340 30734
rect 30288 30670 30340 30676
rect 30300 30258 30328 30670
rect 30472 30660 30524 30666
rect 30472 30602 30524 30608
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30380 30048 30432 30054
rect 30380 29990 30432 29996
rect 30392 29578 30420 29990
rect 30484 29714 30512 30602
rect 30576 30394 30604 31282
rect 30668 30734 30696 31758
rect 31220 31754 31248 33458
rect 31300 33312 31352 33318
rect 31300 33254 31352 33260
rect 31312 32978 31340 33254
rect 31864 33114 31892 33458
rect 31852 33108 31904 33114
rect 31852 33050 31904 33056
rect 31300 32972 31352 32978
rect 31300 32914 31352 32920
rect 31576 32428 31628 32434
rect 31576 32370 31628 32376
rect 31208 31748 31260 31754
rect 31208 31690 31260 31696
rect 30656 30728 30708 30734
rect 30656 30670 30708 30676
rect 30932 30728 30984 30734
rect 30932 30670 30984 30676
rect 30564 30388 30616 30394
rect 30564 30330 30616 30336
rect 30564 30252 30616 30258
rect 30564 30194 30616 30200
rect 30576 29850 30604 30194
rect 30668 30122 30696 30670
rect 30944 30598 30972 30670
rect 30748 30592 30800 30598
rect 30748 30534 30800 30540
rect 30932 30592 30984 30598
rect 30932 30534 30984 30540
rect 30656 30116 30708 30122
rect 30656 30058 30708 30064
rect 30564 29844 30616 29850
rect 30564 29786 30616 29792
rect 30760 29714 30788 30534
rect 30472 29708 30524 29714
rect 30472 29650 30524 29656
rect 30748 29708 30800 29714
rect 30748 29650 30800 29656
rect 30380 29572 30432 29578
rect 30380 29514 30432 29520
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30392 28762 30420 29106
rect 30380 28756 30432 28762
rect 30380 28698 30432 28704
rect 30484 28490 30512 29650
rect 30840 29028 30892 29034
rect 30840 28970 30892 28976
rect 30852 28626 30880 28970
rect 30840 28620 30892 28626
rect 30840 28562 30892 28568
rect 30472 28484 30524 28490
rect 30472 28426 30524 28432
rect 30840 28144 30892 28150
rect 30840 28086 30892 28092
rect 30656 28076 30708 28082
rect 30656 28018 30708 28024
rect 30668 27606 30696 28018
rect 30852 27606 30880 28086
rect 30656 27600 30708 27606
rect 30656 27542 30708 27548
rect 30840 27600 30892 27606
rect 30840 27542 30892 27548
rect 31300 25832 31352 25838
rect 31300 25774 31352 25780
rect 31312 25702 31340 25774
rect 31300 25696 31352 25702
rect 31300 25638 31352 25644
rect 31208 25220 31260 25226
rect 31208 25162 31260 25168
rect 30196 24200 30248 24206
rect 30196 24142 30248 24148
rect 29828 23860 29880 23866
rect 29828 23802 29880 23808
rect 31116 23656 31168 23662
rect 31116 23598 31168 23604
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 29828 23044 29880 23050
rect 29828 22986 29880 22992
rect 29840 22574 29868 22986
rect 30300 22642 30328 23122
rect 31128 22778 31156 23598
rect 30748 22772 30800 22778
rect 30748 22714 30800 22720
rect 31116 22772 31168 22778
rect 31116 22714 31168 22720
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 30564 22636 30616 22642
rect 30564 22578 30616 22584
rect 29828 22568 29880 22574
rect 29828 22510 29880 22516
rect 30288 22500 30340 22506
rect 30288 22442 30340 22448
rect 30300 22234 30328 22442
rect 30288 22228 30340 22234
rect 30288 22170 30340 22176
rect 29920 21888 29972 21894
rect 29920 21830 29972 21836
rect 29932 21622 29960 21830
rect 29920 21616 29972 21622
rect 29920 21558 29972 21564
rect 30300 21554 30328 22170
rect 30576 21962 30604 22578
rect 30760 22030 30788 22714
rect 31116 22568 31168 22574
rect 31116 22510 31168 22516
rect 31128 22166 31156 22510
rect 31220 22438 31248 25162
rect 31208 22432 31260 22438
rect 31208 22374 31260 22380
rect 31116 22160 31168 22166
rect 31116 22102 31168 22108
rect 30748 22024 30800 22030
rect 30748 21966 30800 21972
rect 30564 21956 30616 21962
rect 30564 21898 30616 21904
rect 31128 21894 31156 22102
rect 30380 21888 30432 21894
rect 30380 21830 30432 21836
rect 31116 21888 31168 21894
rect 31116 21830 31168 21836
rect 30392 21622 30420 21830
rect 30380 21616 30432 21622
rect 30380 21558 30432 21564
rect 30288 21548 30340 21554
rect 30288 21490 30340 21496
rect 30472 21344 30524 21350
rect 30472 21286 30524 21292
rect 31208 21344 31260 21350
rect 31208 21286 31260 21292
rect 30484 21010 30512 21286
rect 30472 21004 30524 21010
rect 30472 20946 30524 20952
rect 30196 20936 30248 20942
rect 30196 20878 30248 20884
rect 30208 20602 30236 20878
rect 31220 20874 31248 21286
rect 31208 20868 31260 20874
rect 31208 20810 31260 20816
rect 30196 20596 30248 20602
rect 30196 20538 30248 20544
rect 29368 19508 29420 19514
rect 29368 19450 29420 19456
rect 29366 19272 29422 19281
rect 29366 19207 29368 19216
rect 29420 19207 29422 19216
rect 30562 19272 30618 19281
rect 30562 19207 30564 19216
rect 29368 19178 29420 19184
rect 30616 19207 30618 19216
rect 30564 19178 30616 19184
rect 29552 18692 29604 18698
rect 29552 18634 29604 18640
rect 29460 4072 29512 4078
rect 29458 4040 29460 4049
rect 29512 4040 29514 4049
rect 29458 3975 29514 3984
rect 29564 3602 29592 18634
rect 30012 4072 30064 4078
rect 30012 4014 30064 4020
rect 29552 3596 29604 3602
rect 29552 3538 29604 3544
rect 29092 2916 29144 2922
rect 29092 2858 29144 2864
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 30024 2514 30052 4014
rect 31312 3398 31340 25638
rect 31484 23112 31536 23118
rect 31484 23054 31536 23060
rect 31496 22778 31524 23054
rect 31484 22772 31536 22778
rect 31484 22714 31536 22720
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31404 21554 31432 22578
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31390 19816 31446 19825
rect 31390 19751 31392 19760
rect 31444 19751 31446 19760
rect 31392 19722 31444 19728
rect 31300 3392 31352 3398
rect 31300 3334 31352 3340
rect 30932 2848 30984 2854
rect 30932 2790 30984 2796
rect 27160 2508 27212 2514
rect 27160 2450 27212 2456
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 28368 800 28396 2314
rect 29656 800 29684 2382
rect 30944 800 30972 2790
rect 31588 2310 31616 32370
rect 31956 26234 31984 44134
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 32128 35488 32180 35494
rect 32128 35430 32180 35436
rect 32140 35018 32168 35430
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 32128 35012 32180 35018
rect 32128 34954 32180 34960
rect 32864 34944 32916 34950
rect 32864 34886 32916 34892
rect 32128 34740 32180 34746
rect 32128 34682 32180 34688
rect 32140 33998 32168 34682
rect 32876 34678 32904 34886
rect 32864 34672 32916 34678
rect 32864 34614 32916 34620
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 32128 33992 32180 33998
rect 32128 33934 32180 33940
rect 32128 33652 32180 33658
rect 32128 33594 32180 33600
rect 32140 31414 32168 33594
rect 32772 33584 32824 33590
rect 32772 33526 32824 33532
rect 32312 33312 32364 33318
rect 32312 33254 32364 33260
rect 32324 32842 32352 33254
rect 32784 33114 32812 33526
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 32772 33108 32824 33114
rect 32772 33050 32824 33056
rect 32312 32836 32364 32842
rect 32312 32778 32364 32784
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 32312 31952 32364 31958
rect 32312 31894 32364 31900
rect 32128 31408 32180 31414
rect 32128 31350 32180 31356
rect 32036 31136 32088 31142
rect 32036 31078 32088 31084
rect 32048 30802 32076 31078
rect 32036 30796 32088 30802
rect 32036 30738 32088 30744
rect 32140 30326 32168 31350
rect 32324 31346 32352 31894
rect 32312 31340 32364 31346
rect 32312 31282 32364 31288
rect 32588 31340 32640 31346
rect 32588 31282 32640 31288
rect 32600 30938 32628 31282
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 32588 30932 32640 30938
rect 32588 30874 32640 30880
rect 32496 30660 32548 30666
rect 32496 30602 32548 30608
rect 32508 30326 32536 30602
rect 32128 30320 32180 30326
rect 32128 30262 32180 30268
rect 32496 30320 32548 30326
rect 32496 30262 32548 30268
rect 32220 30252 32272 30258
rect 32220 30194 32272 30200
rect 32128 29572 32180 29578
rect 32128 29514 32180 29520
rect 32140 29306 32168 29514
rect 32128 29300 32180 29306
rect 32128 29242 32180 29248
rect 32232 29186 32260 30194
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 32140 29170 32260 29186
rect 32128 29164 32260 29170
rect 32180 29158 32260 29164
rect 32128 29106 32180 29112
rect 32140 28082 32168 29106
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 32220 28484 32272 28490
rect 32220 28426 32272 28432
rect 32232 28218 32260 28426
rect 32220 28212 32272 28218
rect 32220 28154 32272 28160
rect 32128 28076 32180 28082
rect 32128 28018 32180 28024
rect 32140 26994 32168 28018
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 32128 26988 32180 26994
rect 32128 26930 32180 26936
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 32128 26376 32180 26382
rect 32128 26318 32180 26324
rect 32036 26240 32088 26246
rect 31956 26206 32036 26234
rect 32036 26182 32088 26188
rect 32048 24750 32076 26182
rect 32140 25974 32168 26318
rect 32312 26308 32364 26314
rect 32312 26250 32364 26256
rect 32324 25974 32352 26250
rect 32128 25968 32180 25974
rect 32128 25910 32180 25916
rect 32312 25968 32364 25974
rect 32312 25910 32364 25916
rect 32140 25294 32168 25910
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 32128 25288 32180 25294
rect 32128 25230 32180 25236
rect 32140 24818 32168 25230
rect 32772 25220 32824 25226
rect 32772 25162 32824 25168
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 32036 24744 32088 24750
rect 32036 24686 32088 24692
rect 31760 23588 31812 23594
rect 31760 23530 31812 23536
rect 32496 23588 32548 23594
rect 32496 23530 32548 23536
rect 31772 23186 31800 23530
rect 32036 23520 32088 23526
rect 32036 23462 32088 23468
rect 32048 23186 32076 23462
rect 32508 23186 32536 23530
rect 31760 23180 31812 23186
rect 31760 23122 31812 23128
rect 32036 23180 32088 23186
rect 32036 23122 32088 23128
rect 32496 23180 32548 23186
rect 32496 23122 32548 23128
rect 32496 23044 32548 23050
rect 32496 22986 32548 22992
rect 32508 22778 32536 22986
rect 32496 22772 32548 22778
rect 32496 22714 32548 22720
rect 31944 21956 31996 21962
rect 31944 21898 31996 21904
rect 31956 20806 31984 21898
rect 31944 20800 31996 20806
rect 31944 20742 31996 20748
rect 31956 20466 31984 20742
rect 31944 20460 31996 20466
rect 31944 20402 31996 20408
rect 32784 18290 32812 25162
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 33140 24336 33192 24342
rect 33140 24278 33192 24284
rect 33152 23662 33180 24278
rect 37292 23798 37320 45526
rect 38212 40118 38240 45902
rect 39960 45554 39988 49200
rect 40408 46980 40460 46986
rect 40408 46922 40460 46928
rect 39960 45526 40080 45554
rect 40052 44334 40080 45526
rect 38660 44328 38712 44334
rect 38660 44270 38712 44276
rect 38844 44328 38896 44334
rect 38844 44270 38896 44276
rect 40040 44328 40092 44334
rect 40040 44270 40092 44276
rect 38672 43110 38700 44270
rect 38856 43994 38884 44270
rect 38844 43988 38896 43994
rect 38844 43930 38896 43936
rect 38752 43784 38804 43790
rect 38752 43726 38804 43732
rect 38660 43104 38712 43110
rect 38660 43046 38712 43052
rect 38200 40112 38252 40118
rect 38200 40054 38252 40060
rect 38764 39438 38792 43726
rect 38752 39432 38804 39438
rect 38752 39374 38804 39380
rect 39948 39432 40000 39438
rect 39948 39374 40000 39380
rect 39960 37942 39988 39374
rect 39948 37936 40000 37942
rect 39948 37878 40000 37884
rect 38292 29232 38344 29238
rect 38292 29174 38344 29180
rect 37280 23792 37332 23798
rect 37280 23734 37332 23740
rect 33048 23656 33100 23662
rect 33048 23598 33100 23604
rect 33140 23656 33192 23662
rect 33140 23598 33192 23604
rect 33060 22778 33088 23598
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 33416 23112 33468 23118
rect 33416 23054 33468 23060
rect 33048 22772 33100 22778
rect 33048 22714 33100 22720
rect 33428 22642 33456 23054
rect 33876 22976 33928 22982
rect 33876 22918 33928 22924
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33428 20942 33456 22578
rect 33888 22574 33916 22918
rect 33876 22568 33928 22574
rect 33876 22510 33928 22516
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 33416 20936 33468 20942
rect 33416 20878 33468 20884
rect 33324 20800 33376 20806
rect 33324 20742 33376 20748
rect 33336 20534 33364 20742
rect 33324 20528 33376 20534
rect 33324 20470 33376 20476
rect 35440 20392 35492 20398
rect 35440 20334 35492 20340
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 33968 4004 34020 4010
rect 33968 3946 34020 3952
rect 33980 3738 34008 3946
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 33968 3732 34020 3738
rect 33968 3674 34020 3680
rect 35452 3670 35480 20334
rect 33048 3664 33100 3670
rect 33048 3606 33100 3612
rect 35440 3664 35492 3670
rect 35440 3606 35492 3612
rect 33060 3534 33088 3606
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 32956 3460 33008 3466
rect 32956 3402 33008 3408
rect 32864 3392 32916 3398
rect 32864 3334 32916 3340
rect 32220 3052 32272 3058
rect 32220 2994 32272 3000
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 32232 800 32260 2994
rect 32876 2854 32904 3334
rect 32968 3058 32996 3402
rect 33140 3392 33192 3398
rect 33140 3334 33192 3340
rect 33152 3126 33180 3334
rect 33140 3120 33192 3126
rect 33140 3062 33192 3068
rect 32956 3052 33008 3058
rect 32956 2994 33008 3000
rect 35912 2990 35940 3470
rect 36176 3460 36228 3466
rect 36176 3402 36228 3408
rect 36188 3194 36216 3402
rect 37924 3392 37976 3398
rect 37924 3334 37976 3340
rect 36176 3188 36228 3194
rect 36176 3130 36228 3136
rect 37936 3058 37964 3334
rect 36084 3052 36136 3058
rect 36084 2994 36136 3000
rect 37924 3052 37976 3058
rect 37924 2994 37976 3000
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 35900 2984 35952 2990
rect 35900 2926 35952 2932
rect 32864 2848 32916 2854
rect 32864 2790 32916 2796
rect 33520 800 33548 2926
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35452 800 35480 2382
rect 36096 800 36124 2994
rect 38304 2650 38332 29174
rect 40420 27402 40448 46922
rect 41248 46918 41276 49200
rect 41236 46912 41288 46918
rect 41236 46854 41288 46860
rect 41788 46912 41840 46918
rect 41788 46854 41840 46860
rect 41236 46368 41288 46374
rect 41236 46310 41288 46316
rect 41248 46034 41276 46310
rect 41236 46028 41288 46034
rect 41236 45970 41288 45976
rect 41420 45892 41472 45898
rect 41420 45834 41472 45840
rect 41432 45626 41460 45834
rect 41420 45620 41472 45626
rect 41420 45562 41472 45568
rect 41328 45484 41380 45490
rect 41328 45426 41380 45432
rect 41340 44470 41368 45426
rect 41328 44464 41380 44470
rect 41328 44406 41380 44412
rect 40408 27396 40460 27402
rect 40408 27338 40460 27344
rect 41236 25152 41288 25158
rect 41236 25094 41288 25100
rect 39764 23112 39816 23118
rect 39764 23054 39816 23060
rect 39948 23112 40000 23118
rect 39948 23054 40000 23060
rect 39776 22642 39804 23054
rect 39960 22710 39988 23054
rect 40132 23044 40184 23050
rect 40132 22986 40184 22992
rect 40144 22778 40172 22986
rect 40132 22772 40184 22778
rect 40132 22714 40184 22720
rect 39948 22704 40000 22710
rect 39948 22646 40000 22652
rect 39764 22636 39816 22642
rect 39764 22578 39816 22584
rect 41248 22030 41276 25094
rect 41236 22024 41288 22030
rect 41236 21966 41288 21972
rect 41340 20058 41368 44406
rect 41800 23186 41828 46854
rect 41892 46034 41920 49200
rect 42536 47138 42564 49200
rect 42536 47110 42748 47138
rect 42524 47048 42576 47054
rect 42524 46990 42576 46996
rect 41880 46028 41932 46034
rect 41880 45970 41932 45976
rect 42064 44872 42116 44878
rect 42064 44814 42116 44820
rect 42076 39370 42104 44814
rect 42536 44334 42564 46990
rect 42720 46510 42748 47110
rect 42800 46980 42852 46986
rect 42800 46922 42852 46928
rect 42616 46504 42668 46510
rect 42616 46446 42668 46452
rect 42708 46504 42760 46510
rect 42708 46446 42760 46452
rect 42628 45082 42656 46446
rect 42708 45416 42760 45422
rect 42708 45358 42760 45364
rect 42616 45076 42668 45082
rect 42616 45018 42668 45024
rect 42720 44402 42748 45358
rect 42812 45082 42840 46922
rect 43640 45778 43668 49286
rect 43782 49200 43894 50000
rect 44426 49314 44538 50000
rect 44426 49286 44864 49314
rect 44426 49200 44538 49286
rect 43824 45966 43852 49200
rect 44272 46436 44324 46442
rect 44272 46378 44324 46384
rect 43812 45960 43864 45966
rect 43812 45902 43864 45908
rect 43916 45886 44128 45914
rect 43916 45778 43944 45886
rect 43640 45750 43944 45778
rect 43996 45824 44048 45830
rect 43996 45766 44048 45772
rect 43812 45416 43864 45422
rect 43812 45358 43864 45364
rect 43824 45082 43852 45358
rect 42800 45076 42852 45082
rect 42800 45018 42852 45024
rect 43812 45076 43864 45082
rect 43812 45018 43864 45024
rect 43076 44872 43128 44878
rect 43076 44814 43128 44820
rect 42708 44396 42760 44402
rect 42708 44338 42760 44344
rect 42524 44328 42576 44334
rect 42524 44270 42576 44276
rect 42064 39364 42116 39370
rect 42064 39306 42116 39312
rect 41512 23180 41564 23186
rect 41512 23122 41564 23128
rect 41788 23180 41840 23186
rect 41788 23122 41840 23128
rect 41524 22710 41552 23122
rect 41512 22704 41564 22710
rect 41512 22646 41564 22652
rect 41524 22234 41552 22646
rect 41604 22568 41656 22574
rect 41604 22510 41656 22516
rect 41616 22438 41644 22510
rect 41604 22432 41656 22438
rect 41604 22374 41656 22380
rect 41512 22228 41564 22234
rect 41512 22170 41564 22176
rect 41328 20052 41380 20058
rect 41328 19994 41380 20000
rect 39304 19440 39356 19446
rect 39304 19382 39356 19388
rect 39212 4140 39264 4146
rect 39212 4082 39264 4088
rect 39120 3528 39172 3534
rect 39120 3470 39172 3476
rect 38568 3188 38620 3194
rect 38568 3130 38620 3136
rect 38580 2990 38608 3130
rect 38568 2984 38620 2990
rect 38568 2926 38620 2932
rect 39026 2952 39082 2961
rect 39026 2887 39028 2896
rect 39080 2887 39082 2896
rect 39028 2858 39080 2864
rect 39132 2650 39160 3470
rect 39224 2922 39252 4082
rect 39212 2916 39264 2922
rect 39212 2858 39264 2864
rect 39316 2650 39344 19382
rect 41616 12238 41644 22374
rect 42076 21690 42104 39306
rect 43088 25226 43116 44814
rect 43812 41064 43864 41070
rect 43812 41006 43864 41012
rect 43824 40118 43852 41006
rect 43812 40112 43864 40118
rect 43812 40054 43864 40060
rect 43720 39976 43772 39982
rect 43720 39918 43772 39924
rect 43536 27668 43588 27674
rect 43536 27610 43588 27616
rect 43444 26308 43496 26314
rect 43444 26250 43496 26256
rect 43456 25974 43484 26250
rect 43444 25968 43496 25974
rect 43444 25910 43496 25916
rect 43076 25220 43128 25226
rect 43076 25162 43128 25168
rect 42800 22976 42852 22982
rect 42800 22918 42852 22924
rect 42064 21684 42116 21690
rect 42064 21626 42116 21632
rect 42812 19378 42840 22918
rect 43548 22506 43576 27610
rect 43536 22500 43588 22506
rect 43536 22442 43588 22448
rect 42800 19372 42852 19378
rect 42800 19314 42852 19320
rect 43732 12434 43760 39918
rect 44008 35834 44036 45766
rect 44100 45422 44128 45886
rect 44088 45416 44140 45422
rect 44088 45358 44140 45364
rect 43996 35828 44048 35834
rect 43996 35770 44048 35776
rect 43996 21888 44048 21894
rect 43996 21830 44048 21836
rect 44008 21622 44036 21830
rect 43996 21616 44048 21622
rect 43996 21558 44048 21564
rect 43812 20800 43864 20806
rect 43812 20742 43864 20748
rect 43824 20534 43852 20742
rect 43812 20528 43864 20534
rect 43812 20470 43864 20476
rect 44284 19854 44312 46378
rect 44836 45554 44864 49286
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49314 46470 50000
rect 46216 49286 46470 49314
rect 45112 47122 45140 49200
rect 45100 47116 45152 47122
rect 45100 47058 45152 47064
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45100 45554 45152 45558
rect 44836 45552 45152 45554
rect 44836 45526 45100 45552
rect 45100 45494 45152 45500
rect 45100 45280 45152 45286
rect 45100 45222 45152 45228
rect 45112 31482 45140 45222
rect 45204 43314 45232 46990
rect 45376 46980 45428 46986
rect 45376 46922 45428 46928
rect 45388 45558 45416 46922
rect 45756 45966 45784 49200
rect 46020 46504 46072 46510
rect 46020 46446 46072 46452
rect 45928 46096 45980 46102
rect 45928 46038 45980 46044
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 45376 45552 45428 45558
rect 45376 45494 45428 45500
rect 45836 45416 45888 45422
rect 45836 45358 45888 45364
rect 45652 45348 45704 45354
rect 45652 45290 45704 45296
rect 45664 44878 45692 45290
rect 45652 44872 45704 44878
rect 45652 44814 45704 44820
rect 45744 44872 45796 44878
rect 45744 44814 45796 44820
rect 45192 43308 45244 43314
rect 45192 43250 45244 43256
rect 45664 42226 45692 44814
rect 45756 44402 45784 44814
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 45652 42220 45704 42226
rect 45652 42162 45704 42168
rect 45560 40452 45612 40458
rect 45560 40394 45612 40400
rect 45572 38758 45600 40394
rect 45848 38962 45876 45358
rect 45940 44402 45968 46038
rect 46032 44538 46060 46446
rect 46216 45490 46244 49286
rect 46358 49200 46470 49286
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 46846 47696 46902 47705
rect 46846 47631 46902 47640
rect 46860 46510 46888 47631
rect 46848 46504 46900 46510
rect 46848 46446 46900 46452
rect 46940 46436 46992 46442
rect 46940 46378 46992 46384
rect 46296 45960 46348 45966
rect 46296 45902 46348 45908
rect 46204 45484 46256 45490
rect 46204 45426 46256 45432
rect 46308 45014 46336 45902
rect 46480 45892 46532 45898
rect 46480 45834 46532 45840
rect 46492 45082 46520 45834
rect 46572 45824 46624 45830
rect 46572 45766 46624 45772
rect 46480 45076 46532 45082
rect 46480 45018 46532 45024
rect 46296 45008 46348 45014
rect 46296 44950 46348 44956
rect 46020 44532 46072 44538
rect 46020 44474 46072 44480
rect 45928 44396 45980 44402
rect 45928 44338 45980 44344
rect 46480 42016 46532 42022
rect 46480 41958 46532 41964
rect 46492 41682 46520 41958
rect 46480 41676 46532 41682
rect 46480 41618 46532 41624
rect 46202 41168 46258 41177
rect 46202 41103 46204 41112
rect 46256 41103 46258 41112
rect 46204 41074 46256 41080
rect 46020 40112 46072 40118
rect 46020 40054 46072 40060
rect 45652 38956 45704 38962
rect 45652 38898 45704 38904
rect 45836 38956 45888 38962
rect 45836 38898 45888 38904
rect 45560 38752 45612 38758
rect 45560 38694 45612 38700
rect 45664 38350 45692 38898
rect 45848 38486 45876 38898
rect 45836 38480 45888 38486
rect 45836 38422 45888 38428
rect 45652 38344 45704 38350
rect 45652 38286 45704 38292
rect 45560 37936 45612 37942
rect 45560 37878 45612 37884
rect 45572 37330 45600 37878
rect 45560 37324 45612 37330
rect 45560 37266 45612 37272
rect 45664 37262 45692 38286
rect 45744 37868 45796 37874
rect 45744 37810 45796 37816
rect 45756 37466 45784 37810
rect 45744 37460 45796 37466
rect 45744 37402 45796 37408
rect 45744 37324 45796 37330
rect 45744 37266 45796 37272
rect 45652 37256 45704 37262
rect 45652 37198 45704 37204
rect 45100 31476 45152 31482
rect 45100 31418 45152 31424
rect 45560 31204 45612 31210
rect 45560 31146 45612 31152
rect 45572 26466 45600 31146
rect 45664 31090 45692 37198
rect 45756 35894 45784 37266
rect 45848 37262 45876 38422
rect 45928 38344 45980 38350
rect 45928 38286 45980 38292
rect 45940 37806 45968 38286
rect 46032 38010 46060 40054
rect 46386 38992 46442 39001
rect 46386 38927 46388 38936
rect 46440 38927 46442 38936
rect 46388 38898 46440 38904
rect 46112 38752 46164 38758
rect 46112 38694 46164 38700
rect 46124 38214 46152 38694
rect 46584 38554 46612 45766
rect 46664 44804 46716 44810
rect 46664 44746 46716 44752
rect 46676 44538 46704 44746
rect 46664 44532 46716 44538
rect 46664 44474 46716 44480
rect 46952 43314 46980 46378
rect 47044 46034 47072 49200
rect 47688 47054 47716 49200
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47860 46572 47912 46578
rect 47860 46514 47912 46520
rect 47872 46345 47900 46514
rect 48044 46368 48096 46374
rect 47858 46336 47914 46345
rect 48044 46310 48096 46316
rect 47858 46271 47914 46280
rect 47032 46028 47084 46034
rect 47032 45970 47084 45976
rect 47492 45484 47544 45490
rect 47492 45426 47544 45432
rect 47504 44402 47532 45426
rect 47584 44736 47636 44742
rect 47584 44678 47636 44684
rect 47492 44396 47544 44402
rect 47492 44338 47544 44344
rect 46940 43308 46992 43314
rect 46940 43250 46992 43256
rect 47308 42220 47360 42226
rect 47308 42162 47360 42168
rect 46848 38888 46900 38894
rect 46848 38830 46900 38836
rect 46572 38548 46624 38554
rect 46572 38490 46624 38496
rect 46112 38208 46164 38214
rect 46112 38150 46164 38156
rect 46020 38004 46072 38010
rect 46020 37946 46072 37952
rect 46124 37874 46152 38150
rect 46112 37868 46164 37874
rect 46112 37810 46164 37816
rect 45928 37800 45980 37806
rect 45928 37742 45980 37748
rect 45836 37256 45888 37262
rect 45836 37198 45888 37204
rect 45756 35866 45876 35894
rect 45664 31062 45784 31090
rect 45480 26438 45600 26466
rect 45480 26194 45508 26438
rect 45652 26240 45704 26246
rect 45480 26166 45600 26194
rect 45652 26182 45704 26188
rect 45572 25158 45600 26166
rect 45664 25906 45692 26182
rect 45652 25900 45704 25906
rect 45652 25842 45704 25848
rect 45664 25294 45692 25842
rect 45652 25288 45704 25294
rect 45652 25230 45704 25236
rect 45560 25152 45612 25158
rect 45560 25094 45612 25100
rect 45376 24744 45428 24750
rect 45376 24686 45428 24692
rect 45008 24676 45060 24682
rect 45284 24676 45336 24682
rect 45060 24636 45284 24664
rect 45008 24618 45060 24624
rect 45284 24618 45336 24624
rect 45388 23866 45416 24686
rect 45560 24064 45612 24070
rect 45560 24006 45612 24012
rect 45376 23860 45428 23866
rect 45376 23802 45428 23808
rect 44732 23656 44784 23662
rect 44732 23598 44784 23604
rect 44744 22098 44772 23598
rect 44732 22092 44784 22098
rect 44732 22034 44784 22040
rect 45572 22030 45600 24006
rect 45560 22024 45612 22030
rect 45560 21966 45612 21972
rect 45376 21480 45428 21486
rect 45376 21422 45428 21428
rect 44272 19848 44324 19854
rect 44272 19790 44324 19796
rect 44284 19718 44312 19790
rect 44272 19712 44324 19718
rect 44272 19654 44324 19660
rect 43732 12406 43852 12434
rect 41604 12232 41656 12238
rect 41604 12174 41656 12180
rect 43536 4684 43588 4690
rect 43536 4626 43588 4632
rect 42892 4616 42944 4622
rect 42892 4558 42944 4564
rect 41328 4072 41380 4078
rect 41328 4014 41380 4020
rect 40040 3936 40092 3942
rect 40040 3878 40092 3884
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 39856 3460 39908 3466
rect 39856 3402 39908 3408
rect 39868 2990 39896 3402
rect 39856 2984 39908 2990
rect 39856 2926 39908 2932
rect 38292 2644 38344 2650
rect 38292 2586 38344 2592
rect 39120 2644 39172 2650
rect 39120 2586 39172 2592
rect 39304 2644 39356 2650
rect 39304 2586 39356 2592
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 38028 800 38056 2382
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 39316 800 39344 2314
rect 39960 800 39988 3470
rect 40052 2446 40080 3878
rect 41340 3534 41368 4014
rect 42800 3936 42852 3942
rect 42800 3878 42852 3884
rect 42524 3664 42576 3670
rect 42524 3606 42576 3612
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41512 3528 41564 3534
rect 41512 3470 41564 3476
rect 40132 3392 40184 3398
rect 40132 3334 40184 3340
rect 40144 2854 40172 3334
rect 41236 3188 41288 3194
rect 41340 3176 41368 3470
rect 41288 3148 41368 3176
rect 41236 3130 41288 3136
rect 41524 3126 41552 3470
rect 42432 3392 42484 3398
rect 42432 3334 42484 3340
rect 41512 3120 41564 3126
rect 41512 3062 41564 3068
rect 40132 2848 40184 2854
rect 40132 2790 40184 2796
rect 41524 2514 41552 3062
rect 42444 3058 42472 3334
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 41512 2508 41564 2514
rect 41512 2450 41564 2456
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40604 800 40632 2314
rect 41248 800 41276 2382
rect 42536 800 42564 3606
rect 42812 3602 42840 3878
rect 42904 3670 42932 4558
rect 43444 4140 43496 4146
rect 43444 4082 43496 4088
rect 43456 3738 43484 4082
rect 43548 4078 43576 4626
rect 43824 4078 43852 12406
rect 43536 4072 43588 4078
rect 43536 4014 43588 4020
rect 43720 4072 43772 4078
rect 43720 4014 43772 4020
rect 43812 4072 43864 4078
rect 43812 4014 43864 4020
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 42892 3664 42944 3670
rect 42892 3606 42944 3612
rect 42800 3596 42852 3602
rect 42800 3538 42852 3544
rect 43168 3596 43220 3602
rect 43168 3538 43220 3544
rect 43180 800 43208 3538
rect 43732 2650 43760 4014
rect 43824 3505 43852 4014
rect 43810 3496 43866 3505
rect 44284 3466 44312 19654
rect 45388 12434 45416 21422
rect 45572 20942 45600 21966
rect 45560 20936 45612 20942
rect 45560 20878 45612 20884
rect 45468 20392 45520 20398
rect 45468 20334 45520 20340
rect 45560 20392 45612 20398
rect 45560 20334 45612 20340
rect 45296 12406 45416 12434
rect 44364 5772 44416 5778
rect 44364 5714 44416 5720
rect 43810 3431 43866 3440
rect 44272 3460 44324 3466
rect 44272 3402 44324 3408
rect 44376 3126 44404 5714
rect 45296 3194 45324 12406
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45284 3188 45336 3194
rect 45284 3130 45336 3136
rect 45388 3126 45416 3334
rect 44364 3120 44416 3126
rect 44364 3062 44416 3068
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 44364 2848 44416 2854
rect 44364 2790 44416 2796
rect 44376 2650 44404 2790
rect 45480 2774 45508 20334
rect 45572 19922 45600 20334
rect 45560 19916 45612 19922
rect 45560 19858 45612 19864
rect 45560 16448 45612 16454
rect 45560 16390 45612 16396
rect 45572 15745 45600 16390
rect 45558 15736 45614 15745
rect 45558 15671 45614 15680
rect 45560 8288 45612 8294
rect 45558 8256 45560 8265
rect 45612 8256 45614 8265
rect 45558 8191 45614 8200
rect 45652 4616 45704 4622
rect 45652 4558 45704 4564
rect 45664 2990 45692 4558
rect 45756 4214 45784 31062
rect 45848 24070 45876 35866
rect 45836 24064 45888 24070
rect 45836 24006 45888 24012
rect 45836 23724 45888 23730
rect 45836 23666 45888 23672
rect 45848 22778 45876 23666
rect 45836 22772 45888 22778
rect 45836 22714 45888 22720
rect 45836 22636 45888 22642
rect 45836 22578 45888 22584
rect 45848 22234 45876 22578
rect 45940 22506 45968 37742
rect 46020 37732 46072 37738
rect 46020 37674 46072 37680
rect 46032 37398 46060 37674
rect 46480 37664 46532 37670
rect 46480 37606 46532 37612
rect 46020 37392 46072 37398
rect 46020 37334 46072 37340
rect 46032 31210 46060 37334
rect 46492 37330 46520 37606
rect 46860 37398 46888 38830
rect 46848 37392 46900 37398
rect 46848 37334 46900 37340
rect 46480 37324 46532 37330
rect 46480 37266 46532 37272
rect 47124 34944 47176 34950
rect 47124 34886 47176 34892
rect 46572 34536 46624 34542
rect 46572 34478 46624 34484
rect 46112 34128 46164 34134
rect 46112 34070 46164 34076
rect 46020 31204 46072 31210
rect 46020 31146 46072 31152
rect 46020 25152 46072 25158
rect 46020 25094 46072 25100
rect 46032 24274 46060 25094
rect 46020 24268 46072 24274
rect 46020 24210 46072 24216
rect 46020 23112 46072 23118
rect 46020 23054 46072 23060
rect 46032 22545 46060 23054
rect 46018 22536 46074 22545
rect 45928 22500 45980 22506
rect 46018 22471 46074 22480
rect 45928 22442 45980 22448
rect 45836 22228 45888 22234
rect 45836 22170 45888 22176
rect 46124 22114 46152 34070
rect 46296 32904 46348 32910
rect 46296 32846 46348 32852
rect 46308 32434 46336 32846
rect 46296 32428 46348 32434
rect 46296 32370 46348 32376
rect 46584 31822 46612 34478
rect 47136 34066 47164 34886
rect 47216 34400 47268 34406
rect 47216 34342 47268 34348
rect 47124 34060 47176 34066
rect 47124 34002 47176 34008
rect 47228 33930 47256 34342
rect 47216 33924 47268 33930
rect 47216 33866 47268 33872
rect 47320 32178 47348 42162
rect 47504 32434 47532 44338
rect 47596 42226 47624 44678
rect 47676 44192 47728 44198
rect 47676 44134 47728 44140
rect 47688 43858 47716 44134
rect 47676 43852 47728 43858
rect 47676 43794 47728 43800
rect 47768 43104 47820 43110
rect 47768 43046 47820 43052
rect 47780 42770 47808 43046
rect 47768 42764 47820 42770
rect 47768 42706 47820 42712
rect 47676 42628 47728 42634
rect 47676 42570 47728 42576
rect 47688 42362 47716 42570
rect 47676 42356 47728 42362
rect 47676 42298 47728 42304
rect 47584 42220 47636 42226
rect 47584 42162 47636 42168
rect 47768 41540 47820 41546
rect 47768 41482 47820 41488
rect 47780 41138 47808 41482
rect 47768 41132 47820 41138
rect 47768 41074 47820 41080
rect 47768 40588 47820 40594
rect 47768 40530 47820 40536
rect 47780 40050 47808 40530
rect 47768 40044 47820 40050
rect 47768 39986 47820 39992
rect 47860 39500 47912 39506
rect 47860 39442 47912 39448
rect 47676 39364 47728 39370
rect 47676 39306 47728 39312
rect 47688 39098 47716 39306
rect 47676 39092 47728 39098
rect 47676 39034 47728 39040
rect 47676 38956 47728 38962
rect 47676 38898 47728 38904
rect 47688 35894 47716 38898
rect 47872 38282 47900 39442
rect 47860 38276 47912 38282
rect 47860 38218 47912 38224
rect 47768 37664 47820 37670
rect 47768 37606 47820 37612
rect 47780 37194 47808 37606
rect 47768 37188 47820 37194
rect 47768 37130 47820 37136
rect 47596 35866 47716 35894
rect 47492 32428 47544 32434
rect 47492 32370 47544 32376
rect 47228 32150 47348 32178
rect 46572 31816 46624 31822
rect 46572 31758 46624 31764
rect 46386 31376 46442 31385
rect 46386 31311 46442 31320
rect 46294 30016 46350 30025
rect 46294 29951 46350 29960
rect 46202 28656 46258 28665
rect 46202 28591 46258 28600
rect 46216 27674 46244 28591
rect 46204 27668 46256 27674
rect 46204 27610 46256 27616
rect 46308 27554 46336 29951
rect 46216 27526 46336 27554
rect 46216 26042 46244 27526
rect 46294 26616 46350 26625
rect 46294 26551 46350 26560
rect 46308 26314 46336 26551
rect 46296 26308 46348 26314
rect 46296 26250 46348 26256
rect 46204 26036 46256 26042
rect 46204 25978 46256 25984
rect 46296 25764 46348 25770
rect 46296 25706 46348 25712
rect 46204 24676 46256 24682
rect 46204 24618 46256 24624
rect 46216 23905 46244 24618
rect 46202 23896 46258 23905
rect 46202 23831 46258 23840
rect 46308 23186 46336 25706
rect 46400 23746 46428 31311
rect 46572 28484 46624 28490
rect 46572 28426 46624 28432
rect 46480 25696 46532 25702
rect 46480 25638 46532 25644
rect 46492 25362 46520 25638
rect 46480 25356 46532 25362
rect 46480 25298 46532 25304
rect 46584 25226 46612 28426
rect 47124 28076 47176 28082
rect 47124 28018 47176 28024
rect 47032 27872 47084 27878
rect 47032 27814 47084 27820
rect 47044 27538 47072 27814
rect 47032 27532 47084 27538
rect 47032 27474 47084 27480
rect 47136 26518 47164 28018
rect 47124 26512 47176 26518
rect 47124 26454 47176 26460
rect 46940 26444 46992 26450
rect 46940 26386 46992 26392
rect 46754 25256 46810 25265
rect 46572 25220 46624 25226
rect 46754 25191 46810 25200
rect 46572 25162 46624 25168
rect 46400 23718 46520 23746
rect 46388 23656 46440 23662
rect 46388 23598 46440 23604
rect 46296 23180 46348 23186
rect 46296 23122 46348 23128
rect 46204 22568 46256 22574
rect 46204 22510 46256 22516
rect 45940 22086 46152 22114
rect 45836 22024 45888 22030
rect 45836 21966 45888 21972
rect 45848 21554 45876 21966
rect 45940 21894 45968 22086
rect 45928 21888 45980 21894
rect 45928 21830 45980 21836
rect 45940 21554 45968 21830
rect 46216 21690 46244 22510
rect 46400 22386 46428 23598
rect 46308 22358 46428 22386
rect 46308 22030 46336 22358
rect 46492 22094 46520 23718
rect 46400 22066 46520 22094
rect 46296 22024 46348 22030
rect 46296 21966 46348 21972
rect 46296 21888 46348 21894
rect 46296 21830 46348 21836
rect 46204 21684 46256 21690
rect 46204 21626 46256 21632
rect 46308 21554 46336 21830
rect 45836 21548 45888 21554
rect 45836 21490 45888 21496
rect 45928 21548 45980 21554
rect 45928 21490 45980 21496
rect 46296 21548 46348 21554
rect 46296 21490 46348 21496
rect 45940 10538 45968 21490
rect 46020 19848 46072 19854
rect 46020 19790 46072 19796
rect 46032 19310 46060 19790
rect 46020 19304 46072 19310
rect 46020 19246 46072 19252
rect 46308 18578 46336 21490
rect 46400 21078 46428 22066
rect 46480 21344 46532 21350
rect 46480 21286 46532 21292
rect 46388 21072 46440 21078
rect 46388 21014 46440 21020
rect 46492 21010 46520 21286
rect 46480 21004 46532 21010
rect 46480 20946 46532 20952
rect 46388 20460 46440 20466
rect 46388 20402 46440 20408
rect 46400 19854 46428 20402
rect 46584 19922 46612 25162
rect 46664 23724 46716 23730
rect 46664 23666 46716 23672
rect 46676 23066 46704 23666
rect 46768 23186 46796 25191
rect 46848 24744 46900 24750
rect 46848 24686 46900 24692
rect 46860 24585 46888 24686
rect 46846 24576 46902 24585
rect 46846 24511 46902 24520
rect 46952 24154 46980 26386
rect 46952 24138 47072 24154
rect 46952 24132 47084 24138
rect 46952 24126 47032 24132
rect 47032 24074 47084 24080
rect 46848 23588 46900 23594
rect 46848 23530 46900 23536
rect 46860 23225 46888 23530
rect 46846 23216 46902 23225
rect 46756 23180 46808 23186
rect 46846 23151 46902 23160
rect 46756 23122 46808 23128
rect 46676 23038 46796 23066
rect 46768 22574 46796 23038
rect 46756 22568 46808 22574
rect 46756 22510 46808 22516
rect 46664 21548 46716 21554
rect 46664 21490 46716 21496
rect 46572 19916 46624 19922
rect 46572 19858 46624 19864
rect 46388 19848 46440 19854
rect 46388 19790 46440 19796
rect 46572 19780 46624 19786
rect 46572 19722 46624 19728
rect 46308 18550 46428 18578
rect 46296 16992 46348 16998
rect 46296 16934 46348 16940
rect 46308 16658 46336 16934
rect 46296 16652 46348 16658
rect 46296 16594 46348 16600
rect 46296 15904 46348 15910
rect 46296 15846 46348 15852
rect 46308 15570 46336 15846
rect 46296 15564 46348 15570
rect 46296 15506 46348 15512
rect 46296 13320 46348 13326
rect 46296 13262 46348 13268
rect 46308 12850 46336 13262
rect 46296 12844 46348 12850
rect 46296 12786 46348 12792
rect 46296 11552 46348 11558
rect 46296 11494 46348 11500
rect 46308 11218 46336 11494
rect 46296 11212 46348 11218
rect 46296 11154 46348 11160
rect 46112 10736 46164 10742
rect 46112 10678 46164 10684
rect 46020 10600 46072 10606
rect 46020 10542 46072 10548
rect 45928 10532 45980 10538
rect 45928 10474 45980 10480
rect 46032 5302 46060 10542
rect 46124 9722 46152 10678
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46308 10130 46336 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 46112 9716 46164 9722
rect 46112 9658 46164 9664
rect 46204 6248 46256 6254
rect 46202 6216 46204 6225
rect 46256 6216 46258 6225
rect 46202 6151 46258 6160
rect 46400 6066 46428 18550
rect 46480 12096 46532 12102
rect 46480 12038 46532 12044
rect 46492 11218 46520 12038
rect 46480 11212 46532 11218
rect 46480 11154 46532 11160
rect 46584 6322 46612 19722
rect 46572 6316 46624 6322
rect 46572 6258 46624 6264
rect 46216 6038 46428 6066
rect 46020 5296 46072 5302
rect 46020 5238 46072 5244
rect 46032 4690 46060 5238
rect 46020 4684 46072 4690
rect 46020 4626 46072 4632
rect 45744 4208 45796 4214
rect 45744 4150 45796 4156
rect 45652 2984 45704 2990
rect 45652 2926 45704 2932
rect 45112 2746 45508 2774
rect 43720 2644 43772 2650
rect 43720 2586 43772 2592
rect 44364 2644 44416 2650
rect 44364 2586 44416 2592
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 44180 2440 44232 2446
rect 44180 2382 44232 2388
rect 43824 800 43852 2382
rect 2870 776 2926 785
rect 2870 711 2926 720
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44192 542 44220 2382
rect 45112 800 45140 2746
rect 46216 2530 46244 6038
rect 46480 5636 46532 5642
rect 46480 5578 46532 5584
rect 46296 4548 46348 4554
rect 46296 4490 46348 4496
rect 46124 2514 46244 2530
rect 46112 2508 46244 2514
rect 46164 2502 46244 2508
rect 46112 2450 46164 2456
rect 46308 2446 46336 4490
rect 46492 4146 46520 5578
rect 46572 4684 46624 4690
rect 46572 4626 46624 4632
rect 46584 4214 46612 4626
rect 46572 4208 46624 4214
rect 46572 4150 46624 4156
rect 46480 4140 46532 4146
rect 46480 4082 46532 4088
rect 46676 3738 46704 21490
rect 46768 20330 46796 22510
rect 46940 20460 46992 20466
rect 46940 20402 46992 20408
rect 46756 20324 46808 20330
rect 46756 20266 46808 20272
rect 46952 20058 46980 20402
rect 46940 20052 46992 20058
rect 46940 19994 46992 20000
rect 46848 19508 46900 19514
rect 46848 19450 46900 19456
rect 46860 18290 46888 19450
rect 46940 19372 46992 19378
rect 46940 19314 46992 19320
rect 46952 18426 46980 19314
rect 47044 19310 47072 24074
rect 47032 19304 47084 19310
rect 47032 19246 47084 19252
rect 47030 18456 47086 18465
rect 46940 18420 46992 18426
rect 47030 18391 47086 18400
rect 46940 18362 46992 18368
rect 46848 18284 46900 18290
rect 46848 18226 46900 18232
rect 47044 17678 47072 18391
rect 47032 17672 47084 17678
rect 47032 17614 47084 17620
rect 47136 16114 47164 26454
rect 47228 26234 47256 32150
rect 47306 32056 47362 32065
rect 47306 31991 47362 32000
rect 47320 31890 47348 31991
rect 47308 31884 47360 31890
rect 47308 31826 47360 31832
rect 47308 29640 47360 29646
rect 47308 29582 47360 29588
rect 47400 29640 47452 29646
rect 47400 29582 47452 29588
rect 47320 29345 47348 29582
rect 47306 29336 47362 29345
rect 47306 29271 47362 29280
rect 47412 28626 47440 29582
rect 47400 28620 47452 28626
rect 47400 28562 47452 28568
rect 47504 26234 47532 32370
rect 47596 28082 47624 35866
rect 47768 33516 47820 33522
rect 47768 33458 47820 33464
rect 47780 33425 47808 33458
rect 47766 33416 47822 33425
rect 47766 33351 47822 33360
rect 47676 32836 47728 32842
rect 47676 32778 47728 32784
rect 47688 32570 47716 32778
rect 47676 32564 47728 32570
rect 47676 32506 47728 32512
rect 47676 28620 47728 28626
rect 47676 28562 47728 28568
rect 47688 28218 47716 28562
rect 47676 28212 47728 28218
rect 47676 28154 47728 28160
rect 47584 28076 47636 28082
rect 47584 28018 47636 28024
rect 47688 27962 47716 28154
rect 47688 27934 47808 27962
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 47688 27402 47716 27814
rect 47676 27396 47728 27402
rect 47676 27338 47728 27344
rect 47780 26450 47808 27934
rect 47768 26444 47820 26450
rect 47768 26386 47820 26392
rect 47228 26206 47348 26234
rect 47320 24426 47348 26206
rect 47412 26206 47532 26234
rect 47412 25838 47440 26206
rect 47400 25832 47452 25838
rect 47400 25774 47452 25780
rect 47320 24398 47532 24426
rect 47308 24268 47360 24274
rect 47308 24210 47360 24216
rect 47216 19440 47268 19446
rect 47216 19382 47268 19388
rect 47228 18290 47256 19382
rect 47216 18284 47268 18290
rect 47216 18226 47268 18232
rect 47228 17882 47256 18226
rect 47216 17876 47268 17882
rect 47216 17818 47268 17824
rect 47124 16108 47176 16114
rect 47124 16050 47176 16056
rect 47136 13938 47164 16050
rect 47124 13932 47176 13938
rect 47124 13874 47176 13880
rect 47320 12434 47348 24210
rect 47504 23730 47532 24398
rect 47492 23724 47544 23730
rect 47492 23666 47544 23672
rect 47504 22438 47532 23666
rect 47584 23316 47636 23322
rect 47584 23258 47636 23264
rect 47596 22642 47624 23258
rect 47676 23044 47728 23050
rect 47676 22986 47728 22992
rect 47688 22778 47716 22986
rect 47676 22772 47728 22778
rect 47676 22714 47728 22720
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 47492 22432 47544 22438
rect 47492 22374 47544 22380
rect 47504 19378 47532 22374
rect 47492 19372 47544 19378
rect 47492 19314 47544 19320
rect 47492 18284 47544 18290
rect 47492 18226 47544 18232
rect 47504 17610 47532 18226
rect 47492 17604 47544 17610
rect 47492 17546 47544 17552
rect 47596 17202 47624 22578
rect 47780 22098 47808 26386
rect 47768 22092 47820 22098
rect 47768 22034 47820 22040
rect 47768 20868 47820 20874
rect 47768 20810 47820 20816
rect 47780 20466 47808 20810
rect 47768 20460 47820 20466
rect 47768 20402 47820 20408
rect 47768 19372 47820 19378
rect 47768 19314 47820 19320
rect 47676 19168 47728 19174
rect 47676 19110 47728 19116
rect 47688 18834 47716 19110
rect 47676 18828 47728 18834
rect 47676 18770 47728 18776
rect 47780 18714 47808 19314
rect 47688 18686 47808 18714
rect 47688 17490 47716 18686
rect 47768 18284 47820 18290
rect 47768 18226 47820 18232
rect 47780 17678 47808 18226
rect 47768 17672 47820 17678
rect 47768 17614 47820 17620
rect 47688 17462 47808 17490
rect 47584 17196 47636 17202
rect 47584 17138 47636 17144
rect 47596 12434 47624 17138
rect 47676 16992 47728 16998
rect 47676 16934 47728 16940
rect 47688 16522 47716 16934
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 47676 15904 47728 15910
rect 47676 15846 47728 15852
rect 47688 15570 47716 15846
rect 47676 15564 47728 15570
rect 47676 15506 47728 15512
rect 47676 13728 47728 13734
rect 47676 13670 47728 13676
rect 47688 13394 47716 13670
rect 47676 13388 47728 13394
rect 47676 13330 47728 13336
rect 47228 12406 47348 12434
rect 47504 12406 47624 12434
rect 46846 9616 46902 9625
rect 46846 9551 46848 9560
rect 46900 9551 46902 9560
rect 46848 9522 46900 9528
rect 47032 7200 47084 7206
rect 47032 7142 47084 7148
rect 47044 6866 47072 7142
rect 47032 6860 47084 6866
rect 47032 6802 47084 6808
rect 46664 3732 46716 3738
rect 46664 3674 46716 3680
rect 47228 3670 47256 12406
rect 47504 9586 47532 12406
rect 47676 9988 47728 9994
rect 47676 9930 47728 9936
rect 47688 9654 47716 9930
rect 47676 9648 47728 9654
rect 47676 9590 47728 9596
rect 47492 9580 47544 9586
rect 47492 9522 47544 9528
rect 47308 8968 47360 8974
rect 47308 8910 47360 8916
rect 47400 8968 47452 8974
rect 47400 8910 47452 8916
rect 47320 7585 47348 8910
rect 47412 7954 47440 8910
rect 47400 7948 47452 7954
rect 47400 7890 47452 7896
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47216 3664 47268 3670
rect 47216 3606 47268 3612
rect 47504 3466 47532 9522
rect 47674 8936 47730 8945
rect 47674 8871 47730 8880
rect 47688 8498 47716 8871
rect 47676 8492 47728 8498
rect 47676 8434 47728 8440
rect 47676 7948 47728 7954
rect 47676 7890 47728 7896
rect 47688 5778 47716 7890
rect 47676 5772 47728 5778
rect 47676 5714 47728 5720
rect 47780 5234 47808 17462
rect 47872 8022 47900 38218
rect 48056 26314 48084 46310
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48136 44940 48188 44946
rect 48136 44882 48188 44888
rect 48134 44568 48190 44577
rect 48134 44503 48190 44512
rect 48148 43858 48176 44503
rect 48136 43852 48188 43858
rect 48136 43794 48188 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 41857 48176 42570
rect 48134 41848 48190 41857
rect 48134 41783 48190 41792
rect 48136 41540 48188 41546
rect 48136 41482 48188 41488
rect 48148 41449 48176 41482
rect 48134 41440 48190 41449
rect 48134 41375 48190 41384
rect 48136 40452 48188 40458
rect 48136 40394 48188 40400
rect 48148 40089 48176 40394
rect 48134 40080 48190 40089
rect 48134 40015 48190 40024
rect 48136 39364 48188 39370
rect 48136 39306 48188 39312
rect 48148 39137 48176 39306
rect 48134 39128 48190 39137
rect 48134 39063 48190 39072
rect 48134 37768 48190 37777
rect 48134 37703 48190 37712
rect 48148 37330 48176 37703
rect 48136 37324 48188 37330
rect 48136 37266 48188 37272
rect 48136 35080 48188 35086
rect 48136 35022 48188 35028
rect 48148 34785 48176 35022
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48136 34604 48188 34610
rect 48136 34546 48188 34552
rect 48148 34105 48176 34546
rect 48134 34096 48190 34105
rect 48134 34031 48190 34040
rect 48136 32836 48188 32842
rect 48136 32778 48188 32784
rect 48148 32745 48176 32778
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48044 26308 48096 26314
rect 48044 26250 48096 26256
rect 48134 25936 48190 25945
rect 48134 25871 48190 25880
rect 48148 25362 48176 25871
rect 48136 25356 48188 25362
rect 48136 25298 48188 25304
rect 47950 21856 48006 21865
rect 47950 21791 48006 21800
rect 47964 21622 47992 21791
rect 47952 21616 48004 21622
rect 47952 21558 48004 21564
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48148 18834 48176 19071
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 48044 17604 48096 17610
rect 48044 17546 48096 17552
rect 47860 8016 47912 8022
rect 47860 7958 47912 7964
rect 48056 6866 48084 17546
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48148 16658 48176 17031
rect 48136 16652 48188 16658
rect 48136 16594 48188 16600
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48148 15570 48176 16351
rect 48136 15564 48188 15570
rect 48136 15506 48188 15512
rect 48136 13252 48188 13258
rect 48136 13194 48188 13200
rect 48148 12345 48176 13194
rect 48134 12336 48190 12345
rect 48134 12271 48190 12280
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 48136 7404 48188 7410
rect 48136 7346 48188 7352
rect 48148 6905 48176 7346
rect 48134 6896 48190 6905
rect 48044 6860 48096 6866
rect 48134 6831 48190 6840
rect 48044 6802 48096 6808
rect 47952 6112 48004 6118
rect 47952 6054 48004 6060
rect 47964 5302 47992 6054
rect 47952 5296 48004 5302
rect 47952 5238 48004 5244
rect 47768 5228 47820 5234
rect 47768 5170 47820 5176
rect 48056 5166 48084 6802
rect 48136 6316 48188 6322
rect 48136 6258 48188 6264
rect 48044 5160 48096 5166
rect 48044 5102 48096 5108
rect 47676 5024 47728 5030
rect 47676 4966 47728 4972
rect 47688 3602 47716 4966
rect 47768 4208 47820 4214
rect 48148 4185 48176 6258
rect 47768 4150 47820 4156
rect 48134 4176 48190 4185
rect 47676 3596 47728 3602
rect 47676 3538 47728 3544
rect 47780 3505 47808 4150
rect 48134 4111 48190 4120
rect 48320 4072 48372 4078
rect 48320 4014 48372 4020
rect 47766 3496 47822 3505
rect 47492 3460 47544 3466
rect 47766 3431 47822 3440
rect 47492 3402 47544 3408
rect 47768 3052 47820 3058
rect 47768 2994 47820 3000
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47032 2508 47084 2514
rect 47032 2450 47084 2456
rect 46296 2440 46348 2446
rect 46296 2382 46348 2388
rect 46388 2372 46440 2378
rect 46388 2314 46440 2320
rect 46400 800 46428 2314
rect 47044 800 47072 2450
rect 47688 800 47716 2926
rect 47780 1465 47808 2994
rect 47858 2952 47914 2961
rect 47858 2887 47914 2896
rect 47872 2854 47900 2887
rect 47860 2848 47912 2854
rect 47860 2790 47912 2796
rect 47952 2372 48004 2378
rect 47952 2314 48004 2320
rect 47766 1456 47822 1465
rect 47766 1391 47822 1400
rect 44180 536 44232 542
rect 44180 478 44232 484
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46846 776 46902 785
rect 46846 711 46902 720
rect 46860 542 46888 711
rect 46848 536 46900 542
rect 46848 478 46900 484
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 47964 105 47992 2314
rect 48332 800 48360 4014
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48976 800 49004 3402
rect 47950 96 48006 105
rect 47950 31 48006 40
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1398 47640 1454 47696
rect 3422 46960 3478 47016
rect 1398 42880 1454 42936
rect 2778 46280 2834 46336
rect 1858 41520 1914 41576
rect 1858 40160 1914 40216
rect 1398 33396 1400 33416
rect 1400 33396 1452 33416
rect 1452 33396 1454 33416
rect 1398 33360 1454 33396
rect 1582 35400 1638 35456
rect 1306 32680 1362 32736
rect 1858 32000 1914 32056
rect 1398 25236 1400 25256
rect 1400 25236 1452 25256
rect 1452 25236 1454 25256
rect 1398 25200 1454 25236
rect 1398 12280 1454 12336
rect 1858 23160 1914 23216
rect 2778 36760 2834 36816
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3514 44920 3570 44976
rect 3698 43560 3754 43616
rect 3514 39480 3570 39536
rect 3882 31320 3938 31376
rect 3974 28600 4030 28656
rect 3974 19760 4030 19816
rect 2226 19080 2282 19136
rect 3330 18400 3386 18456
rect 1858 17720 1914 17776
rect 3974 17040 4030 17096
rect 1858 16360 1914 16416
rect 2778 15000 2834 15056
rect 3974 13676 3976 13696
rect 3976 13676 4028 13696
rect 4028 13676 4030 13696
rect 3974 13640 4030 13676
rect 2778 10240 2834 10296
rect 3422 7520 3478 7576
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3514 6860 3570 6896
rect 3514 6840 3516 6860
rect 3516 6840 3568 6860
rect 3568 6840 3570 6860
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3974 3984 4030 4040
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3422 3440 3478 3496
rect 3238 1400 3294 1456
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3974 2352 4030 2408
rect 17314 31728 17370 31784
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 18418 32972 18474 33008
rect 18418 32952 18420 32972
rect 18420 32952 18472 32972
rect 18472 32952 18474 32972
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19062 32680 19118 32736
rect 18970 31728 19026 31784
rect 17130 3460 17186 3496
rect 17130 3440 17132 3460
rect 17132 3440 17184 3460
rect 17184 3440 17186 3460
rect 17314 3052 17370 3088
rect 17314 3032 17316 3052
rect 17316 3032 17368 3052
rect 17368 3032 17370 3052
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19522 32308 19524 32328
rect 19524 32308 19576 32328
rect 19576 32308 19578 32328
rect 19522 32272 19578 32308
rect 20166 32172 20168 32192
rect 20168 32172 20220 32192
rect 20220 32172 20222 32192
rect 20166 32136 20222 32172
rect 19706 32000 19762 32056
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19338 31220 19340 31240
rect 19340 31220 19392 31240
rect 19392 31220 19394 31240
rect 19338 31184 19394 31220
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 21546 32972 21602 33008
rect 21546 32952 21548 32972
rect 21548 32952 21600 32972
rect 21600 32952 21602 32972
rect 22190 32308 22192 32328
rect 22192 32308 22244 32328
rect 22244 32308 22246 32328
rect 22190 32272 22246 32308
rect 20810 30504 20866 30560
rect 22466 31320 22522 31376
rect 22374 30776 22430 30832
rect 22190 30368 22246 30424
rect 18234 3032 18290 3088
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20718 3188 20774 3224
rect 20718 3168 20720 3188
rect 20720 3168 20772 3188
rect 20772 3168 20774 3188
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 22834 31864 22890 31920
rect 22834 30368 22890 30424
rect 23294 35672 23350 35728
rect 23202 31320 23258 31376
rect 23110 31184 23166 31240
rect 23386 31864 23442 31920
rect 22190 3032 22246 3088
rect 22466 2916 22522 2952
rect 22466 2896 22468 2916
rect 22468 2896 22520 2916
rect 22520 2896 22522 2916
rect 22834 3168 22890 3224
rect 24950 32136 25006 32192
rect 25502 32000 25558 32056
rect 26422 32308 26424 32328
rect 26424 32308 26476 32328
rect 26476 32308 26478 32328
rect 26422 32272 26478 32308
rect 28354 35264 28410 35320
rect 24858 2896 24914 2952
rect 29090 35808 29146 35864
rect 28814 35672 28870 35728
rect 28998 35692 29054 35728
rect 28998 35672 29000 35692
rect 29000 35672 29052 35692
rect 29052 35672 29054 35692
rect 29090 35536 29146 35592
rect 28814 35400 28870 35456
rect 28722 35264 28778 35320
rect 29274 35808 29330 35864
rect 29550 35536 29606 35592
rect 30286 35672 30342 35728
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 29366 19236 29422 19272
rect 29366 19216 29368 19236
rect 29368 19216 29420 19236
rect 29420 19216 29422 19236
rect 30562 19236 30618 19272
rect 30562 19216 30564 19236
rect 30564 19216 30616 19236
rect 30616 19216 30618 19236
rect 29458 4020 29460 4040
rect 29460 4020 29512 4040
rect 29512 4020 29514 4040
rect 29458 3984 29514 4020
rect 31390 19780 31446 19816
rect 31390 19760 31392 19780
rect 31392 19760 31444 19780
rect 31444 19760 31446 19780
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 39026 2916 39082 2952
rect 39026 2896 39028 2916
rect 39028 2896 39080 2916
rect 39080 2896 39082 2916
rect 46846 47640 46902 47696
rect 46202 41132 46258 41168
rect 46202 41112 46204 41132
rect 46204 41112 46256 41132
rect 46256 41112 46258 41132
rect 46386 38956 46442 38992
rect 46386 38936 46388 38956
rect 46388 38936 46440 38956
rect 46440 38936 46442 38956
rect 47858 46280 47914 46336
rect 43810 3440 43866 3496
rect 45558 15680 45614 15736
rect 45558 8236 45560 8256
rect 45560 8236 45612 8256
rect 45612 8236 45614 8256
rect 45558 8200 45614 8236
rect 46018 22480 46074 22536
rect 46386 31320 46442 31376
rect 46294 29960 46350 30016
rect 46202 28600 46258 28656
rect 46294 26560 46350 26616
rect 46202 23840 46258 23896
rect 46754 25200 46810 25256
rect 46846 24520 46902 24576
rect 46846 23160 46902 23216
rect 46202 6196 46204 6216
rect 46204 6196 46256 6216
rect 46256 6196 46258 6216
rect 46202 6160 46258 6196
rect 2870 720 2926 776
rect 47030 18400 47086 18456
rect 47306 32000 47362 32056
rect 47306 29280 47362 29336
rect 47766 33360 47822 33416
rect 46846 9580 46902 9616
rect 46846 9560 46848 9580
rect 46848 9560 46900 9580
rect 46900 9560 46902 9580
rect 47306 7520 47362 7576
rect 47674 8880 47730 8936
rect 48134 45600 48190 45656
rect 48134 44512 48190 44568
rect 48134 41792 48190 41848
rect 48134 41384 48190 41440
rect 48134 40024 48190 40080
rect 48134 39072 48190 39128
rect 48134 37712 48190 37768
rect 48134 34720 48190 34776
rect 48134 34040 48190 34096
rect 48134 32680 48190 32736
rect 48134 27920 48190 27976
rect 48134 25880 48190 25936
rect 47950 21800 48006 21856
rect 48134 21120 48190 21176
rect 48134 19080 48190 19136
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 12280 48190 12336
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 48134 6840 48190 6896
rect 48134 4120 48190 4176
rect 47766 3440 47822 3496
rect 47858 2896 47914 2952
rect 47766 1400 47822 1456
rect 46846 720 46902 776
rect 47950 40 48006 96
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1393 47698 1459 47701
rect 0 47696 1459 47698
rect 0 47640 1398 47696
rect 1454 47640 1459 47696
rect 0 47638 1459 47640
rect 0 47548 800 47638
rect 1393 47635 1459 47638
rect 46841 47698 46907 47701
rect 49200 47698 50000 47788
rect 46841 47696 50000 47698
rect 46841 47640 46846 47696
rect 46902 47640 50000 47696
rect 46841 47638 50000 47640
rect 46841 47635 46907 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3417 47018 3483 47021
rect 0 47016 3483 47018
rect 0 46960 3422 47016
rect 3478 46960 3483 47016
rect 0 46958 3483 46960
rect 0 46868 800 46958
rect 3417 46955 3483 46958
rect 46054 46956 46060 47020
rect 46124 47018 46130 47020
rect 49200 47018 50000 47108
rect 46124 46958 50000 47018
rect 46124 46956 46130 46958
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46188 800 46278
rect 2773 46275 2839 46278
rect 47853 46338 47919 46341
rect 49200 46338 50000 46428
rect 47853 46336 50000 46338
rect 47853 46280 47858 46336
rect 47914 46280 50000 46336
rect 47853 46278 50000 46280
rect 47853 46275 47919 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3509 44978 3575 44981
rect 49200 44978 50000 45068
rect 0 44976 3575 44978
rect 0 44920 3514 44976
rect 3570 44920 3575 44976
rect 0 44918 3575 44920
rect 0 44828 800 44918
rect 3509 44915 3575 44918
rect 48270 44918 50000 44978
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 48129 44570 48195 44573
rect 48270 44570 48330 44918
rect 49200 44828 50000 44918
rect 48129 44568 48330 44570
rect 48129 44512 48134 44568
rect 48190 44512 48330 44568
rect 48129 44510 48330 44512
rect 48129 44507 48195 44510
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3693 43618 3759 43621
rect 0 43616 3759 43618
rect 0 43560 3698 43616
rect 3754 43560 3759 43616
rect 0 43558 3759 43560
rect 0 43468 800 43558
rect 3693 43555 3759 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42788 800 42878
rect 1393 42875 1459 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 49200 42258 50000 42348
rect 48270 42198 50000 42258
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 48129 41850 48195 41853
rect 48270 41850 48330 42198
rect 49200 42108 50000 42198
rect 48129 41848 48330 41850
rect 48129 41792 48134 41848
rect 48190 41792 48330 41848
rect 48129 41790 48330 41792
rect 48129 41787 48195 41790
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 49200 41578 50000 41668
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48270 41518 50000 41578
rect 48129 41442 48195 41445
rect 48270 41442 48330 41518
rect 48129 41440 48330 41442
rect 48129 41384 48134 41440
rect 48190 41384 48330 41440
rect 49200 41428 50000 41518
rect 48129 41382 48330 41384
rect 48129 41379 48195 41382
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 46197 41170 46263 41173
rect 46197 41168 48330 41170
rect 46197 41112 46202 41168
rect 46258 41112 48330 41168
rect 46197 41110 48330 41112
rect 46197 41107 46263 41110
rect 0 40748 800 40988
rect 48270 40898 48330 41110
rect 49200 40898 50000 40988
rect 48270 40838 50000 40898
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1853 40218 1919 40221
rect 49200 40218 50000 40308
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40068 800 40158
rect 1853 40155 1919 40158
rect 48270 40158 50000 40218
rect 48129 40082 48195 40085
rect 48270 40082 48330 40158
rect 48129 40080 48330 40082
rect 48129 40024 48134 40080
rect 48190 40024 48330 40080
rect 49200 40068 50000 40158
rect 48129 40022 48330 40024
rect 48129 40019 48195 40022
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3509 39538 3575 39541
rect 49200 39538 50000 39628
rect 0 39536 3575 39538
rect 0 39480 3514 39536
rect 3570 39480 3575 39536
rect 0 39478 3575 39480
rect 0 39388 800 39478
rect 3509 39475 3575 39478
rect 48270 39478 50000 39538
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 48129 39130 48195 39133
rect 48270 39130 48330 39478
rect 49200 39388 50000 39478
rect 48129 39128 48330 39130
rect 48129 39072 48134 39128
rect 48190 39072 48330 39128
rect 48129 39070 48330 39072
rect 48129 39067 48195 39070
rect 46381 38994 46447 38997
rect 46381 38992 48330 38994
rect 0 38708 800 38948
rect 46381 38936 46386 38992
rect 46442 38936 48330 38992
rect 46381 38934 48330 38936
rect 46381 38931 46447 38934
rect 48270 38858 48330 38934
rect 49200 38858 50000 38948
rect 48270 38798 50000 38858
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 49200 38178 50000 38268
rect 48270 38118 50000 38178
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 48129 37770 48195 37773
rect 48270 37770 48330 38118
rect 49200 38028 50000 38118
rect 48129 37768 48330 37770
rect 48129 37712 48134 37768
rect 48190 37712 48330 37768
rect 48129 37710 48330 37712
rect 48129 37707 48195 37710
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 29085 35866 29151 35869
rect 29269 35866 29335 35869
rect 27570 35864 29335 35866
rect 27570 35808 29090 35864
rect 29146 35808 29274 35864
rect 29330 35808 29335 35864
rect 27570 35806 29335 35808
rect 23289 35730 23355 35733
rect 27570 35730 27630 35806
rect 29085 35803 29151 35806
rect 29269 35803 29335 35806
rect 28809 35730 28875 35733
rect 23289 35728 27630 35730
rect 23289 35672 23294 35728
rect 23350 35672 27630 35728
rect 23289 35670 27630 35672
rect 28766 35728 28875 35730
rect 28766 35672 28814 35728
rect 28870 35672 28875 35728
rect 23289 35667 23355 35670
rect 28766 35667 28875 35672
rect 28993 35730 29059 35733
rect 30281 35730 30347 35733
rect 28993 35728 30347 35730
rect 28993 35672 28998 35728
rect 29054 35672 30286 35728
rect 30342 35672 30347 35728
rect 28993 35670 30347 35672
rect 28993 35667 29059 35670
rect 30281 35667 30347 35670
rect 0 35458 800 35548
rect 28766 35461 28826 35667
rect 29085 35594 29151 35597
rect 29545 35594 29611 35597
rect 29085 35592 29611 35594
rect 29085 35536 29090 35592
rect 29146 35536 29550 35592
rect 29606 35536 29611 35592
rect 29085 35534 29611 35536
rect 29085 35531 29151 35534
rect 29545 35531 29611 35534
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 28766 35456 28875 35461
rect 28766 35400 28814 35456
rect 28870 35400 28875 35456
rect 28766 35398 28875 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 28809 35395 28875 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 28349 35322 28415 35325
rect 28717 35322 28783 35325
rect 28349 35320 28783 35322
rect 28349 35264 28354 35320
rect 28410 35264 28722 35320
rect 28778 35264 28783 35320
rect 28349 35262 28783 35264
rect 28349 35259 28415 35262
rect 28717 35259 28783 35262
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 48129 34098 48195 34101
rect 49200 34098 50000 34188
rect 48129 34096 50000 34098
rect 48129 34040 48134 34096
rect 48190 34040 50000 34096
rect 48129 34038 50000 34040
rect 48129 34035 48195 34038
rect 49200 33948 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 47761 33418 47827 33421
rect 49200 33418 50000 33508
rect 47761 33416 50000 33418
rect 47761 33360 47766 33416
rect 47822 33360 50000 33416
rect 47761 33358 50000 33360
rect 47761 33355 47827 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 18413 33010 18479 33013
rect 21541 33010 21607 33013
rect 18413 33008 21607 33010
rect 18413 32952 18418 33008
rect 18474 32952 21546 33008
rect 21602 32952 21607 33008
rect 18413 32950 21607 32952
rect 18413 32947 18479 32950
rect 21541 32947 21607 32950
rect 0 32738 800 32828
rect 1301 32738 1367 32741
rect 19057 32738 19123 32741
rect 0 32736 1367 32738
rect 0 32680 1306 32736
rect 1362 32680 1367 32736
rect 0 32678 1367 32680
rect 0 32588 800 32678
rect 1301 32675 1367 32678
rect 19014 32736 19123 32738
rect 19014 32680 19062 32736
rect 19118 32680 19123 32736
rect 19014 32675 19123 32680
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 1853 32058 1919 32061
rect 0 32056 1919 32058
rect 0 32000 1858 32056
rect 1914 32000 1919 32056
rect 0 31998 1919 32000
rect 0 31908 800 31998
rect 1853 31995 1919 31998
rect 19014 31789 19074 32675
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 49200 32588 50000 32678
rect 19517 32330 19583 32333
rect 22185 32330 22251 32333
rect 26417 32330 26483 32333
rect 19517 32328 26483 32330
rect 19517 32272 19522 32328
rect 19578 32272 22190 32328
rect 22246 32272 26422 32328
rect 26478 32272 26483 32328
rect 19517 32270 26483 32272
rect 19517 32267 19583 32270
rect 22185 32267 22251 32270
rect 26417 32267 26483 32270
rect 20161 32194 20227 32197
rect 24945 32194 25011 32197
rect 20161 32192 25011 32194
rect 20161 32136 20166 32192
rect 20222 32136 24950 32192
rect 25006 32136 25011 32192
rect 20161 32134 25011 32136
rect 20161 32131 20227 32134
rect 24945 32131 25011 32134
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19701 32058 19767 32061
rect 25497 32058 25563 32061
rect 19701 32056 25563 32058
rect 19701 32000 19706 32056
rect 19762 32000 25502 32056
rect 25558 32000 25563 32056
rect 19701 31998 25563 32000
rect 19701 31995 19767 31998
rect 25497 31995 25563 31998
rect 47301 32058 47367 32061
rect 49200 32058 50000 32148
rect 47301 32056 50000 32058
rect 47301 32000 47306 32056
rect 47362 32000 50000 32056
rect 47301 31998 50000 32000
rect 47301 31995 47367 31998
rect 22829 31922 22895 31925
rect 23381 31922 23447 31925
rect 22829 31920 23447 31922
rect 22829 31864 22834 31920
rect 22890 31864 23386 31920
rect 23442 31864 23447 31920
rect 49200 31908 50000 31998
rect 22829 31862 23447 31864
rect 22829 31859 22895 31862
rect 23381 31859 23447 31862
rect 17309 31788 17375 31789
rect 17309 31784 17356 31788
rect 17420 31786 17426 31788
rect 17309 31728 17314 31784
rect 17309 31724 17356 31728
rect 17420 31726 17466 31786
rect 18965 31784 19074 31789
rect 18965 31728 18970 31784
rect 19026 31728 19074 31784
rect 18965 31726 19074 31728
rect 17420 31724 17426 31726
rect 17309 31723 17375 31724
rect 18965 31723 19031 31726
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3877 31378 3943 31381
rect 0 31376 3943 31378
rect 0 31320 3882 31376
rect 3938 31320 3943 31376
rect 0 31318 3943 31320
rect 0 31228 800 31318
rect 3877 31315 3943 31318
rect 22461 31378 22527 31381
rect 23197 31378 23263 31381
rect 22461 31376 23263 31378
rect 22461 31320 22466 31376
rect 22522 31320 23202 31376
rect 23258 31320 23263 31376
rect 22461 31318 23263 31320
rect 22461 31315 22527 31318
rect 23197 31315 23263 31318
rect 46381 31378 46447 31381
rect 49200 31378 50000 31468
rect 46381 31376 50000 31378
rect 46381 31320 46386 31376
rect 46442 31320 50000 31376
rect 46381 31318 50000 31320
rect 46381 31315 46447 31318
rect 19333 31242 19399 31245
rect 23105 31242 23171 31245
rect 19333 31240 23171 31242
rect 19333 31184 19338 31240
rect 19394 31184 23110 31240
rect 23166 31184 23171 31240
rect 49200 31228 50000 31318
rect 19333 31182 23171 31184
rect 19333 31179 19399 31182
rect 23105 31179 23171 31182
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 22369 30834 22435 30837
rect 22050 30832 22435 30834
rect 0 30548 800 30788
rect 22050 30776 22374 30832
rect 22430 30776 22435 30832
rect 22050 30774 22435 30776
rect 20805 30562 20871 30565
rect 22050 30562 22110 30774
rect 22369 30771 22435 30774
rect 20805 30560 22110 30562
rect 20805 30504 20810 30560
rect 20866 30504 22110 30560
rect 49200 30548 50000 30788
rect 20805 30502 22110 30504
rect 20805 30499 20871 30502
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 22185 30426 22251 30429
rect 22829 30426 22895 30429
rect 22185 30424 22895 30426
rect 22185 30368 22190 30424
rect 22246 30368 22834 30424
rect 22890 30368 22895 30424
rect 22185 30366 22895 30368
rect 22185 30363 22251 30366
rect 22829 30363 22895 30366
rect 0 29868 800 30108
rect 46289 30018 46355 30021
rect 49200 30018 50000 30108
rect 46289 30016 50000 30018
rect 46289 29960 46294 30016
rect 46350 29960 50000 30016
rect 46289 29958 50000 29960
rect 46289 29955 46355 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 47301 29338 47367 29341
rect 49200 29338 50000 29428
rect 47301 29336 50000 29338
rect 47301 29280 47306 29336
rect 47362 29280 50000 29336
rect 47301 29278 50000 29280
rect 47301 29275 47367 29278
rect 49200 29188 50000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3969 28658 4035 28661
rect 0 28656 4035 28658
rect 0 28600 3974 28656
rect 4030 28600 4035 28656
rect 0 28598 4035 28600
rect 0 28508 800 28598
rect 3969 28595 4035 28598
rect 46197 28658 46263 28661
rect 49200 28658 50000 28748
rect 46197 28656 50000 28658
rect 46197 28600 46202 28656
rect 46258 28600 50000 28656
rect 46197 28598 50000 28600
rect 46197 28595 46263 28598
rect 49200 28508 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 49200 27828 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 46289 26618 46355 26621
rect 49200 26618 50000 26708
rect 46289 26616 50000 26618
rect 46289 26560 46294 26616
rect 46350 26560 50000 26616
rect 46289 26558 50000 26560
rect 46289 26555 46355 26558
rect 49200 26468 50000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 48129 25938 48195 25941
rect 49200 25938 50000 26028
rect 48129 25936 50000 25938
rect 48129 25880 48134 25936
rect 48190 25880 50000 25936
rect 48129 25878 50000 25880
rect 48129 25875 48195 25878
rect 49200 25788 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25108 800 25198
rect 1393 25195 1459 25198
rect 46749 25258 46815 25261
rect 49200 25258 50000 25348
rect 46749 25256 50000 25258
rect 46749 25200 46754 25256
rect 46810 25200 50000 25256
rect 46749 25198 50000 25200
rect 46749 25195 46815 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24428 800 24668
rect 46841 24578 46907 24581
rect 49200 24578 50000 24668
rect 46841 24576 50000 24578
rect 46841 24520 46846 24576
rect 46902 24520 50000 24576
rect 46841 24518 50000 24520
rect 46841 24515 46907 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 46197 23898 46263 23901
rect 49200 23898 50000 23988
rect 46197 23896 50000 23898
rect 46197 23840 46202 23896
rect 46258 23840 50000 23896
rect 46197 23838 50000 23840
rect 46197 23835 46263 23838
rect 49200 23748 50000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23068 800 23158
rect 1853 23155 1919 23158
rect 46841 23218 46907 23221
rect 49200 23218 50000 23308
rect 46841 23216 50000 23218
rect 46841 23160 46846 23216
rect 46902 23160 50000 23216
rect 46841 23158 50000 23160
rect 46841 23155 46907 23158
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 46013 22538 46079 22541
rect 49200 22538 50000 22628
rect 46013 22536 50000 22538
rect 46013 22480 46018 22536
rect 46074 22480 50000 22536
rect 46013 22478 50000 22480
rect 46013 22475 46079 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21708 800 21948
rect 47945 21858 48011 21861
rect 49200 21858 50000 21948
rect 47945 21856 50000 21858
rect 47945 21800 47950 21856
rect 48006 21800 50000 21856
rect 47945 21798 50000 21800
rect 47945 21795 48011 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 49200 21028 50000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19668 800 19758
rect 3969 19755 4035 19758
rect 31385 19818 31451 19821
rect 46054 19818 46060 19820
rect 31385 19816 46060 19818
rect 31385 19760 31390 19816
rect 31446 19760 46060 19816
rect 31385 19758 46060 19760
rect 31385 19755 31451 19758
rect 46054 19756 46060 19758
rect 46124 19756 46130 19820
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 29361 19274 29427 19277
rect 30557 19274 30623 19277
rect 29361 19272 30623 19274
rect 0 19138 800 19228
rect 29361 19216 29366 19272
rect 29422 19216 30562 19272
rect 30618 19216 30623 19272
rect 29361 19214 30623 19216
rect 29361 19211 29427 19214
rect 30557 19211 30623 19214
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3325 18458 3391 18461
rect 0 18456 3391 18458
rect 0 18400 3330 18456
rect 3386 18400 3391 18456
rect 0 18398 3391 18400
rect 0 18308 800 18398
rect 3325 18395 3391 18398
rect 47025 18458 47091 18461
rect 49200 18458 50000 18548
rect 47025 18456 50000 18458
rect 47025 18400 47030 18456
rect 47086 18400 50000 18456
rect 47025 18398 50000 18400
rect 47025 18395 47091 18398
rect 49200 18308 50000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1853 17778 1919 17781
rect 0 17776 1919 17778
rect 0 17720 1858 17776
rect 1914 17720 1919 17776
rect 0 17718 1919 17720
rect 0 17628 800 17718
rect 1853 17715 1919 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3969 17098 4035 17101
rect 0 17096 4035 17098
rect 0 17040 3974 17096
rect 4030 17040 4035 17096
rect 0 17038 4035 17040
rect 0 16948 800 17038
rect 3969 17035 4035 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16268 800 16358
rect 1853 16355 1919 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16508
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 45553 15738 45619 15741
rect 49200 15738 50000 15828
rect 45553 15736 50000 15738
rect 45553 15680 45558 15736
rect 45614 15680 50000 15736
rect 45553 15678 50000 15680
rect 45553 15675 45619 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3969 13698 4035 13701
rect 0 13696 4035 13698
rect 0 13640 3974 13696
rect 4030 13640 4035 13696
rect 0 13638 4035 13640
rect 0 13548 800 13638
rect 3969 13635 4035 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 2773 10298 2839 10301
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 0 10148 800 10238
rect 2773 10235 2839 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 46841 9618 46907 9621
rect 49200 9618 50000 9708
rect 46841 9616 50000 9618
rect 46841 9560 46846 9616
rect 46902 9560 50000 9616
rect 46841 9558 50000 9560
rect 46841 9555 46907 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47669 8938 47735 8941
rect 49200 8938 50000 9028
rect 47669 8936 50000 8938
rect 47669 8880 47674 8936
rect 47730 8880 50000 8936
rect 47669 8878 50000 8880
rect 47669 8875 47735 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 45553 8258 45619 8261
rect 49200 8258 50000 8348
rect 45553 8256 50000 8258
rect 45553 8200 45558 8256
rect 45614 8200 50000 8256
rect 45553 8198 50000 8200
rect 45553 8195 45619 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3417 7578 3483 7581
rect 0 7576 3483 7578
rect 0 7520 3422 7576
rect 3478 7520 3483 7576
rect 0 7518 3483 7520
rect 0 7428 800 7518
rect 3417 7515 3483 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 3509 6898 3575 6901
rect 0 6896 3575 6898
rect 0 6840 3514 6896
rect 3570 6840 3575 6896
rect 0 6838 3575 6840
rect 0 6748 800 6838
rect 3509 6835 3575 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 46197 6218 46263 6221
rect 49200 6218 50000 6308
rect 46197 6216 50000 6218
rect 46197 6160 46202 6216
rect 46258 6160 50000 6216
rect 46197 6158 50000 6160
rect 46197 6155 46263 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 48129 4178 48195 4181
rect 49200 4178 50000 4268
rect 48129 4176 50000 4178
rect 48129 4120 48134 4176
rect 48190 4120 50000 4176
rect 48129 4118 50000 4120
rect 48129 4115 48195 4118
rect 3969 4042 4035 4045
rect 29453 4042 29519 4045
rect 3969 4040 29519 4042
rect 3969 3984 3974 4040
rect 4030 3984 29458 4040
rect 29514 3984 29519 4040
rect 49200 4028 50000 4118
rect 3969 3982 29519 3984
rect 3969 3979 4035 3982
rect 29453 3979 29519 3982
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3588
rect 3417 3498 3483 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3348 800 3438
rect 3417 3435 3483 3438
rect 17125 3498 17191 3501
rect 43805 3498 43871 3501
rect 17125 3496 43871 3498
rect 17125 3440 17130 3496
rect 17186 3440 43810 3496
rect 43866 3440 43871 3496
rect 17125 3438 43871 3440
rect 17125 3435 17191 3438
rect 43805 3435 43871 3438
rect 47761 3498 47827 3501
rect 49200 3498 50000 3588
rect 47761 3496 50000 3498
rect 47761 3440 47766 3496
rect 47822 3440 50000 3496
rect 47761 3438 50000 3440
rect 47761 3435 47827 3438
rect 49200 3348 50000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 20713 3226 20779 3229
rect 22829 3226 22895 3229
rect 20713 3224 22895 3226
rect 20713 3168 20718 3224
rect 20774 3168 22834 3224
rect 22890 3168 22895 3224
rect 20713 3166 22895 3168
rect 20713 3163 20779 3166
rect 22829 3163 22895 3166
rect 17309 3090 17375 3093
rect 18229 3090 18295 3093
rect 22185 3090 22251 3093
rect 17309 3088 22251 3090
rect 17309 3032 17314 3088
rect 17370 3032 18234 3088
rect 18290 3032 22190 3088
rect 22246 3032 22251 3088
rect 17309 3030 22251 3032
rect 17309 3027 17375 3030
rect 18229 3027 18295 3030
rect 22185 3027 22251 3030
rect 22461 2954 22527 2957
rect 24853 2954 24919 2957
rect 22461 2952 24919 2954
rect 0 2668 800 2908
rect 22461 2896 22466 2952
rect 22522 2896 24858 2952
rect 24914 2896 24919 2952
rect 22461 2894 24919 2896
rect 22461 2891 22527 2894
rect 24853 2891 24919 2894
rect 39021 2954 39087 2957
rect 47853 2954 47919 2957
rect 39021 2952 47919 2954
rect 39021 2896 39026 2952
rect 39082 2896 47858 2952
rect 47914 2896 47919 2952
rect 39021 2894 47919 2896
rect 39021 2891 39087 2894
rect 47853 2891 47919 2894
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 3969 2410 4035 2413
rect 17350 2410 17356 2412
rect 3969 2408 17356 2410
rect 3969 2352 3974 2408
rect 4030 2352 17356 2408
rect 3969 2350 17356 2352
rect 3969 2347 4035 2350
rect 17350 2348 17356 2350
rect 17420 2348 17426 2412
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3233 1458 3299 1461
rect 0 1456 3299 1458
rect 0 1400 3238 1456
rect 3294 1400 3299 1456
rect 0 1398 3299 1400
rect 0 1308 800 1398
rect 3233 1395 3299 1398
rect 47761 1458 47827 1461
rect 49200 1458 50000 1548
rect 47761 1456 50000 1458
rect 47761 1400 47766 1456
rect 47822 1400 50000 1456
rect 47761 1398 50000 1400
rect 47761 1395 47827 1398
rect 49200 1308 50000 1398
rect 0 778 800 868
rect 2865 778 2931 781
rect 0 776 2931 778
rect 0 720 2870 776
rect 2926 720 2931 776
rect 0 718 2931 720
rect 0 628 800 718
rect 2865 715 2931 718
rect 46841 778 46907 781
rect 49200 778 50000 868
rect 46841 776 50000 778
rect 46841 720 46846 776
rect 46902 720 50000 776
rect 46841 718 50000 720
rect 46841 715 46907 718
rect 49200 628 50000 718
rect 47945 98 48011 101
rect 49200 98 50000 188
rect 47945 96 50000 98
rect 47945 40 47950 96
rect 48006 40 50000 96
rect 47945 38 50000 40
rect 47945 35 48011 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 46060 46956 46124 47020
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 17356 31784 17420 31788
rect 17356 31728 17370 31784
rect 17370 31728 17420 31784
rect 17356 31724 17420 31728
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 46060 19756 46124 19820
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 17356 2348 17420 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 17355 31788 17421 31789
rect 17355 31724 17356 31788
rect 17420 31724 17421 31788
rect 17355 31723 17421 31724
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 17358 2413 17418 31723
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 17355 2412 17421 2413
rect 17355 2348 17356 2412
rect 17420 2348 17421 2412
rect 17355 2347 17421 2348
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 46059 47020 46125 47021
rect 46059 46956 46060 47020
rect 46124 46956 46125 47020
rect 46059 46955 46125 46956
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 46062 19821 46122 46955
rect 46059 19820 46125 19821
rect 46059 19756 46060 19820
rect 46124 19756 46125 19820
rect 46059 19755 46125 19756
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18032 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_95 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1644511149
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1644511149
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1644511149
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_200
timestamp 1644511149
transform 1 0 19504 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1644511149
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1644511149
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_291 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1644511149
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_412
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1644511149
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_464
timestamp 1644511149
transform 1 0 43792 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_63
timestamp 1644511149
transform 1 0 6900 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_92
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_99
timestamp 1644511149
transform 1 0 10212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1644511149
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_185
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_199
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp 1644511149
transform 1 0 20884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_289
timestamp 1644511149
transform 1 0 27692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_301
timestamp 1644511149
transform 1 0 28796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_313
timestamp 1644511149
transform 1 0 29900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_325
timestamp 1644511149
transform 1 0 31004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1644511149
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_345
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_379
timestamp 1644511149
transform 1 0 35972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1644511149
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_399
timestamp 1644511149
transform 1 0 37812 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1644511149
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_415
timestamp 1644511149
transform 1 0 39284 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_440
timestamp 1644511149
transform 1 0 41584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_470
timestamp 1644511149
transform 1 0 44344 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1644511149
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_117
timestamp 1644511149
transform 1 0 11868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_122
timestamp 1644511149
transform 1 0 12328 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_130
timestamp 1644511149
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_152
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1644511149
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_179
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_183
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1644511149
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1644511149
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_216
timestamp 1644511149
transform 1 0 20976 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_223
timestamp 1644511149
transform 1 0 21620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_232
timestamp 1644511149
transform 1 0 22448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_239
timestamp 1644511149
transform 1 0 23092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_246
timestamp 1644511149
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_259
timestamp 1644511149
transform 1 0 24932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_266
timestamp 1644511149
transform 1 0 25576 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_278
timestamp 1644511149
transform 1 0 26680 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_290
timestamp 1644511149
transform 1 0 27784 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1644511149
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_330
timestamp 1644511149
transform 1 0 31464 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1644511149
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_346
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_350
timestamp 1644511149
transform 1 0 33304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_399
timestamp 1644511149
transform 1 0 37812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_411
timestamp 1644511149
transform 1 0 38916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1644511149
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1644511149
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_63
timestamp 1644511149
transform 1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_67
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_71
timestamp 1644511149
transform 1 0 7636 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_80
timestamp 1644511149
transform 1 0 8464 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_91
timestamp 1644511149
transform 1 0 9476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 1644511149
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_116
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_128
timestamp 1644511149
transform 1 0 12880 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_188
timestamp 1644511149
transform 1 0 18400 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_194
timestamp 1644511149
transform 1 0 18952 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_198
timestamp 1644511149
transform 1 0 19320 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_212
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1644511149
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_239
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_246
timestamp 1644511149
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_253
timestamp 1644511149
transform 1 0 24380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_265
timestamp 1644511149
transform 1 0 25484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1644511149
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_421
timestamp 1644511149
transform 1 0 39836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_425
timestamp 1644511149
transform 1 0 40204 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_437
timestamp 1644511149
transform 1 0 41308 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_445
timestamp 1644511149
transform 1 0 42044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_456
timestamp 1644511149
transform 1 0 43056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_460
timestamp 1644511149
transform 1 0 43424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_482
timestamp 1644511149
transform 1 0 45448 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_74
timestamp 1644511149
transform 1 0 7912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1644511149
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_201
timestamp 1644511149
transform 1 0 19596 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_205
timestamp 1644511149
transform 1 0 19964 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_212
timestamp 1644511149
transform 1 0 20608 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1644511149
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_226
timestamp 1644511149
transform 1 0 21896 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_240
timestamp 1644511149
transform 1 0 23184 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_451
timestamp 1644511149
transform 1 0 42596 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_455
timestamp 1644511149
transform 1 0 42964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_467
timestamp 1644511149
transform 1 0 44068 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_481
timestamp 1644511149
transform 1 0 45356 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_485
timestamp 1644511149
transform 1 0 45724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_510
timestamp 1644511149
transform 1 0 48024 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1644511149
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_508
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1644511149
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_489
timestamp 1644511149
transform 1 0 46092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_500
timestamp 1644511149
transform 1 0 47104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_497
timestamp 1644511149
transform 1 0 46828 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_511
timestamp 1644511149
transform 1 0 48116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_515
timestamp 1644511149
transform 1 0 48484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1644511149
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_500
timestamp 1644511149
transform 1 0 47104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_508
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_183
timestamp 1644511149
transform 1 0 17940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1644511149
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_203
timestamp 1644511149
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1644511149
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_184
timestamp 1644511149
transform 1 0 18032 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1644511149
transform 1 0 19044 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1644511149
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_495
timestamp 1644511149
transform 1 0 46644 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_499
timestamp 1644511149
transform 1 0 47012 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_511
timestamp 1644511149
transform 1 0 48116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_515
timestamp 1644511149
transform 1 0 48484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1644511149
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_202
timestamp 1644511149
transform 1 0 19688 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1644511149
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1644511149
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1644511149
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_157
timestamp 1644511149
transform 1 0 15548 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_179
timestamp 1644511149
transform 1 0 17572 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1644511149
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_201
timestamp 1644511149
transform 1 0 19596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_205
timestamp 1644511149
transform 1 0 19964 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1644511149
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_178
timestamp 1644511149
transform 1 0 17480 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1644511149
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_216
timestamp 1644511149
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_508
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_147
timestamp 1644511149
transform 1 0 14628 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_161
timestamp 1644511149
transform 1 0 15916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_168
timestamp 1644511149
transform 1 0 16560 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_174
timestamp 1644511149
transform 1 0 17112 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1644511149
transform 1 0 17664 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_200
timestamp 1644511149
transform 1 0 19504 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_212
timestamp 1644511149
transform 1 0 20608 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_224
timestamp 1644511149
transform 1 0 21712 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_236
timestamp 1644511149
transform 1 0 22816 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_152
timestamp 1644511149
transform 1 0 15088 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1644511149
transform 1 0 17572 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_186
timestamp 1644511149
transform 1 0 18216 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_198
timestamp 1644511149
transform 1 0 19320 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_210
timestamp 1644511149
transform 1 0 20424 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1644511149
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1644511149
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_145
timestamp 1644511149
transform 1 0 14444 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_152
timestamp 1644511149
transform 1 0 15088 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1644511149
transform 1 0 15640 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1644511149
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_187
timestamp 1644511149
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_200
timestamp 1644511149
transform 1 0 19504 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_208
timestamp 1644511149
transform 1 0 20240 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_214
timestamp 1644511149
transform 1 0 20792 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_226
timestamp 1644511149
transform 1 0 21896 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_238
timestamp 1644511149
transform 1 0 23000 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1644511149
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_512
timestamp 1644511149
transform 1 0 48208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_121
timestamp 1644511149
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_131
timestamp 1644511149
transform 1 0 13156 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_156
timestamp 1644511149
transform 1 0 15456 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_195
timestamp 1644511149
transform 1 0 19044 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1644511149
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_500
timestamp 1644511149
transform 1 0 47104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_178
timestamp 1644511149
transform 1 0 17480 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_184
timestamp 1644511149
transform 1 0 18032 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_204
timestamp 1644511149
transform 1 0 19872 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_214
timestamp 1644511149
transform 1 0 20792 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_226
timestamp 1644511149
transform 1 0 21896 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_238
timestamp 1644511149
transform 1 0 23000 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1644511149
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_73
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_77
timestamp 1644511149
transform 1 0 8188 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_102
timestamp 1644511149
transform 1 0 10488 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1644511149
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_117
timestamp 1644511149
transform 1 0 11868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_129
timestamp 1644511149
transform 1 0 12972 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_142
timestamp 1644511149
transform 1 0 14168 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_150
timestamp 1644511149
transform 1 0 14904 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1644511149
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_162
timestamp 1644511149
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_185
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_191
timestamp 1644511149
transform 1 0 18676 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_199
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_229
timestamp 1644511149
transform 1 0 22172 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_241
timestamp 1644511149
transform 1 0 23276 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_253
timestamp 1644511149
transform 1 0 24380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_265
timestamp 1644511149
transform 1 0 25484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1644511149
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_310
timestamp 1644511149
transform 1 0 29624 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1644511149
transform 1 0 30728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1644511149
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_145
timestamp 1644511149
transform 1 0 14444 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_176
timestamp 1644511149
transform 1 0 17296 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_212
timestamp 1644511149
transform 1 0 20608 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_276
timestamp 1644511149
transform 1 0 26496 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1644511149
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_495
timestamp 1644511149
transform 1 0 46644 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_499
timestamp 1644511149
transform 1 0 47012 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_506
timestamp 1644511149
transform 1 0 47656 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_514
timestamp 1644511149
transform 1 0 48392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_11
timestamp 1644511149
transform 1 0 2116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_23
timestamp 1644511149
transform 1 0 3220 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_35
timestamp 1644511149
transform 1 0 4324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1644511149
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_148
timestamp 1644511149
transform 1 0 14720 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_155
timestamp 1644511149
transform 1 0 15364 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_190
timestamp 1644511149
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_201
timestamp 1644511149
transform 1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1644511149
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_212
timestamp 1644511149
transform 1 0 20608 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_231
timestamp 1644511149
transform 1 0 22356 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_255
timestamp 1644511149
transform 1 0 24564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_263
timestamp 1644511149
transform 1 0 25300 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_267
timestamp 1644511149
transform 1 0 25668 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 1644511149
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1644511149
transform 1 0 27416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_295
timestamp 1644511149
transform 1 0 28244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_302
timestamp 1644511149
transform 1 0 28888 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_314
timestamp 1644511149
transform 1 0 29992 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_326
timestamp 1644511149
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1644511149
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_510
timestamp 1644511149
transform 1 0 48024 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1644511149
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_106
timestamp 1644511149
transform 1 0 10856 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_118
timestamp 1644511149
transform 1 0 11960 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_127
timestamp 1644511149
transform 1 0 12788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_134
timestamp 1644511149
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_146
timestamp 1644511149
transform 1 0 14536 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_159
timestamp 1644511149
transform 1 0 15732 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_171
timestamp 1644511149
transform 1 0 16836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_175
timestamp 1644511149
transform 1 0 17204 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_183
timestamp 1644511149
transform 1 0 17940 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1644511149
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1644511149
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_218
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_226
timestamp 1644511149
transform 1 0 21896 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_232
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_240
timestamp 1644511149
transform 1 0 23184 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_244
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_256
timestamp 1644511149
transform 1 0 24656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_268
timestamp 1644511149
transform 1 0 25760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_276
timestamp 1644511149
transform 1 0 26496 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_285
timestamp 1644511149
transform 1 0 27324 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_291
timestamp 1644511149
transform 1 0 27876 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1644511149
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1644511149
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_483
timestamp 1644511149
transform 1 0 45540 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_487
timestamp 1644511149
transform 1 0 45908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_89
timestamp 1644511149
transform 1 0 9292 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_101
timestamp 1644511149
transform 1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_133
timestamp 1644511149
transform 1 0 13340 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_146
timestamp 1644511149
transform 1 0 14536 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_158
timestamp 1644511149
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1644511149
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1644511149
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_180
timestamp 1644511149
transform 1 0 17664 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_209
timestamp 1644511149
transform 1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_241
timestamp 1644511149
transform 1 0 23276 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_253
timestamp 1644511149
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_265
timestamp 1644511149
transform 1 0 25484 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_288
timestamp 1644511149
transform 1 0 27600 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_300
timestamp 1644511149
transform 1 0 28704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_306
timestamp 1644511149
transform 1 0 29256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_320
timestamp 1644511149
transform 1 0 30544 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_426
timestamp 1644511149
transform 1 0 40296 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_438
timestamp 1644511149
transform 1 0 41400 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1644511149
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_483
timestamp 1644511149
transform 1 0 45540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_500
timestamp 1644511149
transform 1 0 47104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1644511149
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_118
timestamp 1644511149
transform 1 0 11960 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_126
timestamp 1644511149
transform 1 0 12696 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_148
timestamp 1644511149
transform 1 0 14720 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_160
timestamp 1644511149
transform 1 0 15824 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1644511149
transform 1 0 16744 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_174
timestamp 1644511149
transform 1 0 17112 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_186
timestamp 1644511149
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1644511149
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_218
timestamp 1644511149
transform 1 0 21160 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_266
timestamp 1644511149
transform 1 0 25576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_273
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_282
timestamp 1644511149
transform 1 0 27048 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_291
timestamp 1644511149
transform 1 0 27876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_299
timestamp 1644511149
transform 1 0 28612 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1644511149
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_330
timestamp 1644511149
transform 1 0 31464 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_342
timestamp 1644511149
transform 1 0 32568 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_354
timestamp 1644511149
transform 1 0 33672 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1644511149
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1644511149
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_485
timestamp 1644511149
transform 1 0 45724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_502
timestamp 1644511149
transform 1 0 47288 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_509
timestamp 1644511149
transform 1 0 47932 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_515
timestamp 1644511149
transform 1 0 48484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_91
timestamp 1644511149
transform 1 0 9476 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_95
timestamp 1644511149
transform 1 0 9844 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_99
timestamp 1644511149
transform 1 0 10212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1644511149
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_124
timestamp 1644511149
transform 1 0 12512 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_132
timestamp 1644511149
transform 1 0 13248 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1644511149
transform 1 0 15456 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_183
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1644511149
transform 1 0 20240 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_228
timestamp 1644511149
transform 1 0 22080 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_240
timestamp 1644511149
transform 1 0 23184 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_252
timestamp 1644511149
transform 1 0 24288 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_262
timestamp 1644511149
transform 1 0 25208 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_270
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_303
timestamp 1644511149
transform 1 0 28980 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_311
timestamp 1644511149
transform 1 0 29716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_318
timestamp 1644511149
transform 1 0 30360 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_330
timestamp 1644511149
transform 1 0 31464 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_345
timestamp 1644511149
transform 1 0 32844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_369
timestamp 1644511149
transform 1 0 35052 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_381
timestamp 1644511149
transform 1 0 36156 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1644511149
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_483
timestamp 1644511149
transform 1 0 45540 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1644511149
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_92
timestamp 1644511149
transform 1 0 9568 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_101
timestamp 1644511149
transform 1 0 10396 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_105
timestamp 1644511149
transform 1 0 10764 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_134
timestamp 1644511149
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_149
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_157
timestamp 1644511149
transform 1 0 15548 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_179
timestamp 1644511149
transform 1 0 17572 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_200
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_212
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_219
timestamp 1644511149
transform 1 0 21252 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_227
timestamp 1644511149
transform 1 0 21988 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_269
timestamp 1644511149
transform 1 0 25852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_273
timestamp 1644511149
transform 1 0 26220 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_285
timestamp 1644511149
transform 1 0 27324 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_297
timestamp 1644511149
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1644511149
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_315
timestamp 1644511149
transform 1 0 30084 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_336
timestamp 1644511149
transform 1 0 32016 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_348
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_353
timestamp 1644511149
transform 1 0 33580 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_361
timestamp 1644511149
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_466
timestamp 1644511149
transform 1 0 43976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1644511149
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp 1644511149
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_121
timestamp 1644511149
transform 1 0 12236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_129
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1644511149
transform 1 0 13524 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_147
timestamp 1644511149
transform 1 0 14628 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_153
timestamp 1644511149
transform 1 0 15180 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_157
timestamp 1644511149
transform 1 0 15548 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_190
timestamp 1644511149
transform 1 0 18584 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_202
timestamp 1644511149
transform 1 0 19688 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_210
timestamp 1644511149
transform 1 0 20424 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1644511149
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_234
timestamp 1644511149
transform 1 0 22632 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_242
timestamp 1644511149
transform 1 0 23368 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_260
timestamp 1644511149
transform 1 0 25024 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_268
timestamp 1644511149
transform 1 0 25760 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1644511149
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_290
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_297
timestamp 1644511149
transform 1 0 28428 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_309
timestamp 1644511149
transform 1 0 29532 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_318
timestamp 1644511149
transform 1 0 30360 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_326
timestamp 1644511149
transform 1 0 31096 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1644511149
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_492
timestamp 1644511149
transform 1 0 46368 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_496
timestamp 1644511149
transform 1 0 46736 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1644511149
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1644511149
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_101
timestamp 1644511149
transform 1 0 10396 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_106
timestamp 1644511149
transform 1 0 10856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_114
timestamp 1644511149
transform 1 0 11592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_145
timestamp 1644511149
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_152
timestamp 1644511149
transform 1 0 15088 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_164
timestamp 1644511149
transform 1 0 16192 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1644511149
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_201
timestamp 1644511149
transform 1 0 19596 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_234
timestamp 1644511149
transform 1 0 22632 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_242
timestamp 1644511149
transform 1 0 23368 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_276
timestamp 1644511149
transform 1 0 26496 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_313
timestamp 1644511149
transform 1 0 29900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_319
timestamp 1644511149
transform 1 0 30452 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_327
timestamp 1644511149
transform 1 0 31188 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_339
timestamp 1644511149
transform 1 0 32292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_351
timestamp 1644511149
transform 1 0 33396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_440
timestamp 1644511149
transform 1 0 41584 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_452
timestamp 1644511149
transform 1 0 42688 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_464
timestamp 1644511149
transform 1 0 43792 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_468
timestamp 1644511149
transform 1 0 44160 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_481
timestamp 1644511149
transform 1 0 45356 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_487
timestamp 1644511149
transform 1 0 45908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_95
timestamp 1644511149
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_104
timestamp 1644511149
transform 1 0 10672 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_120
timestamp 1644511149
transform 1 0 12144 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_128
timestamp 1644511149
transform 1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_136
timestamp 1644511149
transform 1 0 13616 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_140
timestamp 1644511149
transform 1 0 13984 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_162
timestamp 1644511149
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_173
timestamp 1644511149
transform 1 0 17020 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_183
timestamp 1644511149
transform 1 0 17940 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_196
timestamp 1644511149
transform 1 0 19136 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_209
timestamp 1644511149
transform 1 0 20332 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_229
timestamp 1644511149
transform 1 0 22172 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_234
timestamp 1644511149
transform 1 0 22632 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_243
timestamp 1644511149
transform 1 0 23460 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_254
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_263
timestamp 1644511149
transform 1 0 25300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_271
timestamp 1644511149
transform 1 0 26036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_300
timestamp 1644511149
transform 1 0 28704 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_311
timestamp 1644511149
transform 1 0 29716 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_325
timestamp 1644511149
transform 1 0 31004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1644511149
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_340
timestamp 1644511149
transform 1 0 32384 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_353
timestamp 1644511149
transform 1 0 33580 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_375
timestamp 1644511149
transform 1 0 35604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_387
timestamp 1644511149
transform 1 0 36708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_426
timestamp 1644511149
transform 1 0 40296 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1644511149
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_455
timestamp 1644511149
transform 1 0 42964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_467
timestamp 1644511149
transform 1 0 44068 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_475
timestamp 1644511149
transform 1 0 44804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_480
timestamp 1644511149
transform 1 0 45264 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_499
timestamp 1644511149
transform 1 0 47012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_508
timestamp 1644511149
transform 1 0 47840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_94
timestamp 1644511149
transform 1 0 9752 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_103
timestamp 1644511149
transform 1 0 10580 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_111
timestamp 1644511149
transform 1 0 11316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_116
timestamp 1644511149
transform 1 0 11776 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_128
timestamp 1644511149
transform 1 0 12880 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1644511149
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_149
timestamp 1644511149
transform 1 0 14812 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_160
timestamp 1644511149
transform 1 0 15824 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_172
timestamp 1644511149
transform 1 0 16928 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_188
timestamp 1644511149
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_218
timestamp 1644511149
transform 1 0 21160 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_226
timestamp 1644511149
transform 1 0 21896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_329
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_353
timestamp 1644511149
transform 1 0 33580 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1644511149
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_443
timestamp 1644511149
transform 1 0 41860 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_455
timestamp 1644511149
transform 1 0 42964 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_467
timestamp 1644511149
transform 1 0 44068 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_483
timestamp 1644511149
transform 1 0 45540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_487
timestamp 1644511149
transform 1 0 45908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_97
timestamp 1644511149
transform 1 0 10028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1644511149
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 1644511149
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_131
timestamp 1644511149
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_136
timestamp 1644511149
transform 1 0 13616 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_148
timestamp 1644511149
transform 1 0 14720 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_173
timestamp 1644511149
transform 1 0 17020 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_185
timestamp 1644511149
transform 1 0 18124 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_194
timestamp 1644511149
transform 1 0 18952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_202
timestamp 1644511149
transform 1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_209
timestamp 1644511149
transform 1 0 20332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1644511149
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_229
timestamp 1644511149
transform 1 0 22172 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1644511149
transform 1 0 23184 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_247
timestamp 1644511149
transform 1 0 23828 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_259
timestamp 1644511149
transform 1 0 24932 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_267
timestamp 1644511149
transform 1 0 25668 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 1644511149
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_302
timestamp 1644511149
transform 1 0 28888 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_314
timestamp 1644511149
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_321
timestamp 1644511149
transform 1 0 30636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_359
timestamp 1644511149
transform 1 0 34132 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_371
timestamp 1644511149
transform 1 0 35236 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_383
timestamp 1644511149
transform 1 0 36340 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_469
timestamp 1644511149
transform 1 0 44252 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_481
timestamp 1644511149
transform 1 0 45356 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_498
timestamp 1644511149
transform 1 0 46920 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_89
timestamp 1644511149
transform 1 0 9292 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_96
timestamp 1644511149
transform 1 0 9936 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_104
timestamp 1644511149
transform 1 0 10672 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_129
timestamp 1644511149
transform 1 0 12972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_145
timestamp 1644511149
transform 1 0 14444 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_161
timestamp 1644511149
transform 1 0 15916 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_171
timestamp 1644511149
transform 1 0 16836 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_179
timestamp 1644511149
transform 1 0 17572 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_183
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_200
timestamp 1644511149
transform 1 0 19504 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_208
timestamp 1644511149
transform 1 0 20240 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_212
timestamp 1644511149
transform 1 0 20608 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_224
timestamp 1644511149
transform 1 0 21712 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_236
timestamp 1644511149
transform 1 0 22816 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_257
timestamp 1644511149
transform 1 0 24748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_281
timestamp 1644511149
transform 1 0 26956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_293
timestamp 1644511149
transform 1 0 28060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1644511149
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_312
timestamp 1644511149
transform 1 0 29808 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_324
timestamp 1644511149
transform 1 0 30912 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_336
timestamp 1644511149
transform 1 0 32016 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_348
timestamp 1644511149
transform 1 0 33120 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_485
timestamp 1644511149
transform 1 0 45724 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_507
timestamp 1644511149
transform 1 0 47748 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_515
timestamp 1644511149
transform 1 0 48484 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_97
timestamp 1644511149
transform 1 0 10028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_104
timestamp 1644511149
transform 1 0 10672 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_116
timestamp 1644511149
transform 1 0 11776 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_124
timestamp 1644511149
transform 1 0 12512 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_147
timestamp 1644511149
transform 1 0 14628 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_155
timestamp 1644511149
transform 1 0 15364 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1644511149
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_189
timestamp 1644511149
transform 1 0 18492 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_197
timestamp 1644511149
transform 1 0 19228 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_263
timestamp 1644511149
transform 1 0 25300 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_271
timestamp 1644511149
transform 1 0 26036 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_275
timestamp 1644511149
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_289
timestamp 1644511149
transform 1 0 27692 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_295
timestamp 1644511149
transform 1 0 28244 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_328
timestamp 1644511149
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_343
timestamp 1644511149
transform 1 0 32660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_355
timestamp 1644511149
transform 1 0 33764 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_367
timestamp 1644511149
transform 1 0 34868 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_379
timestamp 1644511149
transform 1 0 35972 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_9
timestamp 1644511149
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1644511149
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_115
timestamp 1644511149
transform 1 0 11684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1644511149
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1644511149
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_163
timestamp 1644511149
transform 1 0 16100 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_171
timestamp 1644511149
transform 1 0 16836 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_181
timestamp 1644511149
transform 1 0 17756 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_217
timestamp 1644511149
transform 1 0 21068 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_228
timestamp 1644511149
transform 1 0 22080 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_236
timestamp 1644511149
transform 1 0 22816 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_267
timestamp 1644511149
transform 1 0 25668 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_279
timestamp 1644511149
transform 1 0 26772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_283
timestamp 1644511149
transform 1 0 27140 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_331
timestamp 1644511149
transform 1 0 31556 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_347
timestamp 1644511149
transform 1 0 33028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_359
timestamp 1644511149
transform 1 0 34132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_483
timestamp 1644511149
transform 1 0 45540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_487
timestamp 1644511149
transform 1 0 45908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_102
timestamp 1644511149
transform 1 0 10488 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1644511149
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_128
timestamp 1644511149
transform 1 0 12880 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_140
timestamp 1644511149
transform 1 0 13984 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_152
timestamp 1644511149
transform 1 0 15088 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_160
timestamp 1644511149
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_176
timestamp 1644511149
transform 1 0 17296 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_184
timestamp 1644511149
transform 1 0 18032 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_208
timestamp 1644511149
transform 1 0 20240 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_233
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_245
timestamp 1644511149
transform 1 0 23644 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_257
timestamp 1644511149
transform 1 0 24748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_269
timestamp 1644511149
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1644511149
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_286
timestamp 1644511149
transform 1 0 27416 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_301
timestamp 1644511149
transform 1 0 28796 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_313
timestamp 1644511149
transform 1 0 29900 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_321
timestamp 1644511149
transform 1 0 30636 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_358
timestamp 1644511149
transform 1 0 34040 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_370
timestamp 1644511149
transform 1 0 35144 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_382
timestamp 1644511149
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1644511149
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_493
timestamp 1644511149
transform 1 0 46460 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_100
timestamp 1644511149
transform 1 0 10304 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_112
timestamp 1644511149
transform 1 0 11408 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_144
timestamp 1644511149
transform 1 0 14352 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_152
timestamp 1644511149
transform 1 0 15088 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_159
timestamp 1644511149
transform 1 0 15732 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_183
timestamp 1644511149
transform 1 0 17940 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_190
timestamp 1644511149
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_201
timestamp 1644511149
transform 1 0 19596 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_205
timestamp 1644511149
transform 1 0 19964 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_220
timestamp 1644511149
transform 1 0 21344 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_229
timestamp 1644511149
transform 1 0 22172 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_241
timestamp 1644511149
transform 1 0 23276 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1644511149
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_260
timestamp 1644511149
transform 1 0 25024 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_266
timestamp 1644511149
transform 1 0 25576 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_274
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_282
timestamp 1644511149
transform 1 0 27048 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_291
timestamp 1644511149
transform 1 0 27876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_300
timestamp 1644511149
transform 1 0 28704 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_327
timestamp 1644511149
transform 1 0 31188 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_331
timestamp 1644511149
transform 1 0 31556 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_344
timestamp 1644511149
transform 1 0 32752 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1644511149
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_512
timestamp 1644511149
transform 1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_131
timestamp 1644511149
transform 1 0 13156 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_138
timestamp 1644511149
transform 1 0 13800 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_158
timestamp 1644511149
transform 1 0 15640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1644511149
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_172
timestamp 1644511149
transform 1 0 16928 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1644511149
transform 1 0 18032 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1644511149
transform 1 0 19136 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1644511149
transform 1 0 20240 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_235
timestamp 1644511149
transform 1 0 22724 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_247
timestamp 1644511149
transform 1 0 23828 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_260
timestamp 1644511149
transform 1 0 25024 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_268
timestamp 1644511149
transform 1 0 25760 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_287
timestamp 1644511149
transform 1 0 27508 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_295
timestamp 1644511149
transform 1 0 28244 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_307
timestamp 1644511149
transform 1 0 29348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_311
timestamp 1644511149
transform 1 0 29716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_340
timestamp 1644511149
transform 1 0 32384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_352
timestamp 1644511149
transform 1 0 33488 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_364
timestamp 1644511149
transform 1 0 34592 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_376
timestamp 1644511149
transform 1 0 35696 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1644511149
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_92
timestamp 1644511149
transform 1 0 9568 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_104
timestamp 1644511149
transform 1 0 10672 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_125
timestamp 1644511149
transform 1 0 12604 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_148
timestamp 1644511149
transform 1 0 14720 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_156
timestamp 1644511149
transform 1 0 15456 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_162
timestamp 1644511149
transform 1 0 16008 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_170
timestamp 1644511149
transform 1 0 16744 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_175
timestamp 1644511149
transform 1 0 17204 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1644511149
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_241
timestamp 1644511149
transform 1 0 23276 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_258
timestamp 1644511149
transform 1 0 24840 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_270
timestamp 1644511149
transform 1 0 25944 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_282
timestamp 1644511149
transform 1 0 27048 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_294
timestamp 1644511149
transform 1 0 28152 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_318
timestamp 1644511149
transform 1 0 30360 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_325
timestamp 1644511149
transform 1 0 31004 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_337
timestamp 1644511149
transform 1 0 32108 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_349
timestamp 1644511149
transform 1 0 33212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1644511149
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_99
timestamp 1644511149
transform 1 0 10212 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_103
timestamp 1644511149
transform 1 0 10580 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1644511149
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_134
timestamp 1644511149
transform 1 0 13432 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_141
timestamp 1644511149
transform 1 0 14076 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_150
timestamp 1644511149
transform 1 0 14904 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_158
timestamp 1644511149
transform 1 0 15640 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_190
timestamp 1644511149
transform 1 0 18584 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_197
timestamp 1644511149
transform 1 0 19228 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_203
timestamp 1644511149
transform 1 0 19780 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_207
timestamp 1644511149
transform 1 0 20148 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_213
timestamp 1644511149
transform 1 0 20700 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 1644511149
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_233
timestamp 1644511149
transform 1 0 22540 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_238
timestamp 1644511149
transform 1 0 23000 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_246
timestamp 1644511149
transform 1 0 23736 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_252
timestamp 1644511149
transform 1 0 24288 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1644511149
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_288
timestamp 1644511149
transform 1 0 27600 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_296
timestamp 1644511149
transform 1 0 28336 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_340
timestamp 1644511149
transform 1 0 32384 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_352
timestamp 1644511149
transform 1 0 33488 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_364
timestamp 1644511149
transform 1 0 34592 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_376
timestamp 1644511149
transform 1 0 35696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1644511149
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_500
timestamp 1644511149
transform 1 0 47104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_110
timestamp 1644511149
transform 1 0 11224 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_118
timestamp 1644511149
transform 1 0 11960 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_122
timestamp 1644511149
transform 1 0 12328 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_128
timestamp 1644511149
transform 1 0 12880 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_162
timestamp 1644511149
transform 1 0 16008 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_170
timestamp 1644511149
transform 1 0 16744 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_217
timestamp 1644511149
transform 1 0 21068 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_228
timestamp 1644511149
transform 1 0 22080 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_237
timestamp 1644511149
transform 1 0 22908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1644511149
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_282
timestamp 1644511149
transform 1 0 27048 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_290
timestamp 1644511149
transform 1 0 27784 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_300
timestamp 1644511149
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_313
timestamp 1644511149
transform 1 0 29900 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_319
timestamp 1644511149
transform 1 0 30452 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_340
timestamp 1644511149
transform 1 0 32384 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_352
timestamp 1644511149
transform 1 0 33488 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_512
timestamp 1644511149
transform 1 0 48208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_129
timestamp 1644511149
transform 1 0 12972 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_133
timestamp 1644511149
transform 1 0 13340 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_140
timestamp 1644511149
transform 1 0 13984 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_152
timestamp 1644511149
transform 1 0 15088 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_190
timestamp 1644511149
transform 1 0 18584 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_202
timestamp 1644511149
transform 1 0 19688 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_206
timestamp 1644511149
transform 1 0 20056 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_216
timestamp 1644511149
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_229
timestamp 1644511149
transform 1 0 22172 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_235
timestamp 1644511149
transform 1 0 22724 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_244
timestamp 1644511149
transform 1 0 23552 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_252
timestamp 1644511149
transform 1 0 24288 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_257
timestamp 1644511149
transform 1 0 24748 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_265
timestamp 1644511149
transform 1 0 25484 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_271
timestamp 1644511149
transform 1 0 26036 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_287
timestamp 1644511149
transform 1 0 27508 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_297
timestamp 1644511149
transform 1 0 28428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_314
timestamp 1644511149
transform 1 0 29992 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_321
timestamp 1644511149
transform 1 0 30636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_333
timestamp 1644511149
transform 1 0 31740 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_340
timestamp 1644511149
transform 1 0 32384 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_352
timestamp 1644511149
transform 1 0 33488 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_364
timestamp 1644511149
transform 1 0 34592 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_376
timestamp 1644511149
transform 1 0 35696 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1644511149
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_145
timestamp 1644511149
transform 1 0 14444 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_149
timestamp 1644511149
transform 1 0 14812 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_161
timestamp 1644511149
transform 1 0 15916 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_173
timestamp 1644511149
transform 1 0 17020 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_181
timestamp 1644511149
transform 1 0 17756 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_190
timestamp 1644511149
transform 1 0 18584 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_216
timestamp 1644511149
transform 1 0 20976 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_235
timestamp 1644511149
transform 1 0 22724 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1644511149
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_273
timestamp 1644511149
transform 1 0 26220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_281
timestamp 1644511149
transform 1 0 26956 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_287
timestamp 1644511149
transform 1 0 27508 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_291
timestamp 1644511149
transform 1 0 27876 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_300
timestamp 1644511149
transform 1 0 28704 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_313
timestamp 1644511149
transform 1 0 29900 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_339
timestamp 1644511149
transform 1 0 32292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_351
timestamp 1644511149
transform 1 0 33396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_133
timestamp 1644511149
transform 1 0 13340 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_139
timestamp 1644511149
transform 1 0 13892 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_190
timestamp 1644511149
transform 1 0 18584 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_202
timestamp 1644511149
transform 1 0 19688 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1644511149
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1644511149
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_230
timestamp 1644511149
transform 1 0 22264 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_240
timestamp 1644511149
transform 1 0 23184 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_252
timestamp 1644511149
transform 1 0 24288 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_258
timestamp 1644511149
transform 1 0 24840 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_264
timestamp 1644511149
transform 1 0 25392 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_269
timestamp 1644511149
transform 1 0 25852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1644511149
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_286
timestamp 1644511149
transform 1 0 27416 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_294
timestamp 1644511149
transform 1 0 28152 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_301
timestamp 1644511149
transform 1 0 28796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_310
timestamp 1644511149
transform 1 0 29624 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_319
timestamp 1644511149
transform 1 0 30452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_331
timestamp 1644511149
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_343
timestamp 1644511149
transform 1 0 32660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_355
timestamp 1644511149
transform 1 0 33764 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1644511149
transform 1 0 34868 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1644511149
transform 1 0 35972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_162
timestamp 1644511149
transform 1 0 16008 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_174
timestamp 1644511149
transform 1 0 17112 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_187
timestamp 1644511149
transform 1 0 18308 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_217
timestamp 1644511149
transform 1 0 21068 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_224
timestamp 1644511149
transform 1 0 21712 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_256
timestamp 1644511149
transform 1 0 24656 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_262
timestamp 1644511149
transform 1 0 25208 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_267
timestamp 1644511149
transform 1 0 25668 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_278
timestamp 1644511149
transform 1 0 26680 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_286
timestamp 1644511149
transform 1 0 27416 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_293
timestamp 1644511149
transform 1 0 28060 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_299
timestamp 1644511149
transform 1 0 28612 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_318
timestamp 1644511149
transform 1 0 30360 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_329
timestamp 1644511149
transform 1 0 31372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_354
timestamp 1644511149
transform 1 0 33672 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1644511149
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_11
timestamp 1644511149
transform 1 0 2116 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_189
timestamp 1644511149
transform 1 0 18492 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_199
timestamp 1644511149
transform 1 0 19412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_211
timestamp 1644511149
transform 1 0 20516 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_215
timestamp 1644511149
transform 1 0 20884 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_236
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_246
timestamp 1644511149
transform 1 0 23736 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_258
timestamp 1644511149
transform 1 0 24840 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_262
timestamp 1644511149
transform 1 0 25208 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_287
timestamp 1644511149
transform 1 0 27508 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_298
timestamp 1644511149
transform 1 0 28520 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_306
timestamp 1644511149
transform 1 0 29256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_311
timestamp 1644511149
transform 1 0 29716 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_322
timestamp 1644511149
transform 1 0 30728 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1644511149
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_343
timestamp 1644511149
transform 1 0 32660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_355
timestamp 1644511149
transform 1 0 33764 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1644511149
transform 1 0 34868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1644511149
transform 1 0 35972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_178
timestamp 1644511149
transform 1 0 17480 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_186
timestamp 1644511149
transform 1 0 18216 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1644511149
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_204
timestamp 1644511149
transform 1 0 19872 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_210
timestamp 1644511149
transform 1 0 20424 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_231
timestamp 1644511149
transform 1 0 22356 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_241
timestamp 1644511149
transform 1 0 23276 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 1644511149
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_261
timestamp 1644511149
transform 1 0 25116 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_282
timestamp 1644511149
transform 1 0 27048 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_290
timestamp 1644511149
transform 1 0 27784 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_298
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1644511149
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_317
timestamp 1644511149
transform 1 0 30268 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_328
timestamp 1644511149
transform 1 0 31280 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_340
timestamp 1644511149
transform 1 0 32384 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_352
timestamp 1644511149
transform 1 0 33488 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_32
timestamp 1644511149
transform 1 0 4048 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_44
timestamp 1644511149
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_189
timestamp 1644511149
transform 1 0 18492 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_201
timestamp 1644511149
transform 1 0 19596 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_209
timestamp 1644511149
transform 1 0 20332 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_233
timestamp 1644511149
transform 1 0 22540 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_243
timestamp 1644511149
transform 1 0 23460 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_250
timestamp 1644511149
transform 1 0 24104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_254
timestamp 1644511149
transform 1 0 24472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_262
timestamp 1644511149
transform 1 0 25208 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_284
timestamp 1644511149
transform 1 0 27232 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_294
timestamp 1644511149
transform 1 0 28152 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_306
timestamp 1644511149
transform 1 0 29256 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_318
timestamp 1644511149
transform 1 0 30360 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_324
timestamp 1644511149
transform 1 0 30912 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_508
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1644511149
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_169
timestamp 1644511149
transform 1 0 16652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_173
timestamp 1644511149
transform 1 0 17020 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_180
timestamp 1644511149
transform 1 0 17664 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_188
timestamp 1644511149
transform 1 0 18400 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_200
timestamp 1644511149
transform 1 0 19504 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_212
timestamp 1644511149
transform 1 0 20608 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_218
timestamp 1644511149
transform 1 0 21160 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_223
timestamp 1644511149
transform 1 0 21620 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_241
timestamp 1644511149
transform 1 0 23276 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1644511149
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_261
timestamp 1644511149
transform 1 0 25116 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_271
timestamp 1644511149
transform 1 0 26036 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_280
timestamp 1644511149
transform 1 0 26864 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_319
timestamp 1644511149
transform 1 0 30452 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_173
timestamp 1644511149
transform 1 0 17020 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_192
timestamp 1644511149
transform 1 0 18768 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_199
timestamp 1644511149
transform 1 0 19412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_211
timestamp 1644511149
transform 1 0 20516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_232
timestamp 1644511149
transform 1 0 22448 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_256
timestamp 1644511149
transform 1 0 24656 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_266
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1644511149
transform 1 0 26404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_286
timestamp 1644511149
transform 1 0 27416 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_294
timestamp 1644511149
transform 1 0 28152 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_300
timestamp 1644511149
transform 1 0 28704 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_307
timestamp 1644511149
transform 1 0 29348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_319
timestamp 1644511149
transform 1 0 30452 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_340
timestamp 1644511149
transform 1 0 32384 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_352
timestamp 1644511149
transform 1 0 33488 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_364
timestamp 1644511149
transform 1 0 34592 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_376
timestamp 1644511149
transform 1 0 35696 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1644511149
transform 1 0 36800 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_512
timestamp 1644511149
transform 1 0 48208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_157
timestamp 1644511149
transform 1 0 15548 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_178
timestamp 1644511149
transform 1 0 17480 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_182
timestamp 1644511149
transform 1 0 17848 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_202
timestamp 1644511149
transform 1 0 19688 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_214
timestamp 1644511149
transform 1 0 20792 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_226
timestamp 1644511149
transform 1 0 21896 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_234
timestamp 1644511149
transform 1 0 22632 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_242
timestamp 1644511149
transform 1 0 23368 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_261
timestamp 1644511149
transform 1 0 25116 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_269
timestamp 1644511149
transform 1 0 25852 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_274
timestamp 1644511149
transform 1 0 26312 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_282
timestamp 1644511149
transform 1 0 27048 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_288
timestamp 1644511149
transform 1 0 27600 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_295
timestamp 1644511149
transform 1 0 28244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_316
timestamp 1644511149
transform 1 0 30176 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_324
timestamp 1644511149
transform 1 0 30912 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_331
timestamp 1644511149
transform 1 0 31556 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_338
timestamp 1644511149
transform 1 0 32200 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_350
timestamp 1644511149
transform 1 0 33304 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1644511149
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_497
timestamp 1644511149
transform 1 0 46828 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_178
timestamp 1644511149
transform 1 0 17480 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_184
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_191
timestamp 1644511149
transform 1 0 18676 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_201
timestamp 1644511149
transform 1 0 19596 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_212
timestamp 1644511149
transform 1 0 20608 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_216
timestamp 1644511149
transform 1 0 20976 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1644511149
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_241
timestamp 1644511149
transform 1 0 23276 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_253
timestamp 1644511149
transform 1 0 24380 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_265
timestamp 1644511149
transform 1 0 25484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_269
timestamp 1644511149
transform 1 0 25852 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_275
timestamp 1644511149
transform 1 0 26404 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_287
timestamp 1644511149
transform 1 0 27508 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_295
timestamp 1644511149
transform 1 0 28244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_302
timestamp 1644511149
transform 1 0 28888 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_310
timestamp 1644511149
transform 1 0 29624 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1644511149
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_512
timestamp 1644511149
transform 1 0 48208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_173
timestamp 1644511149
transform 1 0 17020 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_182
timestamp 1644511149
transform 1 0 17848 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_204
timestamp 1644511149
transform 1 0 19872 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_212
timestamp 1644511149
transform 1 0 20608 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_246
timestamp 1644511149
transform 1 0 23736 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_268
timestamp 1644511149
transform 1 0 25760 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_280
timestamp 1644511149
transform 1 0 26864 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_290
timestamp 1644511149
transform 1 0 27784 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_296
timestamp 1644511149
transform 1 0 28336 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_315
timestamp 1644511149
transform 1 0 30084 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_323
timestamp 1644511149
transform 1 0 30820 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_346
timestamp 1644511149
transform 1 0 32936 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_358
timestamp 1644511149
transform 1 0 34040 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_178
timestamp 1644511149
transform 1 0 17480 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_187
timestamp 1644511149
transform 1 0 18308 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_200
timestamp 1644511149
transform 1 0 19504 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_212
timestamp 1644511149
transform 1 0 20608 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_229
timestamp 1644511149
transform 1 0 22172 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_241
timestamp 1644511149
transform 1 0 23276 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_262
timestamp 1644511149
transform 1 0 25208 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_274
timestamp 1644511149
transform 1 0 26312 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_284
timestamp 1644511149
transform 1 0 27232 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_288
timestamp 1644511149
transform 1 0 27600 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_296
timestamp 1644511149
transform 1 0 28336 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_309
timestamp 1644511149
transform 1 0 29532 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_318
timestamp 1644511149
transform 1 0 30360 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_340
timestamp 1644511149
transform 1 0 32384 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_352
timestamp 1644511149
transform 1 0 33488 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_364
timestamp 1644511149
transform 1 0 34592 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_376
timestamp 1644511149
transform 1 0 35696 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1644511149
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1644511149
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1644511149
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_185
timestamp 1644511149
transform 1 0 18124 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_193
timestamp 1644511149
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_229
timestamp 1644511149
transform 1 0 22172 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_235
timestamp 1644511149
transform 1 0 22724 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1644511149
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_261
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_284
timestamp 1644511149
transform 1 0 27232 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_290
timestamp 1644511149
transform 1 0 27784 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_295
timestamp 1644511149
transform 1 0 28244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_315
timestamp 1644511149
transform 1 0 30084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_327
timestamp 1644511149
transform 1 0 31188 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_339
timestamp 1644511149
transform 1 0 32292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_351
timestamp 1644511149
transform 1 0 33396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_28
timestamp 1644511149
transform 1 0 3680 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1644511149
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_177
timestamp 1644511149
transform 1 0 17388 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_183
timestamp 1644511149
transform 1 0 17940 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_195
timestamp 1644511149
transform 1 0 19044 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_207
timestamp 1644511149
transform 1 0 20148 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1644511149
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_229
timestamp 1644511149
transform 1 0 22172 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_234
timestamp 1644511149
transform 1 0 22632 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_244
timestamp 1644511149
transform 1 0 23552 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_255
timestamp 1644511149
transform 1 0 24564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_267
timestamp 1644511149
transform 1 0 25668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_297
timestamp 1644511149
transform 1 0 28428 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_318
timestamp 1644511149
transform 1 0 30360 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_325
timestamp 1644511149
transform 1 0 31004 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_333
timestamp 1644511149
transform 1 0 31740 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1644511149
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_212
timestamp 1644511149
transform 1 0 20608 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_230
timestamp 1644511149
transform 1 0 22264 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_239
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_293
timestamp 1644511149
transform 1 0 28060 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_303
timestamp 1644511149
transform 1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_312
timestamp 1644511149
transform 1 0 29808 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_324
timestamp 1644511149
transform 1 0 30912 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_336
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_348
timestamp 1644511149
transform 1 0 33120 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1644511149
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_483
timestamp 1644511149
transform 1 0 45540 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_487
timestamp 1644511149
transform 1 0 45908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_512
timestamp 1644511149
transform 1 0 48208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_191
timestamp 1644511149
transform 1 0 18676 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_199
timestamp 1644511149
transform 1 0 19412 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_229
timestamp 1644511149
transform 1 0 22172 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_240
timestamp 1644511149
transform 1 0 23184 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_248
timestamp 1644511149
transform 1 0 23920 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_256
timestamp 1644511149
transform 1 0 24656 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_260
timestamp 1644511149
transform 1 0 25024 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_264
timestamp 1644511149
transform 1 0 25392 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_268
timestamp 1644511149
transform 1 0 25760 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1644511149
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_285
timestamp 1644511149
transform 1 0 27324 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_314
timestamp 1644511149
transform 1 0 29992 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_326
timestamp 1644511149
transform 1 0 31096 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 1644511149
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_481
timestamp 1644511149
transform 1 0 45356 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_490
timestamp 1644511149
transform 1 0 46184 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_494
timestamp 1644511149
transform 1 0 46552 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_498
timestamp 1644511149
transform 1 0 46920 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_180
timestamp 1644511149
transform 1 0 17664 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_184
timestamp 1644511149
transform 1 0 18032 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_190
timestamp 1644511149
transform 1 0 18584 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_206
timestamp 1644511149
transform 1 0 20056 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_210
timestamp 1644511149
transform 1 0 20424 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_214
timestamp 1644511149
transform 1 0 20792 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_222
timestamp 1644511149
transform 1 0 21528 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_228
timestamp 1644511149
transform 1 0 22080 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_275
timestamp 1644511149
transform 1 0 26404 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_279
timestamp 1644511149
transform 1 0 26772 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_290
timestamp 1644511149
transform 1 0 27784 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_302
timestamp 1644511149
transform 1 0 28888 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_472
timestamp 1644511149
transform 1 0 44528 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_483
timestamp 1644511149
transform 1 0 45540 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_509
timestamp 1644511149
transform 1 0 47932 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_515
timestamp 1644511149
transform 1 0 48484 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_187
timestamp 1644511149
transform 1 0 18308 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_200
timestamp 1644511149
transform 1 0 19504 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_212
timestamp 1644511149
transform 1 0 20608 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_245
timestamp 1644511149
transform 1 0 23644 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_257
timestamp 1644511149
transform 1 0 24748 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_265
timestamp 1644511149
transform 1 0 25484 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_269
timestamp 1644511149
transform 1 0 25852 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_277
timestamp 1644511149
transform 1 0 26588 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_321
timestamp 1644511149
transform 1 0 30636 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_333
timestamp 1644511149
transform 1 0 31740 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_481
timestamp 1644511149
transform 1 0 45356 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_487
timestamp 1644511149
transform 1 0 45908 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_500
timestamp 1644511149
transform 1 0 47104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_508
timestamp 1644511149
transform 1 0 47840 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_179
timestamp 1644511149
transform 1 0 17572 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_192
timestamp 1644511149
transform 1 0 18768 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_238
timestamp 1644511149
transform 1 0 23000 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1644511149
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_196
timestamp 1644511149
transform 1 0 19136 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_208
timestamp 1644511149
transform 1 0 20240 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1644511149
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_457
timestamp 1644511149
transform 1 0 43148 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_471
timestamp 1644511149
transform 1 0 44436 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1644511149
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_512
timestamp 1644511149
transform 1 0 48208 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_9
timestamp 1644511149
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_13
timestamp 1644511149
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_25
timestamp 1644511149
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_37
timestamp 1644511149
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1644511149
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_489
timestamp 1644511149
transform 1 0 46092 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_500
timestamp 1644511149
transform 1 0 47104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_508
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_302
timestamp 1644511149
transform 1 0 28888 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_314
timestamp 1644511149
transform 1 0 29992 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_326
timestamp 1644511149
transform 1 0 31096 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 1644511149
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1644511149
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_7
timestamp 1644511149
transform 1 0 1748 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_19
timestamp 1644511149
transform 1 0 2852 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_31
timestamp 1644511149
transform 1 0 3956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_43
timestamp 1644511149
transform 1 0 5060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_276
timestamp 1644511149
transform 1 0 26496 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_302
timestamp 1644511149
transform 1 0 28888 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_314
timestamp 1644511149
transform 1 0 29992 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_326
timestamp 1644511149
transform 1 0 31096 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_334
timestamp 1644511149
transform 1 0 31832 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_492
timestamp 1644511149
transform 1 0 46368 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_499
timestamp 1644511149
transform 1 0 47012 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1644511149
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_304
timestamp 1644511149
transform 1 0 29072 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_312
timestamp 1644511149
transform 1 0 29808 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_324
timestamp 1644511149
transform 1 0 30912 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_336
timestamp 1644511149
transform 1 0 32016 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_348
timestamp 1644511149
transform 1 0 33120 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_360
timestamp 1644511149
transform 1 0 34224 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_412
timestamp 1644511149
transform 1 0 39008 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_289
timestamp 1644511149
transform 1 0 27692 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_312
timestamp 1644511149
transform 1 0 29808 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_324
timestamp 1644511149
transform 1 0 30912 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_455
timestamp 1644511149
transform 1 0 42964 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_463
timestamp 1644511149
transform 1 0 43700 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_467
timestamp 1644511149
transform 1 0 44068 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_479
timestamp 1644511149
transform 1 0 45172 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_483
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_490
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1644511149
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_293
timestamp 1644511149
transform 1 0 28060 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_297
timestamp 1644511149
transform 1 0 28428 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_305
timestamp 1644511149
transform 1 0 29164 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_441
timestamp 1644511149
transform 1 0 41676 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_78_447
timestamp 1644511149
transform 1 0 42228 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_455
timestamp 1644511149
transform 1 0 42964 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_459
timestamp 1644511149
transform 1 0 43332 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_466
timestamp 1644511149
transform 1 0 43976 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_474
timestamp 1644511149
transform 1 0 44712 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_11
timestamp 1644511149
transform 1 0 2116 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_45
timestamp 1644511149
transform 1 0 5244 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_53
timestamp 1644511149
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_101
timestamp 1644511149
transform 1 0 10396 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_266
timestamp 1644511149
transform 1 0 25576 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1644511149
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_284
timestamp 1644511149
transform 1 0 27232 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_296
timestamp 1644511149
transform 1 0 28336 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_308
timestamp 1644511149
transform 1 0 29440 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_320
timestamp 1644511149
transform 1 0 30544 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_332
timestamp 1644511149
transform 1 0 31648 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_340
timestamp 1644511149
transform 1 0 32384 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_352
timestamp 1644511149
transform 1 0 33488 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_364
timestamp 1644511149
transform 1 0 34592 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_376
timestamp 1644511149
transform 1 0 35696 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1644511149
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_440
timestamp 1644511149
transform 1 0 41584 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_473
timestamp 1644511149
transform 1 0 44620 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_481
timestamp 1644511149
transform 1 0 45356 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_489
timestamp 1644511149
transform 1 0 46092 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1644511149
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_508
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1644511149
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_54
timestamp 1644511149
transform 1 0 6072 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_66
timestamp 1644511149
transform 1 0 7176 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_78
timestamp 1644511149
transform 1 0 8280 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_122
timestamp 1644511149
transform 1 0 12328 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_130
timestamp 1644511149
transform 1 0 13064 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1644511149
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_188
timestamp 1644511149
transform 1 0 18400 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_202
timestamp 1644511149
transform 1 0 19688 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_227
timestamp 1644511149
transform 1 0 21988 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_239
timestamp 1644511149
transform 1 0 23092 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_261
timestamp 1644511149
transform 1 0 25116 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_285
timestamp 1644511149
transform 1 0 27324 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_297
timestamp 1644511149
transform 1 0 28428 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_305
timestamp 1644511149
transform 1 0 29164 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_329
timestamp 1644511149
transform 1 0 31372 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_353
timestamp 1644511149
transform 1 0 33580 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_361
timestamp 1644511149
transform 1 0 34316 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_406
timestamp 1644511149
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1644511149
transform 1 0 39560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_457
timestamp 1644511149
transform 1 0 43148 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_7
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_14
timestamp 1644511149
transform 1 0 2392 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_26
timestamp 1644511149
transform 1 0 3496 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_37
timestamp 1644511149
transform 1 0 4508 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_49
timestamp 1644511149
transform 1 0 5612 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_101
timestamp 1644511149
transform 1 0 10396 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_121
timestamp 1644511149
transform 1 0 12236 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_126
timestamp 1644511149
transform 1 0 12696 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_134
timestamp 1644511149
transform 1 0 13432 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_157
timestamp 1644511149
transform 1 0 15548 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_165
timestamp 1644511149
transform 1 0 16284 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_189
timestamp 1644511149
transform 1 0 18492 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_195
timestamp 1644511149
transform 1 0 19044 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_228
timestamp 1644511149
transform 1 0 22080 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_240
timestamp 1644511149
transform 1 0 23184 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_252
timestamp 1644511149
transform 1 0 24288 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_284
timestamp 1644511149
transform 1 0 27232 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_292
timestamp 1644511149
transform 1 0 27968 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_316
timestamp 1644511149
transform 1 0 30176 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_328
timestamp 1644511149
transform 1 0 31280 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_340
timestamp 1644511149
transform 1 0 32384 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_352
timestamp 1644511149
transform 1 0 33488 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_364
timestamp 1644511149
transform 1 0 34592 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_376
timestamp 1644511149
transform 1 0 35696 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_388
timestamp 1644511149
transform 1 0 36800 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_431
timestamp 1644511149
transform 1 0 40756 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_437
timestamp 1644511149
transform 1 0 41308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1644511149
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_57
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_67
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_75
timestamp 1644511149
transform 1 0 8004 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1644511149
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_149
timestamp 1644511149
transform 1 0 14812 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_161
timestamp 1644511149
transform 1 0 15916 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_191
timestamp 1644511149
transform 1 0 18676 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_201
timestamp 1644511149
transform 1 0 19596 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_216
timestamp 1644511149
transform 1 0 20976 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_268
timestamp 1644511149
transform 1 0 25760 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_300
timestamp 1644511149
transform 1 0 28704 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_332
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_406
timestamp 1644511149
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_418
timestamp 1644511149
transform 1 0 39560 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_441
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_447
timestamp 1644511149
transform 1 0 42228 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_511
timestamp 1644511149
transform 1 0 48116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_515
timestamp 1644511149
transform 1 0 48484 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0571_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0573_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0574_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0575_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28336 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0576_
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0577_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0578_
timestamp 1644511149
transform 1 0 22632 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0579_
timestamp 1644511149
transform 1 0 18216 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0580_
timestamp 1644511149
transform 1 0 19044 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0581_
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0582_
timestamp 1644511149
transform 1 0 26404 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0583_
timestamp 1644511149
transform 1 0 27232 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0584_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0585_
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0586_
timestamp 1644511149
transform 1 0 20792 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0587_
timestamp 1644511149
transform 1 0 21712 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0588_
timestamp 1644511149
transform 1 0 21988 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0589_
timestamp 1644511149
transform 1 0 22908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0590_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23828 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10120 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0594_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0595_
timestamp 1644511149
transform 1 0 12144 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0596_
timestamp 1644511149
transform 1 0 18216 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0597_
timestamp 1644511149
transform 1 0 17020 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0598_
timestamp 1644511149
transform 1 0 17296 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0599_
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0600_
timestamp 1644511149
transform 1 0 15456 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0601_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24840 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0604_
timestamp 1644511149
transform 1 0 30360 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31004 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0607_
timestamp 1644511149
transform 1 0 29992 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0608_
timestamp 1644511149
transform 1 0 29072 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1644511149
transform 1 0 31188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0610_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30820 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0611_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30084 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1644511149
transform 1 0 28152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0613_
timestamp 1644511149
transform 1 0 27140 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1644511149
transform 1 0 26128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0615_
timestamp 1644511149
transform 1 0 23000 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0616_
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0617_
timestamp 1644511149
transform 1 0 24748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0618_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1644511149
transform 1 0 23736 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0620_
timestamp 1644511149
transform 1 0 21988 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0622_
timestamp 1644511149
transform 1 0 22264 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0623_
timestamp 1644511149
transform 1 0 23552 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0625_
timestamp 1644511149
transform 1 0 20700 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1644511149
transform 1 0 17480 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1644511149
transform 1 0 15364 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0628_
timestamp 1644511149
transform 1 0 15548 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0629_
timestamp 1644511149
transform 1 0 15272 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0630_
timestamp 1644511149
transform 1 0 15364 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0631_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1644511149
transform 1 0 17664 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0633_
timestamp 1644511149
transform 1 0 22632 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0634_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0635_
timestamp 1644511149
transform 1 0 15272 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15548 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0638_
timestamp 1644511149
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0640_
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13524 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0643_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12420 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0645_
timestamp 1644511149
transform 1 0 12696 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0646_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1644511149
transform 1 0 13800 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0648_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11776 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 1644511149
transform 1 0 12052 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1644511149
transform 1 0 14628 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0651_
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0652_
timestamp 1644511149
transform 1 0 12972 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0653_
timestamp 1644511149
transform 1 0 11868 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1644511149
transform 1 0 10212 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0655_
timestamp 1644511149
transform 1 0 9660 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0657_
timestamp 1644511149
transform 1 0 14352 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0658_
timestamp 1644511149
transform 1 0 10488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0659_
timestamp 1644511149
transform 1 0 10304 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0660_
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1644511149
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0662_
timestamp 1644511149
transform 1 0 10212 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0663_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9016 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1644511149
transform 1 0 10120 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0665_
timestamp 1644511149
transform 1 0 9476 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0666_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0667_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1644511149
transform 1 0 9936 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0669_
timestamp 1644511149
transform 1 0 8648 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0670_
timestamp 1644511149
transform 1 0 13156 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1644511149
transform 1 0 12512 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0672_
timestamp 1644511149
transform 1 0 15272 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0673_
timestamp 1644511149
transform 1 0 13892 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0674_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11224 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1644511149
transform 1 0 14536 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0676_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0677_
timestamp 1644511149
transform 1 0 12972 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1644511149
transform 1 0 13892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0679_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0680_
timestamp 1644511149
transform 1 0 15088 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1644511149
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0682_
timestamp 1644511149
transform 1 0 12512 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0684_
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0685_
timestamp 1644511149
transform 1 0 17848 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0686_
timestamp 1644511149
transform 1 0 17204 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0687_
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0688_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0689_
timestamp 1644511149
transform 1 0 20792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0691_
timestamp 1644511149
transform 1 0 17204 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0692_
timestamp 1644511149
transform 1 0 17940 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1644511149
transform 1 0 20056 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0694_
timestamp 1644511149
transform 1 0 18032 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0696_
timestamp 1644511149
transform 1 0 18952 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0697_
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0698_
timestamp 1644511149
transform 1 0 17940 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1644511149
transform 1 0 20516 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0700_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0702_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0703_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0704_
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0705_
timestamp 1644511149
transform 1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0707_
timestamp 1644511149
transform 1 0 20700 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0708_
timestamp 1644511149
transform 1 0 20700 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0710_
timestamp 1644511149
transform 1 0 20148 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0711_
timestamp 1644511149
transform 1 0 20976 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0712_
timestamp 1644511149
transform 1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0714_
timestamp 1644511149
transform 1 0 22356 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0715_
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1644511149
transform 1 0 24472 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0718_
timestamp 1644511149
transform 1 0 24104 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0719_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 1644511149
transform 1 0 19688 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0721_
timestamp 1644511149
transform 1 0 27140 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0722_
timestamp 1644511149
transform 1 0 25300 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20976 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0725_
timestamp 1644511149
transform 1 0 22448 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0726_
timestamp 1644511149
transform 1 0 22356 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0727_
timestamp 1644511149
transform 1 0 24748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0728_
timestamp 1644511149
transform 1 0 22080 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0729_
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24564 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0731_
timestamp 1644511149
transform 1 0 22356 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _0732_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0733_
timestamp 1644511149
transform 1 0 25668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0734_
timestamp 1644511149
transform 1 0 23092 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0735_
timestamp 1644511149
transform 1 0 20424 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0736_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0737_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0738_
timestamp 1644511149
transform 1 0 23828 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0739_
timestamp 1644511149
transform 1 0 24472 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0740_
timestamp 1644511149
transform 1 0 17940 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0741_
timestamp 1644511149
transform 1 0 29348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _0742_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _0743_
timestamp 1644511149
transform 1 0 25484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17664 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0745_
timestamp 1644511149
transform 1 0 18032 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0746_
timestamp 1644511149
transform 1 0 21252 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0747_
timestamp 1644511149
transform 1 0 22632 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0748_
timestamp 1644511149
transform 1 0 22080 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0749_
timestamp 1644511149
transform 1 0 23092 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0750_
timestamp 1644511149
transform 1 0 23184 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0751_
timestamp 1644511149
transform 1 0 27416 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0752_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20976 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22080 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0755_
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0756_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _0757_
timestamp 1644511149
transform 1 0 22724 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0758_
timestamp 1644511149
transform 1 0 27876 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0759_
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0760_
timestamp 1644511149
transform 1 0 25944 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0761_
timestamp 1644511149
transform 1 0 24932 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0762_
timestamp 1644511149
transform 1 0 23092 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0763_
timestamp 1644511149
transform 1 0 23092 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0764_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 1644511149
transform 1 0 26036 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0766_
timestamp 1644511149
transform 1 0 25944 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0767_
timestamp 1644511149
transform 1 0 25852 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1644511149
transform 1 0 26956 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0769_
timestamp 1644511149
transform 1 0 25576 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0770_
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0771_
timestamp 1644511149
transform 1 0 25024 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0772_
timestamp 1644511149
transform 1 0 29900 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _0773_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0774_
timestamp 1644511149
transform 1 0 22724 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0775_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0776_
timestamp 1644511149
transform 1 0 27968 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0777_
timestamp 1644511149
transform 1 0 27876 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0778_
timestamp 1644511149
transform 1 0 27232 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0779_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0780_
timestamp 1644511149
transform 1 0 27600 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 1644511149
transform 1 0 28612 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0782_
timestamp 1644511149
transform 1 0 27876 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0783_
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0784_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26128 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0785_
timestamp 1644511149
transform 1 0 29808 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0786_
timestamp 1644511149
transform 1 0 29900 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0787_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27692 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0788_
timestamp 1644511149
transform 1 0 28704 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0789_
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0790_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0791_
timestamp 1644511149
transform 1 0 28428 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0792_
timestamp 1644511149
transform 1 0 28152 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0793_
timestamp 1644511149
transform 1 0 30728 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0794_
timestamp 1644511149
transform 1 0 31004 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0795_
timestamp 1644511149
transform 1 0 31004 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0796_
timestamp 1644511149
transform 1 0 29900 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0797_
timestamp 1644511149
transform 1 0 31924 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0798_
timestamp 1644511149
transform 1 0 30452 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0799_
timestamp 1644511149
transform 1 0 30636 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0800_
timestamp 1644511149
transform 1 0 17848 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0801_
timestamp 1644511149
transform 1 0 26680 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0802_
timestamp 1644511149
transform 1 0 26036 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0803_
timestamp 1644511149
transform 1 0 18124 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0804_
timestamp 1644511149
transform 1 0 18492 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0805_
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0806_
timestamp 1644511149
transform 1 0 18124 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0808_
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0809_
timestamp 1644511149
transform 1 0 17940 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0810_
timestamp 1644511149
transform 1 0 17112 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0811_
timestamp 1644511149
transform 1 0 16928 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0813_
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0814_
timestamp 1644511149
transform 1 0 19136 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0815_
timestamp 1644511149
transform 1 0 17296 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0816_
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0817_
timestamp 1644511149
transform 1 0 18676 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0818_
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0819_
timestamp 1644511149
transform 1 0 22264 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0820_
timestamp 1644511149
transform 1 0 21344 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0821_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0822_
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0823_
timestamp 1644511149
transform 1 0 17848 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0824_
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0825_
timestamp 1644511149
transform 1 0 16836 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0826_
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0827_
timestamp 1644511149
transform 1 0 20700 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0828_
timestamp 1644511149
transform 1 0 19780 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0829_
timestamp 1644511149
transform 1 0 22540 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0830_
timestamp 1644511149
transform 1 0 22816 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 1644511149
transform 1 0 22172 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0832_
timestamp 1644511149
transform 1 0 21804 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1644511149
transform 1 0 30360 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0834_
timestamp 1644511149
transform 1 0 29992 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 1644511149
transform 1 0 27600 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0836_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0837_
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0838_
timestamp 1644511149
transform 1 0 28244 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0839_
timestamp 1644511149
transform 1 0 27048 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0840_
timestamp 1644511149
transform 1 0 27876 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0841_
timestamp 1644511149
transform 1 0 28704 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0842_
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0843_
timestamp 1644511149
transform 1 0 30084 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0844_
timestamp 1644511149
transform 1 0 29808 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0845_
timestamp 1644511149
transform 1 0 30728 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0846_
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0847_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0848_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0849_
timestamp 1644511149
transform 1 0 26496 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0850_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0851_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0852_
timestamp 1644511149
transform 1 0 25852 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0853_
timestamp 1644511149
transform 1 0 25668 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0854_
timestamp 1644511149
transform 1 0 25116 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0855_
timestamp 1644511149
transform 1 0 28244 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0856_
timestamp 1644511149
transform 1 0 27232 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0857_
timestamp 1644511149
transform 1 0 27968 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1644511149
transform 1 0 24196 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0859_
timestamp 1644511149
transform 1 0 23276 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0860_
timestamp 1644511149
transform 1 0 31188 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0861_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31924 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1644511149
transform 1 0 45632 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1644511149
transform 1 0 28152 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1644511149
transform 1 0 46552 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0873_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1644511149
transform 1 0 28612 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1644511149
transform 1 0 43056 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0879_
timestamp 1644511149
transform 1 0 30820 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0885_
timestamp 1644511149
transform 1 0 17572 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0886_
timestamp 1644511149
transform 1 0 16836 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1644511149
transform 1 0 46552 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0892_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  _0893_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform 1 0 16928 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0898_
timestamp 1644511149
transform 1 0 17940 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 11868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0904_
timestamp 1644511149
transform 1 0 16376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 11592 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1644511149
transform 1 0 15732 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 11500 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0910_
timestamp 1644511149
transform 1 0 17112 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 18768 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 7912 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1644511149
transform 1 0 15088 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1644511149
transform 1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0916_
timestamp 1644511149
transform -1 0 18584 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0917_
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 18032 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1644511149
transform 1 0 42780 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1644511149
transform 1 0 41952 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0923_
timestamp 1644511149
transform 1 0 18400 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 25300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0929_
timestamp 1644511149
transform 1 0 17940 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 4968 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 46644 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 43700 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1644511149
transform 1 0 43884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 38732 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0935_
timestamp 1644511149
transform 1 0 17020 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 18676 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 19412 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 10488 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 2208 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 2208 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0941_
timestamp 1644511149
transform 1 0 18308 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 45908 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 15732 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0947_
timestamp 1644511149
transform 1 0 41216 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0948_
timestamp 1644511149
transform 1 0 18032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 15272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 16744 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 14536 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 13616 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 18308 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0954_
timestamp 1644511149
transform 1 0 41400 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 40020 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 32936 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 46736 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 33304 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0960_
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 43700 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0966_
timestamp 1644511149
transform 1 0 18308 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 2024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0972_
timestamp 1644511149
transform 1 0 19504 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 31280 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0979_
timestamp 1644511149
transform 1 0 19872 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0980_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _0982_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1644511149
transform 1 0 45080 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 1644511149
transform 1 0 45632 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0985_
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0986_
timestamp 1644511149
transform 1 0 45448 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0987_
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0988_
timestamp 1644511149
transform 1 0 47380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0989_
timestamp 1644511149
transform 1 0 25944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0990_
timestamp 1644511149
transform 1 0 26036 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0991_
timestamp 1644511149
transform 1 0 25944 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0992_
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _0993_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0994_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0995_
timestamp 1644511149
transform 1 0 44804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0996_
timestamp 1644511149
transform 1 0 47656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _0997_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45908 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0998_
timestamp 1644511149
transform 1 0 46092 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_4  _0999_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45632 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__xnor2_4  _1000_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45908 0 1 38080
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _1001_
timestamp 1644511149
transform 1 0 44988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1002_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1003_
timestamp 1644511149
transform 1 0 45172 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1004_
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1005_
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45908 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1007_
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27416 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1010_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _1011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26864 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1644511149
transform 1 0 26036 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1013_
timestamp 1644511149
transform 1 0 25392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26864 0 1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1016_
timestamp 1644511149
transform 1 0 27784 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1017_
timestamp 1644511149
transform 1 0 27968 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 1644511149
transform 1 0 45632 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1019_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45540 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1020_
timestamp 1644511149
transform 1 0 43240 0 -1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1021_
timestamp 1644511149
transform 1 0 44804 0 -1 40256
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _1022_
timestamp 1644511149
transform 1 0 16836 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 24472 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1644511149
transform 1 0 27968 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1644511149
transform 1 0 26128 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1644511149
transform 1 0 28704 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1644511149
transform 1 0 32384 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1644511149
transform 1 0 30728 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1032_
timestamp 1644511149
transform 1 0 21252 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform 1 0 21896 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1644511149
transform 1 0 20516 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1644511149
transform 1 0 16744 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1038_
timestamp 1644511149
transform 1 0 29900 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1644511149
transform 1 0 17204 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 17664 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1044_
timestamp 1644511149
transform 1 0 23000 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1644511149
transform 1 0 30728 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1644511149
transform 1 0 29072 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1050_
timestamp 1644511149
transform 1 0 22264 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1644511149
transform 1 0 24288 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1644511149
transform 1 0 23828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1644511149
transform 1 0 24564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1056_
timestamp 1644511149
transform 1 0 19320 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1644511149
transform 1 0 18952 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1644511149
transform 1 0 19872 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1061_
timestamp 1644511149
transform 1 0 22080 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1062_
timestamp 1644511149
transform 1 0 22816 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1063_
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1064_
timestamp 1644511149
transform 1 0 19596 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1065_
timestamp 1644511149
transform 1 0 20240 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1066_
timestamp 1644511149
transform 1 0 17204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1067_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1068_
timestamp 1644511149
transform 1 0 18032 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1069_
timestamp 1644511149
transform 1 0 14260 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1070_
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1071_
timestamp 1644511149
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1644511149
transform 1 0 13156 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1073_
timestamp 1644511149
transform 1 0 12144 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1074_
timestamp 1644511149
transform 1 0 10672 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1075_
timestamp 1644511149
transform 1 0 9108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1076_
timestamp 1644511149
transform 1 0 9200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1077_
timestamp 1644511149
transform 1 0 12972 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1078_
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1079_
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1080_
timestamp 1644511149
transform 1 0 9200 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1644511149
transform 1 0 13064 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1082_
timestamp 1644511149
transform 1 0 10672 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1083_
timestamp 1644511149
transform 1 0 13248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1085_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1086_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1087_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1088_
timestamp 1644511149
transform 1 0 16468 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1089_
timestamp 1644511149
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1090_
timestamp 1644511149
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1091_
timestamp 1644511149
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1092_
timestamp 1644511149
transform 1 0 23000 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1093_
timestamp 1644511149
transform 1 0 25668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 25944 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1095_
timestamp 1644511149
transform 1 0 29992 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1096_
timestamp 1644511149
transform 1 0 28336 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1644511149
transform 1 0 30360 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1644511149
transform 1 0 20056 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1100_
timestamp 1644511149
transform 1 0 27232 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1101_
timestamp 1644511149
transform 1 0 25116 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1644511149
transform 1 0 29808 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1644511149
transform 1 0 30452 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 1644511149
transform 1 0 28428 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 1644511149
transform 1 0 30544 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1107_
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1108_
timestamp 1644511149
transform 1 0 19504 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 1644511149
transform 1 0 20700 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 1644511149
transform 1 0 15640 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1114_
timestamp 1644511149
transform 1 0 16836 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1115_
timestamp 1644511149
transform 1 0 31004 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1116_
timestamp 1644511149
transform 1 0 31096 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1117_
timestamp 1644511149
transform 1 0 28152 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 1644511149
transform 1 0 28520 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 1644511149
transform 1 0 25392 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 1644511149
transform 1 0 27232 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1121_
timestamp 1644511149
transform 1 0 22816 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1122_
timestamp 1644511149
transform 1 0 24564 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1123_
timestamp 1644511149
transform 1 0 23368 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1124_
timestamp 1644511149
transform 1 0 20516 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1125_
timestamp 1644511149
transform 1 0 22080 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 1644511149
transform 1 0 16928 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 1644511149
transform 1 0 19504 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1131_
timestamp 1644511149
transform 1 0 21988 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22448 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1133_
timestamp 1644511149
transform 1 0 18400 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1134_
timestamp 1644511149
transform 1 0 19412 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 1644511149
transform 1 0 17204 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1136_
timestamp 1644511149
transform 1 0 19044 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 1644511149
transform 1 0 17848 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 1644511149
transform 1 0 14260 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1139_
timestamp 1644511149
transform 1 0 13524 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1140_
timestamp 1644511149
transform 1 0 12880 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1141_
timestamp 1644511149
transform 1 0 13616 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1142_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1143_
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1144_
timestamp 1644511149
transform 1 0 9108 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1145_
timestamp 1644511149
transform 1 0 8188 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1146_
timestamp 1644511149
transform 1 0 9844 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1147_
timestamp 1644511149
transform 1 0 9108 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1148_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1149_
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1150_
timestamp 1644511149
transform 1 0 11776 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1151_
timestamp 1644511149
transform 1 0 12788 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1152_
timestamp 1644511149
transform 1 0 14076 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1153_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1154_
timestamp 1644511149
transform 1 0 16100 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1155_
timestamp 1644511149
transform 1 0 19964 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1156_
timestamp 1644511149
transform 1 0 21988 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1157_
timestamp 1644511149
transform 1 0 22080 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1644511149
transform 1 0 24656 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1159_
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 1644511149
transform 1 0 30176 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1162_
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1163_
timestamp 1644511149
transform 1 0 18308 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1164__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1165__82
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1166__83
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1167__84
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1168__85
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1169__86
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1170__87
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1171__88
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1172__89
timestamp 1644511149
transform 1 0 10488 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1173__90
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1174__91
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1175__92
timestamp 1644511149
transform 1 0 2116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1176__93
timestamp 1644511149
transform 1 0 33672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1177__94
timestamp 1644511149
transform 1 0 4232 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1178__95
timestamp 1644511149
transform 1 0 1472 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1179__96
timestamp 1644511149
transform 1 0 42688 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1180__97
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1181__98
timestamp 1644511149
transform 1 0 46736 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1182__99
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1183__100
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1184__101
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1185__102
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1186__103
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1187__104
timestamp 1644511149
transform 1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1188__105
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1189__106
timestamp 1644511149
transform 1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1190__107
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1191__108
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1192__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1193__110
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1194__111
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1195__112
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1196__113
timestamp 1644511149
transform 1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1197__114
timestamp 1644511149
transform 1 0 45632 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1198__115
timestamp 1644511149
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1199__116
timestamp 1644511149
transform 1 0 42688 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1200__117
timestamp 1644511149
transform 1 0 45264 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1201__118
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1202__119
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1203__120
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1204__121
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1205__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1206__123
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1207__124
timestamp 1644511149
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1208__125
timestamp 1644511149
transform 1 0 46092 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1209__126
timestamp 1644511149
transform 1 0 18768 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1210__127
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1211__128
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1212__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1213__130
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1214__131
timestamp 1644511149
transform 1 0 1840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1215__132
timestamp 1644511149
transform 1 0 45448 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1216__133
timestamp 1644511149
transform 1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1217__134
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1218__135
timestamp 1644511149
transform 1 0 43792 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1220_
timestamp 1644511149
transform 1 0 27692 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1221_
timestamp 1644511149
transform 1 0 43608 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1222_
timestamp 1644511149
transform 1 0 45816 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1223_
timestamp 1644511149
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1224_
timestamp 1644511149
transform 1 0 43792 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1225_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1226_
timestamp 1644511149
transform 1 0 27140 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1227_
timestamp 1644511149
transform 1 0 38640 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1228_
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1229_
timestamp 1644511149
transform 1 0 31648 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1230_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1231_
timestamp 1644511149
transform 1 0 46276 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1232_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1233_
timestamp 1644511149
transform 1 0 20056 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1234_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1235_
timestamp 1644511149
transform 1 0 25392 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1236_
timestamp 1644511149
transform 1 0 10396 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1237_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1238_
timestamp 1644511149
transform 1 0 46276 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1239_
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1240_
timestamp 1644511149
transform 1 0 32936 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1241_
timestamp 1644511149
transform 1 0 4140 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1242_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1243_
timestamp 1644511149
transform 1 0 42596 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1244_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1245_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1246_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1247_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1248_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1249_
timestamp 1644511149
transform 1 0 7636 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1250_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1251_
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1252_
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1253_
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1254_
timestamp 1644511149
transform 1 0 17848 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1255_
timestamp 1644511149
transform 1 0 16376 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1256_
timestamp 1644511149
transform 1 0 19412 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1257_
timestamp 1644511149
transform 1 0 16836 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1258_
timestamp 1644511149
transform 1 0 15640 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1259_
timestamp 1644511149
transform 1 0 15548 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1260_
timestamp 1644511149
transform 1 0 15364 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1261_
timestamp 1644511149
transform 1 0 15640 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1262_
timestamp 1644511149
transform 1 0 11500 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1263_
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1264_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1265_
timestamp 1644511149
transform 1 0 9292 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1266_
timestamp 1644511149
transform 1 0 11040 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1267_
timestamp 1644511149
transform 1 0 14260 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1268_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1269_
timestamp 1644511149
transform 1 0 11408 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1270_
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1271_
timestamp 1644511149
transform 1 0 11684 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1272_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1273_
timestamp 1644511149
transform 1 0 18308 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1274_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1275_
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1276_
timestamp 1644511149
transform 1 0 39928 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1277_
timestamp 1644511149
transform 1 0 21712 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1278_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1279_
timestamp 1644511149
transform 1 0 33672 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1280_
timestamp 1644511149
transform 1 0 33120 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1281_
timestamp 1644511149
transform 1 0 29348 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1282_
timestamp 1644511149
transform 1 0 32200 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1283_
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1284_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1285_
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1286_
timestamp 1644511149
transform 1 0 46276 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1644511149
transform 1 0 45172 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1644511149
transform 1 0 41216 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1644511149
transform 1 0 42688 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1644511149
transform 1 0 13616 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 13800 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1644511149
transform 1 0 46276 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1309_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1310_
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1311_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1312_
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1313_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1314_
timestamp 1644511149
transform 1 0 42596 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 28152 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 21896 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 22264 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 28336 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1644511149
transform 1 0 46276 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 47932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 47932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1644511149
transform 1 0 44160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1644511149
transform 1 0 46184 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1644511149
transform 1 0 44436 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1644511149
transform 1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1644511149
transform 1 0 40020 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input29
timestamp 1644511149
transform 1 0 47656 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input30
timestamp 1644511149
transform 1 0 47656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input33
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1644511149
transform 1 0 47748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1644511149
transform 1 0 47288 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1644511149
transform 1 0 47840 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1644511149
transform 1 0 12328 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1644511149
transform 1 0 20056 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 14444 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1644511149
transform 1 0 47656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 30728 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 44988 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 27324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1644511149
transform 1 0 11684 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1644511149
transform 1 0 45632 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 46736 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1644511149
transform 1 0 46184 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1644511149
transform 1 0 46184 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1644511149
transform 1 0 46184 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 24104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 6716 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 38548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 39652 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 39928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 37904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 19688 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 20608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 21620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[0\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39100 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 24564 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 46920 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 28244 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 29440 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 15272 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 29348 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2116 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45908 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35880 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 45908 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
